`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p4tmXC8+28B9pJ5HZUg121DZRF6LhciTEerSeem3J9qpChypE0/8Hg9V7+4Xke10
TVe0gQACWkQz4lJNumcNXX56OuSUxiZV34KranuScgr6FzulpL76vsHYY+UTwl/Y
ClsrCbpPC0eVRXg3Iia9smtEmEisbHoxmf8W7qbd5TxwkOMcZ8ZgI0PwDds6JYOz
xxTrUUpkHi5zZQV3PUuJbrYgrwq2JKHcKSoA/3MfECKmUe+BRqJTqKD/EP+JI64E
IoUC+XLUNhlkbL4Yw/MolPy5QZf0zKvaIgR8H43z7v5V/Rieub/tN3VTFa0+y3OZ
0EN23JBszGYFnhN2Lk84qSeilLOim+0IrsJUCIMEseA02BvXb5ONSaDD+wOhOYRB
`protect END_PROTECTED
