`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
stbsi9FrlhrHKbwhb7QvqegKWAEfVWXVRvT5lP/E4bsEwOGJ8kgRHrOyAbo90Drp
S9z6uJGSj+S6PBdI0V1sPi9gEpBNRb65ELScr/gMOEoxa8wWrDJJsWYKGJBcf64v
GzdFhui0HtGHOfCHCc2JuLOX29kvF7DPUQaVSuNNBF3xl1z7hBPthuDUwymXw876
Zpj9d2yMrMcqtOPb76twEHW7MiEpafPujTe5LEthaj8GUxRqPwqMH8oLvujMUsYT
IFd4GJwhFlcovJoEU9sjn+Y2eLAN8xwqTh4hO7OuBL1M3BF1+1fXZ6QtL3p5sMfo
sxSPOumJSsHXhl/hnjQW7VdOBjHAmbQWBZlRXPUnqKcFKjDcia+PcC/0dvanlZeO
Zp+CmU7fyPPhRzvvyZw/hjchMy6TUKC50zyamojOJ2PhXi5bM/O4AWf8RxzqwB0q
+28Bcjjt5n3pkp70gmgeEXTGfpw+99wnrM+zbvxIbtrJDKUHBs+t41XXuv8FPF0Y
4hAGpNk927Z/RbwznYJukucIPLwxqgUCV2P9fJj3yIo=
`protect END_PROTECTED
