`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PJcQs3ALb5lqDcv+SRoWM5byWMOYVlb1l9L32xCodE/F+2tmBB1UBGoOSmpNt92y
0K++VsZjy5d1ARWVcL/l1wsKfzPOyKEY9b32sN5DYUGlnFXodBzm2Lrvbl2l9dst
oDQ6kBRmtWE+bttDVIOBRkokacHHvrXQ4brAyeq1pNVwd+17iDa3AOHDAKmWSFWX
61d0xbjYhmNGOdqtShhRCv4fDLmOI7pr3wyVCHCACytcijxyMjuuDdy0YWHkzWUA
C7wTXunO5VGPdRqVSMcIC7jxjAZeGjbCRSFzOsjDtNpupPx89GvQcJOHrGi+Xxr3
0n3T1M7W4XuFYgq4DztO4J+D+T8tMU/rI3ScRhODFbV8WVeGXbw82RolBgtY+OQL
nLGmffboreDTqDzlSzuA7NIeMciHklyzehfEisMKv0aG+wHmnwJspkdb10+IKQtO
3qKB8UPch91A1WqytUUYIpzBRoHmUYPJeuqCvmzwRzqwPIwb/YwAf7G6oPywKHft
c5YZ6WoWkFDSMdCoG04d0Wst5RXM5VSBobwcZphkeC7E8Ktp/MVfrSvutmfKHTGq
QNTZAmd+SvssEzkFu7yZOu51FMVJPwUNTnHyzzQJioTxz/Z7Zs3zB6eug1jB7IHq
gnyIYU3ZoTs5fJaMbU5EImRc0GgflYq4ZeE21dPtY6DZHDho9ylHLZZOWVuqFu1p
EwpB8ZCZDgvsK2c1EP29p4gpsDjbb/ktWsKWQchRPPUaSeSPIpJAkPsIRaNwYAQx
OmMAmkGQn2s1XF9PtUI38Y8V2ZIdXNCgZvKLqhnNA1gwGGdW8gAXhKI7YhSmYVdX
VIY2p2omXCXrLHDtnk0UhfwxGyrFmWud8LkyKTkf9aU2p5c8LMC+j1/0TtCGKBAd
PUmdD0NHLa0f6lvJFylUeeWvxOJHRWpFhcTg0J97gDRbptcIQq/eU6vJIPjrQeAz
dxReQZXw52vXB8xcv82lnVvMcmH1icxmId1MAfiUDHYLXcL+yDIzk0BEyDV3zQwa
BHUR3eXI+yXwyzGvtwTvIhOq30RJneQeFEKahwyXm7kxmDGd1fKLuJslQaRiM2lX
uMrtp4Mbw7Mc6ZQZk9ulwPjzRJSTmAGOLBWPVdJaXQObaS8pia5QdMUr23wxdQ1j
GpJ1G4QD/og+tFnXrb5MEFdNuN8iOltDh+MADKXjatlSbXONAF1DQidwLSSDAjMe
07A3DKaD67OL8g1IjH9CJoQI7i3kRlTjNfgk+UMXSWyL1qmNy0QaVjVD0uVUBbMW
uxtjTVklFGbjXSVlipSnaSZUTsCsqLhE96q2Eof8fmZIlfc0Vam/uO0zL5wvGzmp
If5Gh4jcEqZO1dGO0ANfZcqJUeh41dLWGai7YTKRFaVFZHHZ1tLJJBzWWxuF3l7A
6pGZtADIVlXFIs/xK6RSqqW5hQ4pXJ1DdDwIcjxqddcBebepYZdYVYpoxy/VfnhY
ignIEQuH+gTOv2ZYknyY+K1S7Rp2tCbQF/3pUS0c9Fsf7gPMlVtj+JqlJV5nQa+j
w9wbRVIX18WQR50PCU8zZiJTNry6+JiZBZl9z9oEoO7bh4zHb4yapM6bjbeeTmQ1
fjP9aM5XS99zhCaRwR7JomVTpOaAxNJK6ZZbypNlLs3YvxlvgGjglUwT+DMtuTWZ
o+S/AllU4K5mFErH4p6jkNyq2+u4AOKbc1m6/QA5hmAxgga1AzcM8rV52/adaU4U
7EIdLmyXV24UBeojcIPr0qW7k44G/TjdvWA+JRopJswAsP9s9rasHaXYwf5IV6co
5q02NGpVzM0Pt+YJH0V4RPferqs3nl4YX7AYv4Vb53DMn+wUHWPqs8PmGu0+wx6N
csqdD9ryqhwi+NnlFzZcfbpMilnZr9aqQ9DZZIwuFeCM0mlHnY/Q8jERrwtlKk+e
uJ6S4n+pE4gw72XD31mMh/j6xWIjPtOIp+obMXZX9PL3U+EKMBTU9jyNwEIt9ZHG
sQVqF7g1/pWKZCderZI0zyavperYQ/i4NTnYQtQjFgNV0X6FaBi69Zp9Zo+lRaIY
9wLHGgWC3dyJZZZnvgxo3XZKnzSU+cLBk9Yxm5kGl3MMp3jIlibkQiI6SS0GOOkW
skeaH7oLQmkibT781dpDAeXl19yz58stcqc/d7DUxETd5m2NafqVKd+tVZ+Svp8j
FbblFILDD5b0ZmBeVY0XRcBCofLHnGl+zdhWK7C2yp57aokganmC8UuHaep2adHW
buRmHpEfkjfczzs1Q0eL5rh7jPd79ovOaD6WTwO+JtPOaEwvmF6yQ3Lhmu0PyypA
ApPsFVFaHadGGmLte81eCvtWHv+cpVs0j0s6LcMXY5mNINiitVeFV4UIUmrId+HS
ggm7BZrnoGDo2sUJceomODR00MEpnIbRe543wEEAOVed49DXgjn9kkqX8oc5GgmK
1fkX4mZvN+ESEcVkjaem+GJOepkl8lXWQZOWYA6pSCOkHT5STO8b3ejZl+vrw2vc
yY5WxGHL13TfkjPD4flTCN1YUDa+FyC2udPClQtoi9CoqspY/2wRoZjegIanFNBV
tsc/P0VhhlbF95ED+2QTDCwTb2pob39Lt6Vbu1AhlGcIV+x07hX6IgaeAkc5fdDb
WLRCLcM8c+5P3aPvzeXwEVSKVXWbzsz2q6lANTiaLq+GJEOWulHpWFKEkXPPoyqK
6aw6xkykUWoZIXigO/1zzOFvRjraXFblB0VVFOH3JtiajPddb6bE2Q/yTVJKDLYQ
nPn2Owa+F7EYwkTxAMbUXoio1NZR9ImuuMslFLn5RjOR41Upd4+ROKz8C5cdbdnb
Qs4mComE5yGxppJCQFnNXhJwX8RLT68dyxKnMIizDpTCsTa/I44Tr/dTRby7ObG0
P18/TeDYIg2JAidw3P/DnHe0MfC2nTYzjEyvcynBRm9LDZhrTq/j58WeYzxnOlc2
d5MhrSygiY1OFNlLgjMVngbpIjK4xD3t5v2Y8e0l7NDCwalRAbWx7WqXh+uWA5lW
1APiUQMH1/apswTvcpvrmX+1PjNQXI35PQgz/uWyuzhxyldU+2L9p3pe8FfFTEPP
68XbwySNXkZjADDHhLJAISlja7b773J9hC3Td/04mAtRM4YHVRf3/CpUX3PQ4jc1
AFyP8rqJjtNrGWSVwrHka/tHbXXf+0HQzYfrAsWgV5XB8ytwOxpIchEeKQUKuRmD
cnBIjms0M3uAF1rxhjR7Gv7JCFTfaSr4dhnekzdhAVTLaAM9Vbng6RKO3niZe+0y
1soAjLOcOsjaVT8hs07ZMO1D8GWVxkt97UpSK1DzDOlFhs4rjeqV35ypiv4OyCGl
bcSFk3RKZaMM9AyG1SgJx4zVwH6bGew1YVEkRyeLktZQWES32TkWpigBcbVyb3Pu
heRxKVSdYkAXWXAcmaehwI7jUdQjZrJpjOqGXHi/JYBNsZ5Z0QBcum10KfjjbFy5
9MPs6u649ZLnowf3MxgUYaT0PWQrxpgRhGTJvqJhQ1FpRlxk4bPs33avMeC0OnBz
jsmzxGTkhn8O61OPDZCPuHaNnXKzVzE3rclWcNMdeQpNnBrjg7PtxM6pUFh5FDoy
9cYjjctEtzh+u6ty8wegs+MkkVszWciEtdfLQTemGrR3enXWE3hgdUu+7s7QqjVH
R6EL8A0zHZneWp95q5gXhHksAITobAxle8NvQi+TyFdhlIgVhzdsP562oWLUuqUw
kerfrvwzaKt1QWrglZg5XdQREVCxr5Pt+BMwdNkeQixByu/g/RhCm3WaPJVjqEpv
BgDm++e3FnxvqO0Pb89kQJCXsbOmvvInkWWLkJ+spMsKqZWdmAkutRTsSoXoqQms
9G4jKoBIRreo5PLe7+f88dccYpZut29O/ncW2Sg3nDolei2YxqfHd9fb2dZxkgs+
71Cx0pYeykVecfW4LwP9w788ceiKbnyO9iI+viuwJIh0wZFYH6Ag5Fo3cqbbyKFI
q1WkhKqhuzDvvDDnjY7sj5WxbKFDdKK91dv1CZ1PxBiH1imxXKT9e5f1zyH39K0O
1C6d6I5Cv6boa9mQSr/jMdSg8havKdxvjXKrhzbgZyHno6GuaykiMyXji93BPWAq
jueAWQn/JrlLG/DNqpg7b6yqlFFAALa9Eo4AE9Dz32hc/IGC1tuzskBqutxZRVwN
8lHRjLb1JGpxe8Pjzept5hYkCHbDqoKKohTokK7tJPgUKHrTwx1tkdKDn9BmIpZJ
laLhx40zIH0jHpbkpk2bpoaB2YRGL5ns873hxwcSHyxPSRwyEzkHHZef91JF28Hx
vG+oQetK+gkALMD1LsfEfkZthNbUAwlORtKeL5TSLS5uuRAJ5hQ1p1j1zswLt/I7
kiKQa12ZlIGmtbXnh4pr6vy0dSjhhTKVwd9h3Dd5AiHK2eLwdLCUwdsDXFwFZQO1
YQmXuDmkY9Uv0zm/yn1FfYWtFbsrLuG8wA9VuCNvn1znqoC8RvRt0Cv+Gs/Vs9pG
9bLbq730gHMDd31RbIG+2Sl9xsu335ymt5b/29ni8nGBbKSHKmJPpuWHEGmW5ky7
oX2L4FPi9HzpPM78wlj41A1W8E5vblgCRgzfZB9NzjqxDcVXYVwJnm5DrQ//7yEA
oUBdrRVHMtgg4QE0xmT3I6iILLpxc1V8CfTyC2CAfi4mXA3du1BiMXu0Z0J4p4qy
aYMyFeO3Oo70GTbJKVzshqKQ8w9EuN1jdGshNM77pLQAPTaFZhLqM7mKY4aElkpe
JRobYWwcaoOB3ZxoP5nf1DESdaGPkwbVZe07EUw2hQAwDcE0Mjq6nFCJ0nhD80Y+
X/KS7UFmkljlRc33yXH7+8Jk0s1UbMhraeOsq3B0h+Ey17IUftExKT7c7YXdO4pa
Ejz1YS4lSyhmcqtpIeg9NqwvkiG1uxh4/xrUv7olN7qVJvbIgxNRebC1ZZwNnIig
ASYvaQUbMTwhrHAunm+fLyDBOlTVKuFgvacocy5FCzPYl2K880woKLgV5xO66MPM
uUGgBmivqux0avim5PlS4NUoJU3Qgq6Li3mYh0sRDtxL61z9Zvy/VYMbibjNUzTP
Tm5aGi2WKQ7zz9wQfx6KkrThVo3CWm/2Ttmc0NaP9/JL6GdTZVaxiC2/HrDHiBmk
BVsjAiOkjz0AjhW8MyF1Y8yVIj73YTfemWyCw59+1KaamhabTCaRE+ZBwjFdytx1
4R9j7OMmxjhjDUrzW+BS4D16gnE+Q4t6zdFFc8YMYHZCeJwmpEfWu2d69rf3sSey
EWMFoNt+R0dfmtuNK496L1eeyyssMR+ULqCwYI4hOWU0vaOmqfuWiETXnJjIVApD
k76VvEBVv22KzUM/8V7yFsMMMfsm9ndylpFruD4PxyWnv1KiePU+mIGl64r8M50D
9kz1VmJnj8jfPo2h8nea1ZAXVIw/G/lyr3zBC25S+OG/URI9fv4pEiT/rVJFnzgJ
Njw+POvBWqDXrVEtZiR06NeGadmQVLpB9UAuNYIpSipe7/ydmBEktbleUllwWY1X
arjnchE1O03VYqXOBpPSb4k8s97FtCnb3aoiDK6CXxbtWg0T9gM7P8+ccoonthnC
594dAwBbIzA6JTTNPITeyuPbkzFlQYOstrGJD5bLuxoY2gbS+n493bwuooGa4rDD
m8HU09wHYb3d12gRe+iWZyPsmHCakLfmDxKznLjoIBFrGH+8nDEw54fHsII2fBQ2
nvsO2fDiJSL5ovQNmvfXwMcM8o7aWme1O9rkHB8+JLJuY02IZOWqfxRvY3IFwdsL
/5Ob7NM3P+pFoyeS5f+hy1mgpzK3ZdHs+hgcoY/KCB51BHkEtxPhp5bklgF4ZlUX
QnLIYTPbBgWS9LqZQDDZnz8S0W4oS5ukgJJDIGECrK5gg4HWauljtRAjzSnMIE7S
Mciom6dzzOKFEGagOGuErpenheOVPjLfY4e4UEt+NUkuY91PeU1AjqaVWZWuUXF6
XIBzHNhhu3D/0+SLFpUCLQ+K6H89aaTL7VnL/4wHCjMUn3vOBR82d6N8AYQI0rjR
OOUX1jUnIoTr3JgfEEE1wua/JIQYEAJF2n91vXg/89NxO3QPP+f/PNkFitCcUz7J
uj6Mwa5axpWW6BMpS21hQtKhccZckzI0ELuRQJewcQcQjdMqu3yhiW416H6DTAtX
Gf67hjv6pcy0F81dXwnaPiBDd68P2K64YvhQHrtEqXQOkx4HkPj8mTolvyIrOorG
q02IRd+FS6VCoDvJh49+pKVsFaDIdyEB+I/WMxiHkDHzT2SlpYXX4sXMiYjp/JOY
i2IoFhjHyMpVdVmwiuTgya1u3YEIz7TaVICYRPA/wnBFvVJKI+OZOw51h+wypxmc
tipssPSAvDHftq3NP5vC9Nuz3O7WZzcVvBDYmrncUlmn0TP921QoIqOt/0KfRYdw
ZmfMLKQzYmyGJe0ogwt1gjOgiCqDDIXsh2H7kscfs8DEwB+rHeRmrdkIOqbgv6XB
if100cFSL6GhQWr93uuILphnS4YXeQISSmGQt1VsWpBWK6xfab7MGP9fDYPhlCGz
+rCXpyjNlnOqlE8fa3hXSXTMwTqnO21TbROyveQ+/L6KhA0KIkCC7VMsuX1cnEpx
Nugp8BXx9uwpQdAHcZiMV6nuZnCMabAxc1/T/5oxLeXOjaapGGGlr/plHMXTpF8D
Ep6k3D3C+RCF2C9DAxN0NnfHs3n70J4EOHofsRmVUkr7Esqyd696kmOiWMyCeO/u
EhPetMuwc5PHQ41j8qTqrWClWRX1H6pk07H7MN9QJf27A9sgdbMcgVWjDFEa6oIF
8JzQ/T2mStr2aYZ5nbhwFdwulAXG5/FT1ii2WiXtAP4fgvcZNM+YRfI+l1F8+b5N
hil1IQF97CNC049b8TwzvYBHfGbdnrpT1yhv5J5cfCznsYBkN1vf8KCdulbl/eaE
GigOQelT+lRKchDkUyC4G46jBvTIZEnhBDCnhdT2K6SpoADENkYkHqR0XDzqKCzp
l4CYmnZqczaZY8Mu/lj7aYUIM40AWvkgtSKB3GxmA5RbKxHdRSGqVToQCxWshODU
e2m3cNzQ3YTCVZ3h4XM5EOA9NdHiKre5Fl+BHd52+ZYB982uNsL/z9hFeLt9w5NR
Rh+r2z1vO5/1onDZqPlF+aelxBpmRYe+SP9Z1LMccnFIDIEl1DkRwwJ0MzJCOiTv
7hO9XMs+Mn0G65uv979SaHq0JEpOzFMyucZVPE4XuCNm9s9bS6RMC7Sf67jSQmav
hArL1TAAAM0xxtI8dV1l9zrk7fYy+uvfuU6kUROh5fI=
`protect END_PROTECTED
