`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QMHkNx2yBWjaFEQu3b6KaqESTIqXAWzXwG5H3qt1TZVTQC91kS411nCQZzif7eFo
+fCNwX+be44NUehicP7sr7bZ7rJwAzGilBYkiLPZN0luzsUXtSqzviI9MVEni/D5
IZB8Dgk+W7I2HpJqNbvWYXoni1IcexMruWQZ/uELy3X3aUwGvvAYypJauK6Rno9I
wjEcfKJR/tLN/CI0AP32gm7fnDKyzBrU5YtX9gjkZRnHXAlMQcwHEhUoHTrel1Rq
mcddMbvw2eSH3WYKH0DiQpfTCSkKwDIaURRhgU/ju6mYSlRcdBJMLXSDnYOUOPsr
JtpkAqEg1XY+ikHn8vVOyDOAqNoK2/SdwvN/Y4oPLk8Q2T6RmyuYOcer+VeTA7wV
pZ4G8/J15Pt7h6/flOc7oa1cf/MtqD9imuKVVDM2R6HmeSP8gNbh728KBcgK4Ke5
ACyd/JwsngNYF7I5PAYtk//vd/pcno4CwoGQwehe1Uj+mRq7zPjjlPhqqRAiOpG1
oevF4scEzItXJwVmyP8YIBTHqlBV9YzeRNvdxl96xRqqqAE2N4xwF/YMPfY34Z9C
b3FoH77vOsM1QTwMJy9H53CVcKOh+tJx/ZRBWzNLtXfVg6OrFahFjdQ4gFD7TuaG
b+zRwGBhQ3UMxcZGlDFrdyChCFOGohddHX8mE1zHgV5ltpthrr7qPG/g9cMs8JnK
H6VIT3EM6uu2Z4G2wvzFB80pR7fFoHz9yCEPfpQ98oIFvV2+a5KXSGySz9y8aHhU
DJOV/yX1k/9XGA1BsVZQ0ep8fbeacnj8zrsPNWSfOhQ7ppUL3sU/jwz1AjuYfhjo
PHYEzoFV/MawDOKPVWUYbePvK9QcZKvOOnRZjI9InwxGetKZLT2P3LWZLss3wnNZ
XphtA5ka+/Ew0PtVkszj4XF2m2x1Ig8kMo01rM+Oxz+QzuO2yptYOoSTGaBTPoJz
vk/Pdp/w5I+4QGx/+5aGDeoN5isy+BFlwPpIsVUmq4ef31jEJYpiEjR6yg+ytHro
kgEiZSiYz1R1YgpkZRczS308B18Z+tlnywPWQi+wV2xNCQRjAeCq7u/rVE7mVeRw
ducR1JKDFX76Xe0hqiYL8Ar4dHsTHkKBH8lcoxaw9stfxlaIzdTtNsLwLetsg+ck
s50OH+8S+LfNUfvLCjb4q2gLHCQsGQ/darivBFciSN3rMwVXpTYDKo1QTwvgMmEC
/eRYN/dOS0PKA2wPbkn/2q7vG8IuWtBBMfi1T+cnC6PCz/LtmzYhhSTAZOySBlWq
Tetqr7HxIPaANZZZHoalejNn/pEs515l3DPn0D9VLzUahL9nmeXlBsyeeMwEoPHc
riGF/Ma+gKSMhdg660OK3aJy7B5MHDqGDeYqsaWD4o71NqG4khrJq9PhluHJHCsu
ZHRBMdl9Yege4n4yrMMZxBZZj+YT+vPofsUbfkLsX93YEEtFs2riOFYTGH7X7OnI
/Cru8rzGY3YsBT5YUBs+sTkd6mZ2Qh4wjRwB+m8I/I1YVpyzO2pBfz7xF6cpYQQi
ylsecwtm/aDGF4MnRZxGnWWj5LF+Z4f3kz6scZIpbZgy2p8l82LNL9E2Q9qhH5DV
A/hVErIE3GWucgdhHWzLRVUCei6YzMXybndTu+TAZ0v/HOOn0SQeLRxCIOXRoLNp
+aKRy06QjgCqAa1zYGHJQzrM4ABATOCVpwZxZAkHIqVU68xkZgORcQY2nWzWB2/4
e7ui48VZtEGZ6EYFTx9H11tomt7OowxCXVMYDZTtVSzMg5HvcHZy0+ypEUO3fshO
nVEVGdJGJViSVY2ZCLBV8nutdkqWxgwg5BxfYaWeYLlnyjK/y6E2sLFM9YE4X/Aa
zi9zDU6ieeuNT1bzFt3hQ+7YMp7oPsKOISa0oLN2DPmW2cMErzTceEZev/7yqllW
I976Ny+spRmz94BPag82uw0ZF+POjMzRNh8Ydibh/Vb/y15WFzLpV7vgDDopF7Zd
A5RWZHeZnjpZA7gk0WyoY4WpQKAlL2bZyItTd3ArYqkRpNVeJRLfwXwK+2jaDI41
R0XviLKG+qJXNtGI7lmSqL8RAzN1vbr5ZYNqWhxJHbKKX3cG3hJY0gFS6tJgi12B
gH3FqE4RdUEmfDnLoZrbp+CweIOoDakxRVVJBNqcj0XpXUeU1/3Sm47xrTzJlzmc
yuz3vt2rwqF7i7KLXgsms0SIGyNcuMv5nIM6r7suq1dDGKkSmc7QAE25g9U+DNlv
Lct3PjQeqaNOrMbbC0xucuhDb8rAzo/tMfRD/3FC6WLVV5RCba4UsQpCkke46LUc
9uCFncb/MYnvi6K5BaQNJM2osXJ+zen7Z1hRS5beV4kAYlFuicEgczMtNJM4WVe1
V4h4y9gjF483MVqBw/8aqfKUp4dCvQj2zLk5oYYgyBdHJcw65/x/zwKQf/rvw7Bo
GHVOAW8FhvOp9K7/SvapAjS2g4ldZtovXvaWAHbICujBrjtN+59KiJFiQ/G1SC7x
UBFRYgyNtf6dsIlpPD3zhd0rIRcjuE/vOOYY+i3Yefyl0AS2DPXER0BwjJVE32Sq
koZHHVJzk/AKYcw/ZTjR7gA392zWvIZ2NwDKfE2JFKXDPIiDqHmJ4Pou6kPozcoi
Eam4NvH5OouHpi50OvNhzXh5Aq7dnmkBPyX9BIsWQRnPZ9nUFtylKL/s3b4eG0yU
KGWoSUmtJWM71QDZXzuvJKNsj0uMUleTcfwltWcSDx4w2thoFuwC6SKvzI3HNfYO
3adAgW6FdmxQA2Fm4No4UUhHWNa2qdukpFRrXZrfvkLRVFZINAcCFY1QeADMLFzO
KvZMKDEV/Emj6QeIpVNq3lPwcSf144JqYO7hp9UN10gRF3eiMmwLCNuY4K6ZDfe0
V47Hoc1EkzamS/FKiA1qvf/oyz7G1tpXaRg3/zRPKF0jp2Kmf/SWBRZIubE4mvPE
SR0+km4gOQp4EVmU1TYxzzDluvh1rXgC3Lp+1plVJrEQ2tNSjCw+bhXf3GqgMQBj
BfR6ww+GNV1DB4Z0/wsRReBko0w2osbZkuYDJwrED9yjCZk0cOIuAaFJtPQAW4xy
s9DKr1ZbrDyIkcCVHibWs1N9xhEFVWXpIIRzrla7dNNQb0Fz9cdFZXZXiZdlwrG2
rmEPsbtRiBx3nq5maRUftWlz9ivq+RP0c0elJkLpAO8pMv6z/fNmL9PFxDWPpw3A
ptOcbufs0+0cWtXW0ueuS2o868lkgQ8C7oAHiRC/h8lLbgZrewRlmeh/nlbzmXXx
foRqMc64jYRsTsgaFBplvBKG3T4cWugikxC5ICbLKCd3f6Xc4w+Iex2Ft91773Aq
dGVeyBcXZ9e4CHpN84B6T44NDprq6Il5/vibY4hKPxATwMAO5dgDRWx+YrvnOuOs
rQaVQHJ98Ucht91bvPEqyNE0Fma9pnTQsJ4hpfqVD7u/ZBy+43DRgHY3BgXeFTBN
oj8kXLlsZxWFXlsNCEgj1deHwYQi/oTJvimlKtctmZpi8s1lCuI9zLzPt/f9u2Om
LNgG24gOUGKGK9PlzCfn1lJWXETkWM/mtwceM5hExx8L6VKCjka9G/c321Pn5e2/
1sVRuSxSSfiOadvpqW1E1f+UpMCYqs6C0keA63DEf0cCjequMbQk1i65/gTvDfpf
CsJACu6jCqJelyKMkkC8jGtVCZ3esuxhwd8weTl0gFL9dX89oG4a1H53xSDHbzTH
seGef9OvDPSJ0pTisR7MIbjMYoB4ZGbBDsMLRdV7mZsdJKitm/tUNt12u60smnJx
eWb/afNi9SjiBAztIMmTB9NoY10BhgqVzP9vGsuLDb9IEFleT2FYK9IQWubaCpEC
pjTJebEC/XjdBV0H/Pw8mvvk+VuRgTxI7ls1U1Fe+I7gZaBjFp90EXy7qJ9yS+xM
wHrb3odU8d838n4acoq06wEltGws7V0a1xnvFfQPFCpeixPOCVQjuEyE9QSamWLM
4Jqlj/owdWvgRIiq5hc9OxJhpODdsEZIfKOJU/4vVEGOWzHj+Z+Uedroj90Tx/aS
QBGK1YbsmjvIwXiUCw9gX9Gdc/9C0R+cxmL9NyDxtiM4UAXx0MYi6a+/mVGZM6gn
sDMCRUqMetIPfCnlQ0aDe1Xkt6QfYT4PqhNiU4bJv185zpz9GF3besyuqJn5looH
pxmtsY7rjifdXxdFYpZlGWmeYam5Z4Gz4r6iyBdLEfQveQQg9S7Q6ZULj0m5S2IX
vuT0EDcsbNR9IkL9lAFMyWyGw41HgLUBstw/kCSZIt3FsNbcKmrz++SfRpkKig9h
TDvYS9KDqDSqjj3bkZ2MnQFZ2Bf+kT8HQIfyz5u2APNkWjzrha6uBsSHm2r4eTj+
RQ3uZY6zfmxVnyiGzZ9t7TzW1z8kXPEMCqJU3jKL3NbTrzO1YGLaELmQHqi+gAAb
VJ9++6FRDzdXSq8eCeGsniTaZsukcWvuUC0/l5nBiuSrHUMwzrA/bhW+1hRObiV8
vtjG1h1E8bzb1D/corvis0Tif675bgWOLGofcat/0eDOvyCJYsp2W37BNMzz8SVY
0gzZuexjp9tnxmLh3+jFJiCpgDGgnXNrwvbCubWjgvGGXj7r7z1J21hFSF6q0YoM
5VtneSWA2efkM4QX0CyeRerKsg5BNuX+f0MRWL7CMp+9Qphjw0LIfQOgW9R1mlLV
K4tg346Gk0Nt6v98YJQ7SGyzRctzi2z9H59DQf2f+V5Ds39IPEIbmWTaaaMNlgc8
L2w+IjZ/L5CfPh9Lmzc69DLlY4DJpx/+uBi3IHZAqj5ikb2aW47IxxY1PUVi9wfl
LmmKzjcVX8bcQJGJRpykamXGeCCQKDVf+nzqR0BNdvaJdpbyS7qjmiEuUwyUjaht
Or9ad+nMU3rMy+RAgZx/2/lAY9it+me8jWJEo/v0l0NnRXEjZ2zqpbCMJ4AHFUKG
XQPif3AxgodOj7Of8b6q/g7r6LnXEM1M3ngbu8wQfXjre0LkN9soVB1R5Z+rDZ+F
2yBGtRb16seqMUJLOmI9XiJFHj756sAhopYuhMUAGfNYsTfwcdoxxFEs2wDcGmY2
tUVX1XTnFWQybKlSFBNs7dflbv8acN70nfrZllyxpPgNulN3yRxsCpIoNvDFVLIO
dZE6MkWjnrXxlSxDbU1/VwRKE0uQDUHq9hYhktJxUqY+36fDMMcbY3oWHWhuHjjV
ZZ0/qe2ApWbHlANBD8DxjjZLUB1MHBUT2rYyF5YK7idaCT2twMqz2IVr7jQ5+7zM
pGpvk6cs3q7wJLAtLJuFsyM5p6JEXj05vCWGQqGLoD5aiOygpdmVFpgDYf2sRin3
lFuKJmoqBe/23Jpm0wK33vluepkCRsyM614ky0/FVJvG5YhZ3pWKe2Sn9ZGtu4Hi
J2x/3orgZCBJSTUV1ErBmmDulCe5/OIth82xXp9OfPMALCGfcSogMlYRvUus8ZwU
X1NdZX5sMmJka/qv+nHXhSOJ9rbtRPW6mtwj0xZIpos4YpdpA24MhCCGuU+CzrhW
llbHqwLint5UByTRyEZQtbp7UI2N9to2QTCtK6P9fbd9UdPziTNa3gh2p1thBdLq
bkJz5/vFaYF2G7CMeuHAEN+/QuJxsfH/epNZ8Og4Jhn0D0MJ7OSE20lDm1Xilywr
WBdm/aOQBCz+3INwYQg9IynzIX3VMCos5dfC1RkYfHvZYMy35F/yhBHU0+zYtQpl
wOOdNHWPDKVGuEbqJsGuWRZmxXD4qqA3vhYllFevbaATlNIeqyS4ThtI/pLsdPSq
ML5RUxIoLdfrAn1g5BQzf/430PIG1Oai1hLKSX9TAZuf8VKJNYOK9RrMlN2VoVT8
PcWmRq/HvGpYFll8xJ6Ob5FyFsbCQvyxFbVeUPmBVlgNDpTjgovC1cgNyce2au2l
T43yxYEDF0XpeZWl3BWxAa4k4kOL32Tekh/3g4vbfh9v+FkiOzdvYmw9Neu+W9xl
DVOqS8NTd7SXzYLsfE3wwKzfL1hUzayq0H2j44JhJksIAY+Ys6Xw3j4K1yjMv04l
Rq3FZLGrT0F3G3Cbr18Pbj9wKs2dRQhb2rDoyTNqf1XKcilMZ1bCUO66PYW6yKpw
6CNTakAKswVE8K/w47VYKhIUmAMHtjhrpfYoHO+v5KJOxYF3/o3MKE87DYC2TV5N
pmg/6G7WON6QWsg9mDELVTCdqIaSzZZnrL94cWGEPKy+Y8ZnySs+M2VebaOBwEfd
OYTlnG3wcwto3bTjRiFv7XV+mwOx2A4w5j3hRVWZ0bLQSdIecDf5kioMFAxBp/62
GP8i3VDrHAhrStCKUrQ7VSUrCzuDPb2tUDCWEBTXlPXPTuAFiLHcNvgjT4I1yX6o
ElRRZFryucDps+7QBIsciA8G4h2mHD//JCC1yDLzgeWVf3AXWMPSONIa5xc2VzvU
Bh9EaQTudU+X5JxjyaQjrBh0Gm2Qt9v35Srpyy7IwmQqCJhQW0hendgsVjAhSktY
0oe9InX5l/bXI8j/QyulAnF+qF5/m44utZ0Ud3pH/1FdoDDYi0gA8068Jb+5XELd
26zjI9JKZmWVSZzDwnnuarumXWuC4GBNWEwh2ud/XXXV5YU8403viTIqPC79lcsv
Q9EVxNWAqH6146Lf4wB2QzsLuBB3mn3dv15Rb5mP0B/gai8YRQcLW2ZmMYr9uRD2
gvL2ns41NMNo31biTyUyt7DsepfNj1XVdgWCB+CuxoNnZTyuw/cYABcfX3I5VFSc
/g3FDvYhno7J3JC7FXUoVZJ7zguvPLZAt7+tu9xoduQUI4PmRbM1+5/RN5/1gDTt
x8o8jxvrF/TtWiro2L3NSCXNyvhxfoe/oY/3Q884BMC430vhuXcK1pclG8Qvd6cV
DSomXg+AetWstr94Nr1/m5UQrDABt6TcUgTRdAYVz3Jr1EYmBCHfPsWvJRdUYMEy
m9kGZW6rl8+H7bkfWPJEIW6cI3sT1PuEDz9AMoF0wBa7o8Y6wHyieZfq1CKb8HkU
EJUUJNZZqVFPkhADiv83+SbjUaqS6YV14YpnRtYYArFCMyMUOitJa9/4aPBsYDXE
+hiOgT3fsjyFc262uUbqBiYTLWB5peXaRmo1NimM7K06UnyCROC0//uTT1mzlprJ
KdMg1Amwwm+xI7hpXLFYhw7h3XZT677PJF3YhiSQe9lqZ2FZzclucKZ2LpzBDnha
D3k0yT0AkJ1r+/SbEDdEsckZ2eEaS/qsLpQ77aKZRDJ6axoO9AB7ZsDyzzkLEBzC
TLDKYeEH/DGDuHGoZaRYoD1B+8l9e7T2ZO4dDJbJp5fwVwjj560KP+cnG25QU8jG
1TOHVmqH5Ti0FvVKSKKwfOQMGFHd5wKTl5ir90NPhHRrlE+OAihB2aFMzSIlyI28
VzhrcNmOdKhc9KP+2AUp2CIWGhCddLke+k5rTaRPu1mKKh+2J8OyagXMvdF64hDu
FGFoe/FdwYBJgcvt6QR+MCuZZqYoKMFFp6ACJ5JPYU0ZD+Ektj3HACAmU1rz8iuU
RdRmcEGO6Yij9tE5diGNOjXT73jv0m4Y9L2t57zYJ+4SYGGhNDPhhFC36XXk1cws
MJ0rM+Y3nPmxOC2yqprxAhYxVFIN/FFqmt4lWiaMb/qZyEeBJNL92e8ZuZBpwQKN
5a5FT1RSWPqDUZ7SHyv1KKxn0OvtBnuRYxbKCZRMFqIXVgf1qRraMEwqDqtyTMLU
koOEOzcCD8CdHWPqL8czXhQcbOYL5iYFak6BjJU2G6/2xIdDQdmWZ5lt4UZe2C7Q
v5qal9sN5u7wIZG2IQarsxHjlpGH6BwzdpgKmPu86pnZgL4+tMAx4meiJZn9IYg4
QHIax0O3WcqIMfo/+TZPcsIwcOZnAy57CxXVI+v+Uq+R/4iuYneJMX6ews2XZG31
RM2hEwmBZvZ/DT4GQbm4SMMY9pYQiIEMghVzOqOxtxy9qFP9tHzdMehyNcWgyujB
+1LIJh43L0u7854byTMXo8PQUoQrxpJ8XXcAyfU59oi+70mI9sEjlyyKxE+i8xkd
2V797FA4rhw9n8P8KfGdYDjHZJdcKq+O8DJknMU2+KsOIJdPkywFtnf/SlOUuhNU
SteNrN7wmWL48fdimUwbweh+LFNpOePcTJvHwBAH9mnRm6Wj+CMrVSH12X9MLpZP
qqjgC+/HFSm/DEPEO4oTdA/paEYJGWMU+aj3Wf4khrbR15FGEhop02XW/kkRNpY+
OHZk88IkLEUSMV2URWyjqDQMK699DIFKC9SX7+qKjYwgpazWvQ5yQn5OAIWqBp3n
/aitMRpvD6toD0+zrr/1Icf472G2mzS4lJ3sPzSWa7b8NBxG9O4mJw63763R5wdK
kopVM5UNN/sXg9EUx8zUL2wDF2DZ3zyyjvfBEzuSnbHQXf8A35I4jCd0uysnmjpD
Kmb+UK45fUopVpYzLYdOzWETMR10m30BHumUU+t47NltC8d4GT3jcIuYzPkGI0pX
5cnqCCem7cDwgifWUx22M3aG3+nUDXgd39sEqHbRxJPEqMNA9fNLKV3IhCr/9/kI
bdTJXy5s50nW2KfUELLfbQuy+ApQ0Gy3WliRaCUnj13xj397lvz0KAKtaYMde3u6
mY58m60EFniUVcubbemPu5xeEiZ9j5pNXAkwpupvUhXMB+74DgLMuOeA956Z2qSS
L/fnylQhC7DTYsSq1RBuhUnlwxr8Owr/Aa/eiSrP6nD7CmiRw41pEwmgwAwIi1rW
PKD21bfSEZYl6wM5z9Yp4N3jAzQF5Xc0h6zIJbt4nM9SxhxTqQNq61H03403RY/k
cDLgtMbOibvJVYCBTxMs4/4Vz2HJh28yK8Sf1eri042O25TwwMTqwUerPx5zr+R2
JyLZ9tamEd5YM2L+VT28D8fS/uYooBo6BxoSVH+ptqo6PfTpfUplX+EXZYuFtWO6
PcreWt2AHTMyMv7rDY+UAzqNQeDXbUIGGCSsQ67CJXknrUwcA6FanGsR8zeAaWxn
7qUjowriMdJcW3cVa8kkDYaKXchzDz1Yh321ZNRl4Xxf6OpWJFEduMm47doiv2an
E08khUT2m+1C++ITuK3dssmIiZLDXB1xdS6KJ9Nft/m2lw0mzK49y/a7qoM6hv4f
C5mTddEDcbgrbT+yvsxpk1tnzKks614sn4b7pp1bufOeTWQDwKfpH+p4QoCMv0HV
jI88xQJYQVqIn8PASZjhK/FJz6KN/zL5Uq6GzuWG/qLQkMkQwor1LR6OpH+5p6G8
s40AAQqabJwnBhtT31hYaFobHp7RMub8ar3sEOHLGcODNSgO4GG+Iltr4GAIK8d0
edMd2em+8mXOoTRb8ZrgUddRDedfIo8/BBgorh4yWc05x3Gj3Fdfcigaw6MhL7fN
rZc+yMYNSz7kuUYOe7sdEWs+KK7DCIf2b/HuG/qjUab+yI3n0r/VZQeZ/j/UhO/d
wH+JbAIWp/xNtCsIYEK9nplcKWKJ+FfJPUgykNuRXFoIY71vAb8m69QXc0dYg8Zx
zCV3fPANs4E6WUhbcva4SHZPB8w1Q69np7xVhjCWgw4T4iuw+RF6KDpe8oWDJ3jF
uW9KuOo9lxVwdiSZq4SymDzC9aOFkeKCuQ8Q2+k+J9fSHJyusvra6Pjn6ClRmEzN
S4vbGPLUDUg1MxEtV8vwT0TX5NxZ1Pda1qHpiIRQA5AhWYZJz/MHtczfR9MoSaHC
+Ltxb5m2lnvudav7UDhtE7+ao1arBqX0eouLpq/CIYHK9SYRfpk3eB1VTn+tZ2iR
WG/8fVvjp73ZYourVVlqA6Ey71lnBSlGtlZhaApDDKHnVMTK4vmXYWk3qnu+BVR9
kLlh9m2XNVTQWrF2syi9yoxOvjyxkEUXOedDNsOszrXuT0YUjGBAyaw+XybeWXRt
fEK15QEuRt6Dm0tR8+et6a43Jq9FOTmRASpIlufOctJ9cxUs7oOH1h7JSn+HRGPk
MibI3rlfZwGJDJdr/T27Pk/t1gk+htbEHJVR4953ZxYesMPF/HS9Xwl4mUXvNcpT
y7o0luCs9+xLZngae1ycOi8/fhycfzeA4hYckkkgAuJrdbye5HaekYiDr7OHhLCV
AGKRP3ZcZycQCrfiFVor78rajOhfgvyYgDeIrVPdZog4Zsi0egYZbbt2PGI1xr0b
V1A4MPEwNpHOl3o2Y0eOY2xHsuaA6KAGZ0w/nagh1qr12mIJH7QLkoZtkTfpaQRI
BqQS2Qe3g/ScrtyWmOVgYy3fPmga4D+3HmCi+5bsSLZV2ZPSLcgGar03IaHmsFFb
TOiX4ncmfViPhCUvgxs0Cw7X1Ch95HbvIA1WNHKTuoaHumYRCy2zbW9h9XC9YfyM
+hgzZv+18I91CMKxqkFxEvmIxQf8kAP1iQVYMEUqhfXkQHI7GD016HZ82PhMtHi/
H95EI7sFQf4vl1V0eHAznHXCc08dgnyYt+w+Cgg8p+pxcHzfeoEvAfVFL4ToftFT
EY+2E+PqL09X9YOuaF4gKEnuSRScaul058pj8to6OjSyy+qVs63t2Pnfda2U5CPK
Xn8A0RaS392updxir35p8AA1cW9sMJ6hQ+hSEdLmrC5yLBEvrll7O5s2w9/Uwrwd
SUNeDa1qCAlM+ddNu5Q+rjdXkT4tgI7vbvia+fZP4LxFQZu23EdB6LROY6r05NH+
8R/+d3XcU4L6ZpflQnlrYzNvxPYgl2Jm+YNGM8Qphfwbfs2RM4qSJ/WU158GHEZf
FMkigfBHfzmdIvvUVQnaXZ3dKmtgIJEbUiLiBljZFWipeQMJp0+gfNIqOOtrl42P
2hVxCcg5AIgHFuyvyfIOmOwzytD64aj7oXrZmPzUvHfoBCp0WCmvHJnkbMobx0hl
E2VKrhNLubHdU2pzAAuHPbMIuKacC5ohJ4xKpRwpMAE/2Pydpy/CiVQmySyATSeL
4olltMekwr2IP6O1Mnjy2HAyOzHh+68Zjev2QMWf1ES0GCpTBIx9RTyELv1J6r3D
YYK6D3F8pIyhFCU4tz6iv44cQYVdjRhhJO+c/WjEHrblTT4MWGgx7wzVGTpAm5i+
+vqCzrM76IkHYqlaYpepYlhQ5zvoSLj9pZlus9XSYYcLSbAAXIoOJLZmBuZ0YrPd
XhhaINXlYd+5wvZv4SWt5e8Bg+MQvQ8gRGuRkzdnTEkzfJ9vBybc+qfRYTT5NZUe
+tjtNtlcmJRkCKeC2FpeRrvE7dmSvcEQh32g08RT6iH+jVfU5zNa6Np/fOHFMV4U
pDs/tL485I0EtysCwo8KiN3VPWURdfWIGvanEGsgap9Np6Phv0uPcAVcUZELRrCo
CK8g+kFWbHD5vLrhNc3edk00dlyvWNkOhn8A5qLCrRgaPsErQa7sixWizVMPHtjV
+sdULScWJBiyTHUQCOQY6Wzp3PyDpdDtX5X9iz1CngtbBARiXdHmm3MK40VYA/Jl
IcMgg+vsXgLmyvhAcLtsKrEKbWiRQ96PYj3llDr3AYRwNVgWcRfJV+tP/EMoM8Sv
ebUfE+eZJnX6Zg49F2Ue5kW3C/nMEARUH2+avL0etKwFgNYcYWf8AnpqpwgmhhX0
/TfFim7YruNLruw3bTw7Q6GBEQNQNiOGKloyW1NpoC+ht/GvGnvcfvT01WUuaJIf
aJzMJ2OZgWOeOZz7ekHoLl5aq5ZjezAeBUjG91Ts0k34fwzxLOitV4CFJUyE6WEu
R+fSJCqsUq5QUeonUF7RSaUVX+IXjNIkcw/6HZ2cZzx1jVgMK/a6V94VoEH7ARDt
RLy9G9ZjaEmol6mRQhmxNIOcEjCj/wHMWLStklzdqbiQCakHeTPT9DT2PbogWwAu
0Bh6YwZuYWDNzTBbIUhgrjO3p09e077lJD3BY/nIMs663h65HIRX4ecahkzBU3pJ
zvrZ8qO8Ka68NkuNpfmgmGa3YJ0IjXX6OkpSycp9zklgJ1ryxW5F4M+hTc7MdFg0
Oh9dJ+EhK7jBhRyU3nvWanC80l8++8PaBndGodd39339ZiidvxhXaOWYBg9Cnxzp
h86GAhXCz/QlYOUvvYb2UZ5aE8wiL7oEfUj1ajqrFFIB4Eg1Ci9+htTdGWV5G9+0
knGkVd18oKqYJ7ZxFJ6serUmyR8hP9BF6/hanYHi2o8p0LuFVbI7e5fl9doPxRpi
cI9yy7FXPSFAINuRRHvhTAuuwQ25p9C+9jBtEszdCa1ljAljHD7YEqRLvqPAVY+F
emDWnyJqDGx/qbsybMG2pIf+SJIXglQCg9ea158si7j0xBjOPsbuvETZNfEb570G
39tNOmZiYvKzc1YRdV7s9yxPLeIzu2U1LWHBYThgc57UjiVJMKDO3xvs8xsT3erS
z3dmYFiu6i8lEbrzEsN9xfRG03jEXC/6iZhdwjDJ7iEwovOi7MlwiNvg6WEZtPMc
VOO4pser2KcDbAoCvGvt7Z/DRl8XNSlGiSv9IB0r1/44kX7ITd+BRSEaGqOW17SW
rdr9KRUxtzZumcijmu9DXSYrShsIwQ//n2kmUmSsFgpnrwi4ylXOa1TZac8HaWM1
qAXPQlgbLdS3G5ykvGhmf5n6uXbUKJtpiBqycyDo/CjwmNhK36ScRenDeuH/18cL
pjMg74lT2PnkdcxEoE+yz927A/kqr0r28YDPm5deHvu4z+BZ34AnYogV1WRSr3SN
PeN3PuLXowbGAv1q8E2b9zDsRlDdn/p4d6agsRj9gIEcuIWVocrBjs2mpy+uOomv
CbBXlfmHspj0E59kxBpSNZZPXduTjo3hWEb9c4KQ3x3pagBvrD0xsdmMz8k1N9go
X9suRMBvTUPK+hhHni7scU6TWMOlB9Z/7xmXyswfAC2H7xUJxYm5GTn1FV20pc0b
O2Yb9wYX1Gto291AniQJ8io9CaqllBPmAg365oeqakSFHCosmQ1zljcVt9KnwIQI
fd6iffeaehtVqO4GJsZ8KVHhYIF0zOamDt0bveVyiAdYSSb2vsu9pTk7Z1WFerpN
Rj7BQ5plXu/Oun8D48XqTqHffggPHUtPWMNzIuqmB0j7PBPaW3mmbLf1vC29JU7K
nmotN1LP+qlAbSXys5EjOTXsZPfW8O7LkqfoORSvyB/Y3ueK6fZ+TAr5XxXFAmok
+fvCOeUWF/ysH3RWMSir4ua5R5fpMYz0ms4YU6nOgKxjDvxv+vgABDGoa3omVpgE
+ZynMGu8+ITHoruca5WLZw8vqdyyM1DQVh8vgiLXkprTdFXMd0pY5jN7rW0wWlkR
dlTQBs48bhYO5jdyVt5SVtyJT+mBMO6zWwraWq479lS9sJMUOda34/2hMYD3vAYO
jP/D01sFP6NuLz9SACpAZqbQ+TISBaka/DhcUjSkec4esllEnIZir4NQerFgxzbH
w94b/oGMjK/TjQG3apPkOXRbDzjzA6XJ/WKAwZfWoi69On5HJx1h5Q+LSfFPFySE
M+qUbGEY/XPLOtZJ1nFrytApqxf0ExgRG4gecFHwWfF6FfZmSS9mUFFH9wZ+iy4C
Fz8yYT698EmnWw5n34T7SJZ/G48LzAoRI2zmWCynT2R9wlBULxFtn59eo+K++0uA
SJBHaLj/iNVxl+uFDvTBgj5aIwRF0miCCR0odXFUUAx5fA22aUv1TeyiLWt+/oem
KW0c3fwZBkyKtsT+a6YAYhAvBgMYb2XSvrfc/WOgR1ASUimnli+3ibEaxVEkb70P
eZXB7g+GTmi+z+BVh/VzTnXU6UT9vg4m9I5UVg2OMfZZF7DihD+oe98eahHdDzyG
KGTD9mo+61K8v1+gdSORZzWcem+gGWTLtlRfXcs62B7SjQlLllQ+XvewhOkmL3EB
nTIOWsriy43CmBD2ItPjsGCQNcYd6waoxNsPI0s/LUjsUMNwsLroPFr0AVZfZKBp
joDA6w4qmVx0UPiGLFrXCbfXe8Sw2+s9M6PCMOy7yzEJuIBiSGn6yBiOQZIld38J
yqXy2NUVZvNPiXhH2lInSDDX/lUTadJwwSC2SD4lzmYEZw2npBksPxaOzu0CWDoB
nDwIn41X5khZIApQypU2CbZAsPxeq0kDoftxlZzn1YXz46ezbdmskzaey0rwVcGc
uQjAe5J8TGtakLSFgssVWUjZEXSwoB9irGelXw91DuCDgj4U8iP8010TIsY4mDr4
gHMXOXjBUvytPkMp7Soqp4LZvQXm7XFhtEQ7BNK6QS3ghdVlF7zX0uZFJWED9fbD
k88C3hfEJFnSZqgIa0U5xx1o9OYzs45wCxAd5qLMAkjZB5CIWJOYmOGR3PBnim9z
HTLpdasdUnx+obyG6xCFRaaWDG0M5IoKIpKSrEtnilQD/mXG5+d2GNM5B4/seCJ8
`protect END_PROTECTED
