`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vJGLBy7Ap2lty/9nvkHo9nVo3JB82G+ByoNyG+lJNtYk0mmEXdO76evDJ3xvE2pv
D9TOPXn05YIzUdMu7WjfbWWW+165PcFWUOWdGQUehzrymX5/Pc8FVac2V0UCZT1E
BV2ujbvX1dy0y2GcYAtMzlhHfa7U/UrnLJLQD8ROhjmgeToEsbzsJA84/7QsUKmw
sqlJYzCv3O7scq9ziFowZr4tAvNsrGY2Injx9B9c3k9tfYznqjxgBsQZyxMPFgWJ
ssD2F2TeMHpNXJSwu8WihIupzOtF9dWef9QcMKT2ll85XtGjeKcTMjORc54PlWgV
u36buwCv9sWPgpAmK1koJICSJemZep+paz2EwssxJNvSLViqh+mWUDZlXBvULlrl
TCZ/d+7Asrh2v8uNlNLJsBlD0ictH21p6HIVOrNtZhEtf4MiLFlzo9bzSoQJu3lx
p0cUBS2qv0T0xzadoRr18BJ0MQ+RD8ARzxSte8yAeo+bBP/x4VMZ5Bd8HD6hsyS/
o8/SKKJ0rky2X17hmKgNvjKf1A0aDWa2dfTPVjj9S0sW+A1Bhv0t4v6Lk+T7J29H
5a+2nXP8e7ozkUKovdoWrF9WyJu538jV5it+5d0aMAAggQmsZEY/Ax7NTt0hl6Qk
Ub/uNq6qEDXmUpTVC2eGMT8YsQ/KIOsYCz/Jt1dqCdr65RFGHw9MnRJsYeV71Rch
bykuqZ7ED/2LGlXGethbtPoUzRxpfNWrtphLQML5xi+KXsEYX4JOJstRRv+zIxEf
wC1jR8jIyxNYIzUCrQhyJh/pgRfAARwCxCJ+2dhXZPcdm2oz1Yoe6Z1T0iUQqyhd
+qQn1ZJzUn0WdW9N/U6sdMoW3rFjMYewRJXO5gDnv/5jQC09nLpsE/pDYuk0tzkz
/UmjmsvzKf725uj7v6Zsme72543UER7SKnRffMlEaUikwJ3Wzu6Y6GAgXxeTCEIF
qLBfkD70Vo9ZfRTpqATxcxT4Iqv4UIiOy0BbQCM3SPBjCEuCf7EVmm+2xPFSz8Ww
88HR56YL20ZNIKMoGN0inPHJho4sLfpfOlGgOvFd8rPhO9NZsU08cTAOcIMEzAgY
rvuzjzr3Cb7WcHC1v75PAcfQ+auZFnrb52sJaexor9i+PXSYsvQVvkenD/UtQFmA
nkYyFcv2H59tF75WH4TmdqVSvS63FkUDIsvsGzEMOX05vXwMdUO5jwe0vSEPFkT4
af7GEP8Its5fq7FCGpmlLil1zRI0JDwVweyevergu3fdc42UyCTrbWqa7zORXOua
ULUUGwr4ZPHVbUdMNjzFsckhvw/dy73ov3cChhrl1P9vroL/DcH+wEeBzDM+4Wgv
v6njln3i2g1+DwQU+ypcJpF/ikQ47ry+CS4m65Kqj37ehx3VvudsDjZGvGUsPkUO
y3wUE6D7bcqWMdLmOloq+pePEB8mSkcWpyiwCa67j7Nz4iq9v/Tj2iD2mAvUYp2q
G+XIw5jz6s4nVih/IPzlNdgZLAYoNatv8ZsVyybM0sn9QsA5EtGEF27UCDpHXxy+
8W7UG3ey/U3j6fyzeasPahUV2AGr32hVMGBnCrROltRTuBSCAr0aLmxDp9NuFKAa
1trHtPFjp0t1uWv5edCI5woUapPyZVrFaH4kh3AnRKIzws54CYg5JK9xyWOwX4Ht
ZOqzjeFLwA5TQQBsWQbcDJk4L8IDN2YHxypcO+g5O+5QUfx5XZcnb9kJbmTYu9eA
zNhiu7j9tgp6nOrnLt5nVVA6HZSqeW/pjUDtkPvHtlbQ1XLlyXCheFVaMqnX9u3n
9HoplaIYucuqs/m5nsDr59WEqRU8G9Nif9rG6HIuFWxTgeAhimwKcphUNQujqib+
DsKq4LtPOlyvX9YenzxlZn1jPVh1I4kS8w+R8CN+4UoQUscvK6F3SvkzGb89ZkZ9
dO8H3SFelFCvskXoS9mDe+zPutb4exO/LXrA1bvaU2I/V28Dgu95TvKWwhimtrHC
28I/F2GIvtn2/x15KSHFMjJg0ouVGbK83xPXE8+kWRWTibMEK0NjI1Kmj+m30XDk
bcZ+u8llTFaVbhz3aWANjpOsHemWJfXQcd5CxhB5rpYOxvIPEydb5eCpIHr6aUg2
oJvo9l4Hpg1baKBASBf2O5FpRO0w6n6aWPFaany3aA+rDGyYSimVjO4Dww8dgIqI
ShRzkNhfb3NB3GY+8Ayv0DR2mRMffGqEMnUj0aTtn8SRmEX7cQRD78ICDPkSOh5g
2H6RU4PPU9kQa+QLDMDKt97B4B2OJiBYfYCjI4YSqSZUvS8WuR2bOhL24B++L4dL
F7TvlzJ2IjjmAqCuOzs8AmHrZ/uU/+6L7B2WH0YNfTeFViRR82k0IEYGHTccOLkH
EEqaangLFwsnEratdbNvS3xmVSp8ATwhCBCxxP49OFIHw8NbxYT21ggg7Tch8zgp
tzYJloM1CAyF8U/hzjAqLxUZJma1jUwnd0KOkt+t6GZQQ25vN7IhNmtVThNBP7GU
RX576qVMn+v5vXFOGCwj8RRy5efIVaJZk2aBfkqkNlMqMDYSe9PUVTJnybavh42W
PJwgf8Sfz9FwJ1zcZUaY2IhRv2965wT2ecHV91XfFD3bPRSHKgTedyjBbE2sG7hQ
rQiLLMH2BuC5xGLWQDuL6zN+vq3OTsCEiWGEzkzooyvx24U5/RJpIdq3sZKRiBcM
muo1Zr7XED/UJyRgFT2rhjeATyd0qOkF0CH2sUf1gUp4l/xsBkJ/gTr0trtHzSHU
d7rqnRktsnke3EsGPgDSERaz+NFeEUMJytl6f+t99gAFTh3Aek//z+pzWcSEUdd2
pN6ByILn0MuPBHaE5OhhGYuVvBjAJEKBcFBIN3TdC5SXVf8Txfq7vEFPLYpameIs
e/+tP+RaqRz0SrNL7iZ5bBR0Ij/Iq7UPQDPFUkVM1GDJJZRws6c8pNSFdnr07hfn
ABCli/772I3OgReR2Rrn5R5RaUqecMui8NhMEWW0sOphmplSxXLTRgUVuE+l/88t
hSNSY3j9i19cXhau2JjM/wl3Dz8jYxVL6BsFwBjxN1/acam2AF8dGu4ggBsYNqo5
7rjRa2ndnJZS0+sAzYt1Qpe+0Eut8g6dAVo+iTCWNW6DWUPuJfgAAwtdbQRPrSMa
o8Ml92MERriWXBDCh566nmT+Q1iNudyRRo4ytFCT1x6hUxEG/oBJNw6Yx37N7MTm
/Zf64hUD4fEz6mSa+i1R6rQTopLAnb5C48BpQyNCfgNelSU0YiW+77nIV7600oET
Wo5rObNh+ZfbHOgeKXJoKVzeQARmwfQQx5MjaxUL6TNQwh4pSbIXyNllxTrBhvyo
PG3a/zMA38PvOm4fcCCKNb74WCsmC9gWWErM6awXO1sRd6LgqHhh9a6bku2kdCVg
OmKp6x6D6E00zesexRvRSmJOLCLcZeRTJXC/bBeGOLGauSbwPPICYmvt5GqiVOwy
9MvPPrrJWm/wyo/bS0MeJHn/TkQCa6O7IUKDnc2xNofFd4Usc4j1U27pqUkxX527
wQtnZ0IStCcr7GGik/3bNBM+xgs6KVvXEFjz6LlYqD4h9AhRJAy1nZn/wrgpj385
uAWqiDIs1NmyXtWam2wK3gIQE8xt1no7xKN6JVnWhQSMRKCPTPd8PI7yiVqeq2TM
yhrvroLJfHT20SyWzajo8BKrMf82peU2NEHUd3esr8H89/Ufqqv+9cjFeoTgDBRY
v6S+Fb5wus7f0G8NSY/kjfUfQ9DIwpUUDriWII446YyqKF5iV1zktQWeDP4IJ7m1
OGhaaAQUqj4zMRECo9T95ADFLEoWmirYWcUwFB1xbeTmZwuJpCaqpdbz1EnEU3YR
12in8/u562CpTwUZzUAox/rMY0Mk9m/qzFC/40kK+B5hnrNBsgEYAE6QzH+6oRM8
VkXk062PdY+RWDqzHLigBQPGalG9cFux9b3omXBh88pTS5puc4yigXcNmHk4vbQ3
y/tPHLJ30pYFj+1m1z/XJttUCw922KSZJla0jnh5Sd2Mt2O/chxvdRVut6jB3tYQ
O7KYVMSYr+au4Sm7EIhit60OmV3b7w2b+blbf4o9l1/2jf2EZJrWZjTgxG/tn2JQ
W/61kIEIdLzcoCrK1jTSkKNmx4Ut1tXXX3p1XMHTVHcmJHkqEZM1DZM/6UyKGhAo
EsYTUEP+vnL1bbuYCNiq25twWL8n+kEjd/F0d1dx3sbRFeSyV3nXIsiI1/R1FTiZ
9bGK/5qbT/2ya0s1XJjmxXOLw4Vp1PPZ87YBGwo486rflF+JAd+dgz50BDCS27SZ
FFnUlFOYnG1612FWJHrWwc1/hATM4gaaOJP4zYt4XkhMO3vqtbXLBVHaM67WuXo6
oBGTMuSShuyZdqY+BIqwttShDnXRV5VimOgcJ2RvgLkUmt69ntbbeMwe9oRGstRF
R17uEQh5IvUNVfHO1Aac4qaf54qQUX31vTMgG2NogXHck0JqydVqGOR5/eOp82aR
+Vg9Fw8uSQ3LMQzI8Oud3CyLX8+O15QsS1wUUP/2ZYpOAH5LjlRGC0lDBv2svyHF
bunvOtjK+SF+Zm2g5BRZXspQtsfXtA3c5rprCYOIV1p1snHzTLeqeZ8nigryqJpe
YWtpRupJ5i0bZO/oQJa3sotNBgg3Njlfi0z9S+oQU1QafRnTnZivYpkvvwm6pjxq
abrZiQqx2DGuT00eztDxuH44DjOwHEfoZXePBdEYIxCbMsSoxPo3c72INEvQSW0Z
NFresdFZZe2cMihd9iQx8u8Znwdb0TyKI6K79DCQ3ORtm4WNJJZ4xZS1BvkWGjuz
NS9g8SRCJNkHxTx6JawIZt/HBqIkVY+9pkSirh0fvGGn1CPrc5ULGpCnquprf58O
f3QhVAifIGUwqgDuSAxpIwLSY16L7FW0HoN05tiH9aLwdhc+g77ZFMPfflRsJXtI
XgDuXowtxkuIpNpv8fqxU8CrcKAG7ZZmWE+kvQVAbSDet3LUZeKcEpekN8eQJ4nj
ZPMOmCNl2R9gGwpsp+vw41yw5/C/2oddVOhqbwQixenbLm5qEIY6MvUmjqEAa4lB
aj+mi3RVYVAt0D+X2VOJQClcAJei9WWrx1PIKzi/kgMoXLn6AXupTFg1dF8CyCPq
IYlAgxndmp+BaLMenlSUl0rc/oy64RE1TVz074h06bGMSo79Hb5Z8u8sxZGVuMBe
iNpGK1JDpLuL1I+oY4YZ16OSR8vhxJhHg/flqoyAr1nXrhb+jKoWY0NqfpEVwkEv
P20/94gSMCKWxbLbs+trqesm+snBxYAlaUh+dhVz7qPBQBt5DEZxBnAZqkior8jI
xFG8QzewZkfvbL4tWdBJKmN8U3GjUEX0gpJH5VkmYWAtoiRSNWYkEg0QkYPoNWWA
JLr+7YiwcyPUvZngkD501qnl/vNPr22wriK8nqPreGxSWI+81GAFZjWxefGjp33y
ZyydI5NcxLz6zfV1om7bg/QylBjX9PUXXNsG8JpMAeil44ighVbX8Mtnh5gqKfH/
AmIc3vRo3tGYzHUaX3pZvukroClu/ZO0ZTMOC6qlVLNZgrRbla4aCPtTL8TDqxwv
CqVUOV+mFbTWej4XxitgH4V4t/tZLQ85rtJbxZ5gSS+7LoUHrIpCbqRZwXbmLuGS
IuKK/Z5Hr3S78TYdtOliQC/KoMAfpe0cnVlRYgTxITVktxuCa5HRIJeJo6JHt1GR
q7ntQNvXzD7aGjIxeukMCcUtMQBL2p47aSog0b47tiVOSnPsPo1cEXdUP0cBjptG
tDGZRKbTxNRnhwGfIOO3tQ6IP4YDUbl6u2VD1FZqCUc4Ylsh+yyAM3Iw63tj5PSW
nnKu/A22BmcrVa+agnz8T03+uaXnzZIsibxhX7OzkTUYQ7/kqik/uWhvq6SM7l1e
0pBRFUdA0GzLAkE7P4uxfygZ376ONEnGATGDeupKHNSdNj08pmR/1WucqVZP4IaJ
lPEba8H7dxBAX928iyJKEMnuKGF5O+xjJAeDGlj9YidJd1pP30DJeu3aOL0iU1bh
Q4LdgbElkjvB9IMHnT2mEbhtIZ20KLN1a9vIuab2XmgF1WeHOv+lRp4PBQFf4eLN
aoyUsnfXl4Bp1ZdSpgVxU/uWETzGzPN5KphyuXXOwg9g9Ai/fN4qC8SUJqY66eGq
a5inest0i6pp/UO5Ci3sshiJur+RuAIBhAzALNvJRT/zxblqSXBDDidXH62t/pAJ
NbvI7X0Sgjm2yAc/ohvYkHf1SIGr95nVuh6rSCeniBCrOJKjjI3A0YXBl3Xc7UKf
Gf/kFF6OxqWuTciCtWuy7CmV0kn1rmDIsB2vBppHD/+U4V/0d4QccFRglap+nd2p
jhBmXWyKE6lei0JSi2vM6AZ0GMJnCUnTinlO9YyCuckbHo6pmh9AWUJD9EOHLx/g
ZMV1GGPASSzA2dKIUKjraS84EVY6E4v/Lmn4LwYjQoSe58AmxcI8jFJd/VUuUDXr
juj53+Qa4FZ/kTqqDljCqwni1thdxu1q4jXgccq218NE4o7DXm8hsorQkcXc3sWZ
sj7cjaKT4Ta60sQj3UDqWoTZGrpTJhiLskJ0SxLYrhpxifHzevNFYGoyY/FmdwgN
UEsTd5GpN7YpE69NjUphie8hVjfH6ZW/FOuVOLc7kHshVNPF6KcSVMtQhx0sa0Rz
BLephmPr204AyJUbdvOy7P2gwrRRlYpa64k8Rp7+D96DZ20uHqd+haqVms3VGfSq
daV9ccWmV2a5VXgzA5E4pCoeyu7FtAI9i5WdksEb4SYgpU6yIb8mq/1lDwycKNVN
UFDQZugZ0K4Ti2XXRo2Wznc5nHts8pX1uarRLEt/Cmd4QBPSHi+5Fu66sOdXtRBt
1NkmlFUj8+fsdejImf3CNjs9YJ4d3ZY+pigAQS2ZtMuC/MEq0uadcEdbtjOGbe8x
aVs30i692hh9gGMBzijJkavvnxExLfmZakvYiXfJhKLGDvlKh+ujJaUToduVa5L8
yYNHD/woP1ptOy01i9do5CxzaLkAsz5dHMtzQaTMtQu8fcAKUd5uIDQ+1rXAftVx
LgfxwBeHcheeyAxeMEQRPbdr1VQWoTTMDq/wrqmCvTutga+fEas2WDOPTz9EGEE8
RalqhD0TcGu8rKzh7G7ce7vlgPChbnccoDgWOd3zrrMcpxREW9JbWC4La/bCxU3J
g7+yG01YwoK0ziHjXt1gGRP1C5fS4caN+6gLo1yt9K78YRXoA7V//H6YgMuung9x
DufE0rVLMzEhzfYlj0kQEqa66u0d6gSHGgtzd8cK5skuW2o+ML3yQXGyUvkO7axx
dAFwTgeQKnxGOiX646WQ4Bbf/yjvf2eI17S43YUES8lAJvOv7N6WiSwc7GrX5fEG
NSgL0MQNdTh8pKqKdxd7awUvxF8O/LWKfaCjnvKtMBMocoapJEj3ragdB9j4F3wl
xRkv09VtkoRxeSbV5eXP5BQUHrPIMZUDARQCAhw2U5Q+6YQ8HJ2eqAoeTP7n88Q9
ml+Q0QxsQQOsLB6bWJ6Accg4wXY5wP3BmceTKVsdOTiiqXuRESOEqsJVoZqCrRZv
WbwK2xVA1MTN92ZXqPcXxg==
`protect END_PROTECTED
