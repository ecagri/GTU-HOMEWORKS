`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0kJQa3EoLGsamMIAR4TBN07OJx60R9uJWBvXsyCLjMpRg3xo661HI1vYbcd2DdPs
eOcz6bY8Bq73qo/s4CV1ZbIUWWrByIriQfGcy6Sdkm8CVADJiCt5OnV2mfsZH3pc
XMKMvFq7mZJW+Gjs3Bgg0DVp8y07gGj1y3W5qcRz5BA2TTbUo+kED4UuaZGrsaV1
clT4JhUV5xIILZeTBOASDC6ZMsprzaxEZDjLQNwAlCDaiyhEQAn7wbG8QBHjQnVP
LCrGnu9yHyD18seVPfRNdsDrIlsIpT7Ws4fekM64jKByD5xB5uq/t0wxSURwxFor
kh+xj4s0eDe11NtkVDt9xG6kabcYHjOEovnybpt8xFbR7o+fXwm3VIXnqTtHl8AM
p8xcTzK7RqEAgipFQ4h/u67hhPQMuvttXAx6ew3Zc7NnbRB7x9RVaajRTuCX0QLy
gj9kCI1sIWLUWeAZBDjYz3qtKwaK7srD7k0osoRxGFtlka+cDROyxZMgHUdNXN6D
sm4M2ulh+d8cfKCzzKWmZACwkma73LjB16qAX/0ONYa2/MNAXYQKYX35MafwQz9J
5uPnDZ5LalTfWtbAW/jk9bt7O8NtdzIs2Xs1ej6asmkwAN4BeFm0L9AYNODaMZu3
oj18Yplizd5hhrrFisV0uejcKcUGcTpniE3mXkmGR8W7fo1M9GQ9MqhJdF+7VoQQ
vdP15H+Kh+d4XSsz59E7QiYpqAXY3rM+d8XCAfMv2y5RtPYiYXPmiIvcyNuLBjMS
RIAR+tIzX81/ohU7SngP7qIkmd8vI60u5Q05q82DXQD+VWn7EeVp9lQVz/DQovBR
5U0vj+sYbsdwMKfvS10APUyisxA9+VZA3RBoQAWL1N5Kiz2CPgm6Z0KN5JmQymoQ
chgyLv2YdV7PEnmYlldU49blASmKXAGLbO0j1BOs5seFCBcRgARrJubuVD3/FLxz
kJU04TkYxSyXiow6iE+M7JBe98TFXsQI0z6a+Yo4iMhfs69iIzdbUO3GPxWAv7q8
J/0MQDGtV6YCN0ieAyRQicdyavUGPCsy4t/WBud186k/lKbEMXqzToMnKeYABhRY
`protect END_PROTECTED
