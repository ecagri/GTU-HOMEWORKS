`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zHQmOqN67vrex9WRbjPdR7M8U+9w1aHqRucutPSxeKZJa9wIcKYg9e6p2A+N2JWY
cuH/K+s2BKIbDqJg0CaTLYcoFgr56zGWmmMXg855fM0UBI/q2D4UyMbV+Q0Pdw4N
LyA94dXwL6w5UdPEmUFttgAiNIzKaLK88Sn/NfiHLy0lIKXBDUuAugSU3Lri8B6d
Xf9EeoAm12GI9tGthI2HR9GIDnpXGSXKQI+XPnLCRljV7zBPJyKgsTSU7ykKAg0V
kUND9XzB39sf47EyrVVH6lnMYICmwPclm2/cOHg4sA5D/FrY75Pk35FJelLmnf56
zWV0fcnlAQ9IH2azfGxarvZj3S0QM7Q7kRY9HH8zZafIEZ95S2qE5TmTZEbAGz2N
9nSbdNWXtxtshm8lAp5wtBFOCV8ZmMIRbDfuNDG0LX6KmjR00hxCam2jGhqHQCA3
jhXVW95d/5qz4Svvkfj0qHs3GMdA2MCTdqmdkVQTZ0wgl8TfXuNtObazyGCD6n9L
4urpBA9OKPCRxIyTXi03R0pg9ilp6zssfscZsM+2k92sglxerulKavPtEzodtlOU
FbqS6JeN3cRdfx5fxItvTGkQIc3btFMp9SBVcLEXibggddan7ET8HWdvcFdW23wY
S7xaAbgAgce9uH8j0vq4r6XOZmjXz8DVnTe6HM0tXNvkpJlISIB0zUweDAGb2eDy
noRA80vX5wWTXXpBpWnrMSuSwqd+/TYicFpJEetqixcxxYnp9Je1WhN1nbtDSUY2
jtJjsZq3k5w5WKsaeNvFDY5Sp6gidyzSg0UCqzPjLUGOCqFO2etENPkwU5560i7/
4VyKIt1QvMhr6XZFOMKBPlXiTVnXq2g98WitexJjtcw2JUEhKRKrWomqRZoIVosx
aBwHW+0MJN2ug3KFKSgPYiGBqEKjFVJvFABeEWQpaWW+19mwSbNqeeDKYKb83bBN
nOKqv+llzRUFWfzwGmihBgnta95XUCAOL0Hu8fcwTKigBXNzujlqwmpSYE5c5hUr
fRAaUpAJZy5+nHx0vA3fW2IqUiBthmT48EUTorrwXpW0yPd01QCfOO7spcz5HtaI
ZIV4PgHMkMW2ijE56IX1PcGvIhRSZ2Tu5M3DBcyPxQS+HGAXutHfL0IW5YeokCw9
kAhPLNHNp+QPlJrpUGmD9Q==
`protect END_PROTECTED
