`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kKYWvMxTiscmkkZTT3UGyF+nV1hc7x7b9VyeW+BYzgEvFKCe22Bprj7DFP9ZGHzb
KFiwjVKs70IurPYUR7NJelhzCWgVmvyZpRgM0Qt6hin1hgvY6KpjSW4AggDE5emb
mJKXcfgbooM+VoezeA3RysrBAinM85sUmi8gikWl37q8l1zmtrw1TnzNJbQNKuy8
mQ/w7RIV8Xmu3xYkxiHewLsY8JyTrkfIAvMFn7BfISiy6PDuwNC3EqtQE3Hr8NDs
LXD1Af2/ASulnz8K4roqUSqwuH+Pb57LmRlsQ/LyvpbnlEek3ihq0Z/JE0RSqX5p
/voUIblWusk5H3n+N+z7H9jPzRjF4UdNgT9gSe8ghFNv8xqsEu4v/gT2iXq31yjG
PDAtG0GV9elvxCvnXvzRFpHX46zz3OGQfuf/c/qKRXTSXI7R9BX3NR2EceZSjunb
xNZzXE56eW0loza+pcl7M4f7w2X1I+gZ70TuwLSK1TFIrPtp6fD2hk1JYdQLPZfg
Y/kzC+h5Zy7jzcdLTCpuRGitej0dGleCVB0a0hliKIsZXWt2VKkTrMTZfPlsMeCh
ESKurinWxXZlSu6Pm4w0tzrgFFeaddjTa7bdY4DLIjsAI4I67P99rieJzf9uK73H
5JJHGXNtNpAJQZec2IuNXdVBsv+zaqg2YOIgIwzo7PueaFzOLSgHUcUpmyHr/gpJ
zz5uQn0An7klu9tEp2tZUZXtL+Pl0x/cqi9tA6VlM4NtcTeFAU2r+uN94wX/mLwN
LcCoBEAnfJEXl/yeWDKT18VVqL9GY1X1gA7FT7LjY2ljgMUZspEHocqA+BNGtG0W
5jHaHtLV1OzuZwpEnZC+a+URu4wYyQAb/kaaVTbcGgTRi8mY7mMEJMbKSRy+7ccI
rxmCEFDAYC4LAmzMvediBU6atee9WLl+V7wLtP68FFkMbAUs9JdP1wdHcRoC4JmF
3Oe1c956coHQmFIbhYKMDejYZS5FiSJm/gbyKhvc1Eh9O9sc4U2lgaz2QMn1MIYC
3G9tArX5nutqEso7JBvrnAfzvJ/t2E61oFWLIQDhNj7dZLI9dhe2ksCb9IQ/xecl
zbJje22Sx6YsalOGUkQfm0IEfejNrYIFn6JBDkOKUi6h8hdiW0ulMMdeCKW+ABtT
FWDqMSTV+dwvNsUDpQoTpaKzlaHP+KNGHovtaJxjZSsDTxhVway/3EMVp1dD0RbZ
cIGvqOzzIN+jFD67GDlpDXzhcdEmT3bms7JuGLLmXn2znAifGchoTEQYtzapL/af
yET27NcgXu7KrdijyCoJw3i7oK7HB/rJYc28WadriFTlUijkpi34xsc0zo0fAMZj
BuCNpJGMocQ44rXD8pT7aFYlZRIQwT8fsnQC15CPB3kVKuyteREyzIfiotgpZUyq
yUO7cfJ4tJ0PPKcDURjgLZ1unYnEymkfmDhW949w7+FfVqmN14JZliDTBToeH1Nj
H0fvTyk8p2yciInTnrTM13CDIwwVjaN1bpWbq0aXtOnUFyzc1tXldxltw4+dfXBc
A/W36rd2wfHj8KvC+Clq/MQt1Jep1ZVXDpOjRm78zHgoKzVnOgu/OtNGOVnjnGo/
FV+2xAslWICh9CZk9k86CQI8SvkrjqJMWcqhxjkRrDwWaTgHDzyuLcjhgKUCr4mN
71IaW6Bd/5SlUkMGx3+e5Hc2hi/19/ZoLij5f2wjq8EddlfDFJheFAAJ3LpSWX/R
EPW8PIfa6VrUoexnIvlIUithVfJkX+8dalWoAkkb9U0O5YYnkdG6vIDbLo5HFoOi
m8x94BmVF2RW48oMHVFOpga1n0+vVRt25/BuuP9La0T/wDbgkWQ7tSZ540bf9nsB
DYf9onW+zHKq8jL1ch6qenXNl0jB43nYda+PdL4mlr+h/Wi6svi5ilKE41v0RLCa
sJxdk5kB951lcKxxHoPgLemhS6sVTxtuGFONkMcgtbBjbm4q2yJw2EZIPVvgqLXa
MmfnnRHpXeIcfUqFJTAVh+jIe6nViWhIMDe8zps04lz3jG/0iXlCVGVWrKkCKeX/
FBqNGVTIXV/r8srCh/fZMuKl/Gf9aNCHCZ7dGtdTH/y0V7Fx6ULijYPSJEeTHyOw
/zCXSWtsXL2wZQnVAs5yi2ITcQsIQ/WwzTdf9zjCbe6bmtIPyGM73N2S7w6vgN1m
jrocEPeEIugf8lC1L/oeJ1gT1MkOlpMSLQz2a7hHsWYSr/UWIv5juVurMgZZ3TqF
LnyDzfwZk9v5j7lFdMTFDzLCWzKPTycDvyo+TCew9FXq8FuRz14tr50fLxhFTEW+
lOrxsYK5c7w4EeWohs1l66IwL1R4dI2vE7bctULwT7YnSrj43Nfw3eF1tnV47P0x
FtP/pHTkiWvA20SDboYPddfwsQYAQpv0oGsVewPruwXey3whZUVAw1akrp4FaEFM
78rIAdw37q6xrG3tAtbZtZORiFCciHhUeVpMcP2zfbiMefzHbOaY8v20Fe0r5a+S
nxSaENSZKmsChc+vQDfmwFAkuLpda9W6OQrROo0SauBKg/734As4IgFmLInUFnRg
F6ocecPKi43Oowg/Cf+FWWqF0YlX0TEzDyQCyBJeEUBWXEkU0o5/dm7vwQNklbpM
RtC91c/GkbLQxA6WDGp7Y8GRIsH7LbRDOD0cnU3+Z5/3O9dp0H9WU7elCLKvF3+h
fo4ELwr+8QBtjkZIR5zbhLRi6cyTIpOCet5iUqGDAysxA8gKs+5jLsLV9gtnnDrd
bXF3+BrPhLHxVx8Oa3nGWPNHzs8AlznRKgTidIqC/dbuC8tmem0MMNLOCYXG6vjV
Br3d39THjw1n56LOAX70tP4AonsVckY2BxItLLb8QyduN/DJu9Y4pyFPnFn/k5Lm
qsVfRpHEErtefymD8m+MJbOskQ1LorehXPal8riJsG5yDC6XZsGvW/lG1w1etrBk
+qwo+seiar3az60u1DGUSXsPlc4SHDKRwhAjfXP6odvaKmQbL67F6s6MoCBXu2m4
Ns3Ob9a/Iu5MFqFKKBIqwPMLAqt/oXIcDScOQ3tAkV7BTcIspm/Py/3TiIGMS9C1
WZtvQifhu0a0MMYbbXKy2SL/+PYi4paRt9z5sBekxpUJ5jHxKvKVofkgbB2XTiad
s24cQKWsaycM7pCNVKA6wREieCzHLs1Ihip+OXGc7a09nEpoygjYavKsECVl/BJE
mx/3BYyTqWw01NPrD0zuzSaGe3sCYfUOSsb3sTHWCrNL8gAg9eSwQFgjgySuyNV/
4GSaHsjKsnxdKCmPIEC6PmnO6SKosRDZetzjNQnjM8MEeznJj55H+UY/JIGfKGCL
gqQ2QgD98xN7XaJxAziWrz76tOOZNtKwSPBEaVqk3DTePR+w0ClG6hfW1nvxSXOJ
l/2ORR1Bb29+7hOIyXK3ZuB6tQldvotlPwS3hrXjyxnWeaO74eXm/nRyHYTJLAxs
HEh5G58qpns1ylLa7m4j6+Vzf47xJo0P+JtasAKwLMVIALPMYGGopbGaT1xbFss8
4ar9ugUySmpI0XRFn6SI4W9JK/C1D8nrCReMRPgQb2COzMYywYkF4lhJnFSsrDD1
qNyMVUOFNBf/hTwGyPAPKa+htp3YNzT3tmxOCLRvG3sbBoJJCFDm921ZxdSn2G/O
Xo2Ch7fU1ddWEVIRQwK6eNAylxq4hrZHY8lkT0DpKm/6kBRl4fbsQmB/AY3x0gJV
2Fs3f2L49gjPani133oJjrnbuVaMQJxYSPqXGBiKh4F8YY84ZTh2V5m/kl3dnPQ/
BsK00Wp/WBR3jVqo+8raATVRf5riVoy8u6zkt8Ru2irJ4qBCRLwG7gQaRVg2tvMF
gjUmaK5PZe3U6vMB3eK4fUokez34n3LPrbIPOldFthlcHj/O/Knb1jerK/N5jSgn
2bjGT2yMcPqYl6o3N4xu8DAuUxEZFwp+jaeoCn0AT4Mqn1Jur199C0AjDza/C3sn
AvzsZMyjiBdHzjqfSxuVAb0s9p6NsvDdlcKgQFmsDLX9sdydKemQSdc/K4BZNZwJ
C21lZULPZYWjvkDD3PZAjbL2u2RYT1nR892023Rk0DAWlvEW8JTbfR7KgIAG7saP
jIxFniN25lz7oPG/9M+mjUe6ZAXU/hTbjUN6uHya+phdDB3JLK9MgW0l14nezZI9
gEyl+3DXcu8qpEcIyWc8RJsMPoYkhBcIxNrc1M9mEa03ITWwoT8gSa75/s9778BF
/L4wTPXzl2EDMBuunWxkWuch/LHQhHjOSi6sfRtonVdXnBvs/I/Cnf21BoF/BqBy
3WgsAaPH1rRiETcwI0ACMz8hi2li8ejd/0BG50q+bIlms0AoOSZsBbnI54A+2IM8
IxlwPiJcUxzDCyVg69yFTYrLvBYZte5TAv5LlO+RKEWIEJnC3vI6Qo2g2FzjisuX
NJU7dvvBFcNKmJEmrn9Tt0QKI/onOyi3O9DFR/mzGgpf5HhTRDEhTbMpjSkbEHaF
GqSnZh0HNbmgMCXjLMZK0d1TzDJPDSGRWZBOFoSvCMlKNLcOIwp8a7Yudkw3xdf4
orSROxRe6alNsOH9USpG8ZkSQ6laXs+YFuj5FTbruKaDHrI+1grSfGveODq4pihX
WZ54xpNZYaPx03YwvwhzllR+KnO9n3NgOs73qIfNA2jAMg6nX+1nvmOV30y0v8ru
DUdi6tpAlI34nQYFmmI5yhjyCfVW0QirTB3RaFlcGRuB03Y1fmCRJHJykhGEhB01
EkPXg0DWQrZWgoAeDW0LhkChcgKBYEgxcKAQH+2Y76u3OdiCTzB98JkB0ckUoHY0
v7VM3BSwnP6Sr6JFD7D+14gDXvK6hDQkBHXe6VYyomlQRw0WZ8p9GNEaSi7fPX4g
+EUWpayDnSo8zwdlP3iAya3goHo2TiZo6h/eRoJHQHypgo8UcCmQrmBFVwhGOoqe
WHyEFT/ypC3JyDdciE/Lx1Swkboe5cGZ5cp3WKjbi4pfYYVzdv1eJDv+XOOWI6uF
jLTkE90/rkx52M6lOZytUJaDHm5kYqJ80qsD03DSXSvk4ZhmpGT85fme49R5yhyS
hNlDdm9yb/HYFausQH69yCnoysunKuge+hFkdUi2TubkAA6FCpGxnaYAjRXCi1LL
zv6KOD2fLYLB0AFTv1wcrlBEVR/TKkEbdjDiX1IFos+6yCB4ktkKTIFT6xsciKWX
IBd+aXQxKcfpfutq+tCE7sViYgUy7dDGi+fVaOcu5rD6bwDUiVUzVB7CBNs8XEke
XWCMyGe7Qm7EJm61v7Uazo2mVMu4fOoczTmLxCMIthBoyAvViH5kH/nzsZ5c72W5
tXlzYZdeq52EzgaK+sbbCQWugLZHx9m+h249gcBrG6DLg0tsPF1rXwyeCTIn0vSf
dB50eR02BFP5n4e+xFaJIqQyIoNfQHLkmIR1QW6B7tYMd/YMED2zJWm5HerKxQ+x
rAt4QEvuVxCGjK1jbIJo3smgkr1rLX7fgPlUGgNJHOHWKgaGsh4Ft/RGX2nO8M6P
ZtV4X3aDV6dqgQss2Q+x2nMsDBxWauc6z7oOXs2CxWJ8YT6PcuE367xE9fHrbKYZ
BBScCLqmsAVa0b7q6vU94rksgHiO1xQICA/sOVrS7B+09SSyc579qztZi3U6Ngvp
Hk4tfJTnRMVcr+EpWtcd8SvbApTOsMD44opkUoPvlSTsuzU1+0g3XLVjgE7JU2ec
7zn7DlK8T2WI4NG/lT4sJC3AX45lMEUMHat7b1H65CjjbOtgfVw8ir0wfhGPU5pd
DYHgCeE3pwXRumIH/+JnViUnZxxoFTzGmHCnto1QGfqciIpAL/Nl25B8ZITycLiA
fZjScQUtT8cdHXkjGjNBWEvOSFpgf1OH1slG4gW5eqVa7IjKKg9SplAoWaquV3Om
Po74GJGS+5Hw1cLI3Av0zm8ZaXxY3nhIyPtlYxMuvHgn2Nf1hoCTqXBSNZsoru4x
25Ph9zC/lFbIbPKNKHcEW0kBo0MU63s5A5akZ9GS40wfHTdVQRKkOz2DpHRH5V44
VBuowznWDzdmJUgBZ6+Jv9iN/QFwbCYxsMeHbkeMgNs+bIantvM1rY90gtEdk0eL
/os4kWvSl9CbLsD7i17zoOSFqAtm+ByObgPwnBzQ0aDXGaEUXLgfJQILzhkoCbB9
plL1BaYYXxX8iZa+pb1YnbO/IbUQ0ZoSnJSeiZ8Mw1rjVfX6dtfWXox49bW/CfBm
x7bXFU7XcqlcJESvsV1I5Zx7yCM8F4ZwtjfqEAuxL9zir5okWA+l7HaMQc59luVY
X4r3BoeLSGq035cFT5fB6z8NYDl20VWPP4XUefkRcjbQxl0dnTfaL4CGZrCK037B
mXim9Ir9w6/YuxVh+puQndg93pq0iD+S52LO3xL6Y65iIip3CPon+RfSXM9KAEIg
ESIcr5FY00p/7HAFvSOpBM5MVg4+G9D60Jb3VLaEjI6zAvET9pyAzWuQbNwFU0tG
KcRA2NxmpLZ2Cjz1HFzxZkurVHDeSFn4Y8vmn1nBy/l3OzvitCsdmEp0pe6rG9QK
ZJKeWMslkVu9drRfE6Emth0TCofBiUiT7Pc6Mjs08rh2BEG3u9GpASxVkmOWSEDT
/Z8izqXsm3LEaKbMfzfCyUQd6uixxnqXOsuh0Hv71bJ+zZ5+3vXQvhjTUH9/MkgT
hGU7IF0LTX8ZmuTCN8v7Qxduw6U8A5EzfsSiRVDK3fBXLPs5Jle7xfakSiW8JfvI
JL4cUX+NwYgbfBWprYV3ZFsmGGcpFlmgUKlTcn+A6XASdQZNrY3L0awe5NVEmXRM
pmK89cE8eKXXJleKtOOk9svePseFQIuvFOcuG+FwV4mEQhw31KdXaeFjjixOu9rH
FfYSCba733hbP77ddOEX/3XJDONqhsSWyTuf+tGsVHMgOC/lBm74l1NSYPIW4idy
gpaKMkeuEd/3foIAzXD/TNwD6HDb5kv1unpxMyoDfG8LtSLPy6KezF529neWRwvL
TdorkEuVlWVDj3bmHWpSogMHnBU1xC+ufmqmiHc69o/qI93ELWPNkEOgRdyvneuI
DfEyh7Jv47mJ7kKaHCM9qtz4RNFWc2dZQdRqImC79exFQHRQNunD2tLgAB1ZKqAj
rrQeaC6ORxOW/7zq4E8SHT66zglo5xaPOKnLWaY30whdhyaTG5epQS9m5hoT6PiU
d2LdG9yEssxKCPgQMzvRTuYUqDKud5cwwC/vZVfpOzDBfL9QM5hQfh6G68qkJFtH
Hk5pxuv5X6Xf2zGndMP21OBxpp/e6xa8kwMLz16bEDm6mFo1DDXOy7XX8IXzwpsm
F8nMW3eWETxADKACZafViazgMXAweEkgeI5pPVdNK24D7ULDx6JQZ5KfC0DREFn6
VFMiEjAlYNl8KkOzw1vbdSh1grY6yQOoiJB4adf0ZVfR2XiKWC+9YjwitXWyX33F
R/iBrFg52HnV4j40101VMz+/NQ0LRlxmGWs8jr5rihCyLzhKtFgYIQdodKVTNCYb
RbKTjog7ForMagVazOnFJtfNGFmilgB155ltPqToaDTlz4ALYeTVa7Oo0Swm7hst
+if561LSmRdrFRuE6wMIGGbZ9FHwIvMdQdU21hoYAchaAFiYNqe8b7ulsGsIbq3+
/OCGfZ0sj1FBvxdGOhLQ7wUYs1PSbI3ol+42PqLF6c6081oECbqIXAEM4yEYIeg2
HSk9C+NL4S/xi9rwJF6FWHMfjlWEwvpIat2KwFrKXBAQfBtGi9k1Jyx6Nk8dahDe
FRmvWG4szcPXGnyioe94htLnKVBc0d4TsI84qXh4oFXk9kEEbnQNBGh2L4QiJXwh
3qQRvF8OYi4OGTg/dUriEhDemgunwqyU4lIh2dk5dMICNuyvQSYrKmjXYwaCRaUu
k2wpnB5K6VpAYaHjYyHc7CKSkq+/epSBDJZUNaN/q2boFFa6W7XkhiJlPTnUmL89
2VVofv2Azmipwey7x3XtJLHF0zenTTICKagUBLXJzGUogmzSSSmtjC8X3/6r5pEf
XG4u4jF85amKC2g9/ywlo4mMxjebOvQM+GGiTkKQOW94y99ayLA8eW9icQ6XwmOa
WrmqHSJoG87SOew5oy6cg2Aahygwqx9BcgUazXTEWnR+/vcXb5uSQPVL4JuQyvqm
B8UpNrh5dXAwIuyj62KN+3aeV0y79iUIHWIaj1hBPek+tzn1U3Ssznt+DibTAZ7Z
BtL2P7gI8x3H2oMjEwf49jFd9MnISnv96FbHj/jyltak2YYUKZOKU5ui6t7ke2qr
bGbvnGlxEg1J96hwpsGPd5ocTwbs6Lw1iTfADREcjFeTtYdDk9pDX4NNGqerWci1
Vq0B06vIFaLNc/tX2WBOGWgecHQZcVPS8FYjr3AzzWjaOP68vnpCEmQA8Hx87S0K
8QIVEkRn/9lhkR24u1lm+Bc4eFKkpVnpRcE9H4wdwu00ngVh95+3XNw5QIRDqUJ9
UxmiNMVneeCJKk8ZfIePH1enVt2VPEPPDVHuI2vkrzk/ZOlnaaGQ30DbZYd4u/9+
os2f9/B2dELKVWfKA6QVoQ7s8tmQNN/+3V7dSfYL9Hx7ubr00JjBa3xe8jpkTvLM
SG2XyJZpSeB0Fya/vdVhxahY+eLNrX6Y45mYL56LOZ16mZ40VZ/7s9BNJARU7vai
FT/NgCaZY64PcoITJ2UGQtIu6yaiaacA6MvaRhe4DKclaMZbOeSNYl+XoD7KL14e
Nu//VpU532Q4QquIKtCuUOAEL0a0TU1wIoEpj2P5e+Ay3Y1QlLP+FcuI/YIWAIsm
YAXZWv/cDD3iazbNTO3xhiwBXNk9jn0E/nr8wQKBgkOf9odHHqbuwoHCGgs0rf6p
0v7n8YvpuVNyJk8v1mbbPXoQq0UWfVnMDHPNMkh49HUFL2B3qEAunqASUmuPAsOr
SIVoy2AP7vzeijPkJFGrn83sh56fq16VVQuVxcFhccltPbpVeHVprHLK+NrVGEY+
EA2+SQyVofQa3OO/f284xk1mIhLpbvZZIUG6a0ZdjbiXX+qC5nPvfI4ueg9zsCKI
Bi0vlziJj8LtG5G7t58MjSYhtkqy2d/6It4V5TQVn7Jj6dK7H9aL4jwUr5avhAu6
G1fJUFdFPg0xKNF3/DM34nUkL2aqTlNHdOzB1MdTfqTAVLgvffP7veFR0sbSF6UJ
sXn/7tNBqwSiqzyu9UWh0T9KWrMRFLMIqee3ha9u4ntvOJ7OFrt5BBo1lMRMpYYP
qM2ZEfDIbif/dblyg67iKqbQQKPYp2TPOD3cQFbf/blW0e8lkMzx0vtpfpiSIn+p
yaUuM3a4SQZtA6cVbgQXqlUyeNNAqt497rPR2fy6E1pkwacIwNNaZ9f2Fj1ljBaW
DsROsecAO4ZsUmbO9KlkzOMutD6xWHR9YZsOeGPnt/Q1lDu5MSX2Y1p/+Uh5tz3x
VG0TOyHzkMVQHyZ7lqvRFDI7KmDCf7lRWYb+syTt45Zlv4CgFCL5IrZz3Z3ArDse
NmcgpkVXT69ZxiQHD9IgeA==
`protect END_PROTECTED
