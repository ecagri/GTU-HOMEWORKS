`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Uqv/vN2EUlZg0Khee55Zx1kstslosi9K+OpmbM/ZJpzHkxa4Okts5mhWjGHILlr
LMBoL2FNj1oWlTVaPnbprbon4MOP5OFG+lILoxAgoxW+Zqc7fhLDMZ/GGdDeMo5m
hItt7e8ay9T6KqpGF/1AnjQnp5Y/MaDi8Ewckl081mJTpDj1m5vITGazGrzR8+Pd
EzDbxOXlhVn6xq+g6IrBGFrkvMX7C/tVlGjXzmeyPeHQqlzV2VWdEMJ3XSfQWenk
05zEsx5/0RHFzo2o5hInTguPzTfgWkK3YTdNjZKwcNotgRFUPg1xEjEOgH0OwHjY
NcQ693h2bBSNC691aeLyj1Fm9bPL5+FIW1Fo14jVBjVeU3UqY/pf1RXqY8Hdmpr2
TyfZyQlSKkcEnUco9tUcWWKUnb+S21LTDrUmUbL4/jpGXwp3/TtUCHmbFSa+PLFY
nco4sUBvvoL4IaEXsahSeNHaIDcpo5Xge3i5qIj8h988s3S/UNurBWQfg4zbdN0a
3CnbIy2/Ib7CG6w9SnEfgIW0VxbMhIYQ+OA1UcsoVdfX5fhLV4ZlWrmQbExfqjBe
J3bBskzlKmDCsNw+Y5yZhzHCL5ggR59fa3MRvwEReGYlmHkrF9ConkkV4rxyo54t
chA+6WOMZO7kKC7yBVdSG/Ae5xq5n0z6BQSUbgQ9y+dl5vNY9Fz+vTsCsWlAohaZ
jjzgr47DM1l119+Iesu03IU5ZGdv2tn+bpCh2C0kVwAg/zZN+/upp2v+Qanw4kGX
lDclCw+zF3E7VNymprFdOB+1SIO65X4gYfxUDlEkQrpHfrJHTXswwrRYhJ/j4YxT
hRZYKeyWUEt7qKWZY8JLbwYZ7ahFs0IO5ZzBtpXtoHshpFKTqsA9IeJCTi/48dgY
CifkbAP9DKsPWl2EW7ZuMng8xIvpD7jDo8LdnHQN9Zj+Fqc0OY7AGXvzAsloje97
7pZrhtuMvy3LllG/WCsfPFPqYAU39wHRPkcWMLjKd/tbv83gz7jGV7wac+NXhDad
f8IW7n6hWMaHPZidh4cfUrN7VOgKpPKuZvMSvE7u2E4kiRFOLspjarAitajZOcDA
bZDenRF5jMnEAaNFTgHtmPIpfi/9rzowvgxlyRg4K122wmf1EkTaFAOI/6VCRCMl
EER3fWJ/Hm0uIcufT1tNf+gYB6ccfOLdb8uX7F7ZOJI4F1Tng62Nfe/pgfyv/HW3
+1djl7Ag+ZpNYA8ve9dSLppRG7uXR0vRKTpjce01BWW4SVSAIcT0OeeloTTl0ZGW
JGZiKTxCt+1CjX7VzooF9TTjyQgMHU/MdJuhwJF3EoZ9ggxhTF5U70+lZH0he5Sv
7KHq8fU4WHBKfTpUVcf1T7Eyi8giQBmW7nkTVxOYe3bQ/aD3rxNteRYTpAnbcl1P
nSaxN/+vF3ln+UOxPFRfKRg4pIRcXyHMmpDzKt9bDiB0a+59ZcIBdZGY/Y5jHE07
Xifz8f2UG6AOl8SV6izdBMvkEBsgduqaCetVfm4RbNkKuiEk2rr2kEUfdG7iyW7c
xVa/R6KnllF7PpACaUMq4GnybtN7PaVI66Iz26KTAwgg9t1VQNP1F6E2P9PgIZ/m
6K1mbDHidGK6Z0bnRFZuaLxfpP4HZN3Fo7uj6uz4MQCOG0npJsdmsOee0LTLGbOv
6PfUhLUfWsXonh3dXC57ILPb1xmu5vnObPewX1y/XGxFmoxB3SEJ0le6ev4b9FIF
KSr8RMNRALwSQvEccxO12GXdekHZFlQkiUaIES211kXYGnzQUrzAIoqRJNcoWV1S
3Oi4Si+sMcUSkHjFjjoT5mnLKRrxOO9fcn9qERTyq9lAAYvap4cfP20yVp9DLpJP
wM2DFWdb9KfrpUPybvwSMPbvxARDxaSn2rKP+o1bX1fME/Pm3HCjpkBt+hrBm81o
WM3DlFFclBehLM0K354f/6Y+UFSLN8iBMKZ0moMxE0XE/7toCPaFnKlTOubBuPeN
2VBsal2bxrocByY70pJFOk1ECt1T8vSHj3hPt6vgU5fAPAEIP5HdkP97Lo7BEdO+
4at3JB4kFxeeNOuALpb/Fkb7eCxHOVKaEY9HJCR1/aDfHn3vRiU0zrD6sMLbV6R/
dW2dgIrP3gbsCoAt09RV6j7gUrKXOO1OTrjWnMhPwzNzlTT9nypsqggZS0mCFgYQ
qol+o018+on676DMGs2OHUPUCC1W+OOpA3gkPHifW2hxWMqwzDQb4Zaq/65pddnu
Qw0xyiIFc3xOqrxi+fqoEv8O1Io1Wiyg8j1d6U9yxFRdjr+87H2KOHTsd7tYrnBz
o5w+/GJWFDbJkyXqsQGSVxmh7PVRU3//MggLcbdYhEE=
`protect END_PROTECTED
