`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bx0f+AX9nSSNKVFxZ61UkonyH6qhLz7xFfZ2DAdWF3QSEOO8HIBBMPIqn2LStUeK
I+bs4DqfWem0ogLT5gGau1tT3jj68oQvlspi4HCQQKgDcsFNbjAIL0wu1x8T9ehj
TUfY1I8nFsMr8K0fTeb4Ty3Do7JwEDi8BwJqxRWrtJkZJasOBqBEG5S+C4EcpXTx
GXp2in3ZRzGlFTZIhKiUyZJj8CzbmI6ZlBoB6c5EvRGM+RiSIAyPGVeBhAQGkSCa
UMjPkxK8+EG53G4mld0CTxcUHAqUA7DG5wJXBQEmk17dc92l61GmOOOxJXk0vaDI
jAKb29LTJ1holFzKRt0r7YrAANGOBgFcEnSuGB+Vhxqu0Vqf3VqR0K9Q1j3SM1vk
3F0jCFOEJmWBKKGOLYPOFEnL67x3GGcgGVLPy0b4NlP84Xn+j/6qZkJ8SEAH1DV7
LWXrzsW8lcWUv5YG3993kFzHedlF6oF2wqsQrh+09bTol+IuzbMl7HFW473X4iHG
5zkEzYVDTTSPxJxxvKLs57o43UcK7d46Z79b9Qca5dBuvBW11rYFFcVcEpHvqqwl
Ctt3GVP2EZHPgn850iiSg3uB50HJRiYGhO6WzLnxq65ppSuL37auNyJ7X/fQzOXG
iOQUO7zJrJ2dBQhb7jMh4mT0ObVL4PQgVb0jqvVnSKabNhQ8RWyYy4LsGNbcTG1D
5Ymh91Y+2Jq2Lm1ixj7eouZPe8wOFtpOjt51vGHgejNkYr2aiA2l5LnxqK0kMI5E
5Gn8pPbWCxjWtbcC2+lzPRQpJvO/4Qfnz7EJQu5d25OEAGiKtM5ClKlLj9974I21
ZbtLDyiOte2Kv+BNnlDi//SCGODsuC0mVzYOe+qNjYmwtO39NoE82AQcgJ1I2Cj0
6hVkdvEOSyw40CYaVL7/k0bIPcv/aUiNhXCxCXpRVvHFTpn4hCA7+BG/nAiWDUAi
JLm6U0MI6ULr1kO0c5kuDsq7R87YlftSxKAewN9z6INe4GVNu9YzIeCLnCnQJvgv
cUcyhOx0mD2RaH9ZbP2MEAyx00pGLf/pwYA5DXJpkLwjK7G2uwEHA8j5JOATrseE
c6N1bCvuzOUt7kFfmcLsX5BBTpZ7ht6srDMCM6kqLGlMkplI55XhFPMXfV5EWtLo
Xdl+aYpYTUEYafkpkY8yhQbInIbJ+qX5ZTYaHg2/2SmhN2snjmKWz31n9r+OzTJS
5BMVYiBG6YQwTobKn+kWd8L0AZZZTvSGn2ZhjEwe+g76uCV6fBKl8XCU5VDUyBdJ
SaKsxvTLq9pwjwVud03kOq5IZauUFe4L3ar436Lo0kolx4FybV2hXZOr73eZ3B+T
rUkr/0tm40HrV0MRTfb04feBO2BoNYwqM/23/0n+IEfR3dTLh8/ZUsiXYzAXBu+s
pbkMlXQ0DyjVmcO5LTVh3qbSzKYDtghIjptobbzjoLgCEuOnDtbXdzl8tqTmfWNo
SpTrRUfdVL1lHmhOYkpEligOA1Ez/QQfII52W9B4EjshHOXXx+n7zqrLgV1jar7E
f4ZWoV5+5hvZQj2RQrBysHgHf0ISjTZc0J6a2wHXbgQmWUJsiIAlVBegrfoUGoqf
qSInvWXuAHq/wu9tihr1jOCL2lmG5MSNHFzl7fwPQriBCsi677kN6PG/GuSMcUbw
PDMehqjSE4OBP0ZVhD4c0nJ7IgEYTzFQBbqq4I1plnfL9VyqY7QUXNNiYd+QgpQT
H0T2StcqzM2MjZqu+Il5aLIe7W20bTl0uBXTL2LGLBzZqoXdmiJ2+eUg9yGhsNax
1Bmr8w9lz6FjfNoRKMlYd0vERqB7aDnOac/cgANDMSdjatLJ3Udolo1OEap4/5vP
86pWZD/NF66lcFSgjWN6Xo3BbxR5LlXiL/adtAORxBNrtSRDKAG8Cz3/BG+WM2eO
ATLey4oOwP2IXhxpKkJzjYFARvx077cqvvtm+MlGe2WtMwBdQWwBecthAFKt8p2f
Y3iMnJaL56HSXn7M4GRjkSnh1R7d/RrEcoUtzI9y63kOEDVKlogS0Ndopmb9EDb+
YGX+zUQjmDFYgwH7qKD5xsfwwpF++j0U6yqHSShBhKTfkuAVAvo0r7U5noLlXXOT
2PcHCoLQwx2zzBZMQPFDrkCxPf1EXST1ypRvYzW9BHFPqd/F6DJMeZ7HOB6x+tE6
fJ/Toohqt6WZVEf6hWl78kWJI5YgfnnJRkip34oTpDfBaMdOJReVJVeuKincMiUE
Y1YZHXfok++x/0cLkN5wTTaFKxPO7UwJVLxf5pVlfZLY6o9mL9KP6fOg6cC+Db8D
poBvXi2vUZNAQrrmb1tRkmi86+VFVfVUz7IBI0gfvJP9VwL4D9PJo+2FBm96nm3N
cjlSHIyEiFAzCBCGT+n3djxwckP4L7HeoAUiY4/fvFl9AiwFVwkR69jbZSxQ9vxk
1ujU/ARYaH7xKlz9IiK8bSMSM0EZ49X58jP1ZZR190vgTmqkeYRP8ThEmFNTF250
3WfQpChOpFayO083QpapuPPKSKtGh3Us0uNz65pcVaEyjqtV6sU9nnEvoGD5BGKT
X2/YQu4G2K/gytF6S0TDrQEYd8i9mHXSDd8BnCLBF7I3yyGIaumBPTj4tdp6UxXM
PheqJLTb6Uj3qAqCNaPbCD2VuK2Tp30zWCbSlI/kFfp+iA3Hdo6M0M9ULMgLZxQo
XluoezI/UwetRJMDvTKC3e3KxftBrbfH/owaswUi5D+Qd/1GikIABvZPKPZznUOy
AeMnUXgYx7rj/vNlmoRLY6FeRhgXMFOlOb3glwa/AeLpXNGsM24MSYf8DFfRR8XT
WxWSvIz2o/TrerCoTQik8BayV2c7A18PHXFEaOv5nKTevG9O2i3P2n4wNs7E8s2X
ScmQi8lpT/DSgGwvWA8oVzvqmyCGRk3nziMgdcge+1K2vyce7BVVJSO/Hc1OyHYd
mBaevZwYmDxHCSrHdpETiIqkzh2ooH9izewiOVNnsfbg//h9z5fFWpc+xwtGj2ol
9UQ0oSKn9PxRwC5ec16yK06WsT8M4pt4eYdPAK8Jwt2KEweSUoR7wHIHXxNGtJhe
BA2KommWtIBdUSmUbnM5bzowbMss5JMBsGEAOFf2U+GBQhORGUydDuuAs89dUdWr
GyDuJmyQuxlKnaaMe23jMTNatRUWiRLU4ntbd7enHYj1wL7Z0C5X8CP+gf0o5ynD
b3Z7Zb4DsWf2PI4UJdl9V4khphN9LrS78S1UyO+/KZ3TuFpc+wdfMDklp3rO9jZi
0EUUK9KhyjS8v3vRNsoh33f2v3aZ4N4z9vBVbDnogXn2qLQe2xooMwC6Agh+jtRs
3JvHRrxmHHjuq7OLNoXk8pLXeh6O/tYeiOACQjk0ZlxSnszMFx4TDG2ejF1q8rdx
KrksZW8l5U1tQsGcjcFdd0Xj2VQTTbQD6lZWvV6vE44OqgbZU5PebEtU3rClacul
5kxKd5OnAOMlblK9GnRs1+YsISj+5oWCCcBVyle8XXgUjv+0m05xLxTRytb/tdJu
PbUL4q0EyRadT4ObzbPQ76kLb0YdUJiYerH6l9xEmdBUBNEwJrS1h3a6hxSzHrV9
o/yw5G+zBOSkRqFSkN7oG9jFDmO00siC9X58YVjA3OcKPssUgxg5uGTMtWrXUNzo
BmxHccVIcXKRILRq2HRHDoqMBj/Ij+w3+d1QZdb4EL39tgj//X8qjkgfXtGqxzbC
/+mBdaMoQWxEMXKTiMOmNWnAulJvFbYLLl8SSvCvga063g43gyoXF4fKGbNiqSCa
t/3GpNcMYA6nvotlAPNjfCaKbLxluF1T79WyqwSM+L1R2zo1w6aiSUUa8AHp6LRk
Nj7eUVkOrMqSA1h18aBbUVUr3HdyxMy8ENXmZrcU34Xnok9+yWpy0sts35VgAwGz
uG7EYmIJT3a4VEmLxQJQSQ4GjzEsZR8W0XU5F4fE1rIOUojEvD4os5MaZPayiLVz
CJxA85XvMvHfnwD60uedfqTpIUmGL2sEZ64GEDw2e3WVh8RZLIRo2SFy4jk9jzlB
FBbaXgVNn948ZOAP2fP1M23eEdKN+LKEYHv4W2aMOKJFFPXdOWy68G4xuEIhqQfn
ndoF2RHvLPxf4Dkvfqol72JJ61NZiPMfXJd9OVhbXF6zzTWUJQmaQaP4mda/ggJ3
Anxe5PGoapl+WqMX5BicPWGNw9h4sBsn/6hiuILNG/bQPBmMLtSjT5Hva/jUBZDB
7fhxErVqKqPsLwH9Q1OpeYowjrebQOT9jkR0qFKyqTh1b+jDjjYsTVT/JxDThHYB
B3pSudptHcP+B1pqouoLVJN8j7+dAaTceLWIMO6QpK6Kn5xd58iCyEvMJ6oTCCdQ
VMVbdYE4lMAtS24nu/XgWxNPCXZ3HTNYry+cX+an3JXlziBMqIlHu/EXElgSqawG
WsWV4ZAchkC6ZnSeANSgwiThfi5YT9glV7JeLGdhEum05GozA9OKavBEuX1YR9+a
iJtZHYQJ29oulLbKQ4fAbIc6pcW1wVo7DAveiI0QZjWeLlNWdX38eiLWLLgiJjXH
34WsJ7CpFZFg7AaJ+0LKfxNtqvIpLnm+7NyStDyZOU8VcocKHRs+xIea1NZ7RnF/
QN7t3zZaGM3XbnGTZXqQrlOi6JU/Br+2IV81sD5yGacOIfUCZvwG8fko6iOZ1UCp
sPzhJlzD+bzFfwWRwF0B6N9Zg6ME1Dx4OOKZM1uXbpVEYgDfpuppRPFlOnC3mz+c
1MGAxFkYuJqm5ZnVUg4oCNH72LcsSlb9T8e13hji5BAtM6hO+4OAEU0TclTrMdEQ
w+VgqhJUJDihVEtBJcNiXj3oBmoB84sIrQz93UjYQECxbrOcJ8VIGu1gR63xUfnw
Xmnau7oKkwSe6dNnRzcIUgZ7kE48VCEUaTf1cwFY2/zDZ/t6kY+kd4QgZABBFRlA
maoDhSbEAhP/+4eYA7ollLp+DGESCNeqyaCnEF4ljuaVQE/6lOgXtFZ0JlMuEcHT
wT06M77+KotBUa8FZ+PkL+1C8dwG+8wY8vJob+qjlxdAEHtE4e2XPHe+S3zKGeh6
CIYqDLbZ292PptnIysV0E8SOPzygMvsFye+9ibfKqpm62VE4K3uDmWoGyfeiYoQV
YTQNJYA1HcozKy2rU7bTy9/OWOjEzXNhr4fcRrxEYR/9zVR4+/ptyEtpo3Sh6EWQ
1v65RlvDSe/PdHZBFhi5RvOn9MN21nao83ry/4zTI5E9jBBGw79lJRNJsnUDHG+t
/khRpiHCSSts+dQ3aX/YgeKZP+SRAAw03rwwTq1V8vNx8b0UjJj3H3l37JzULjdN
ryjEMqMa0n8JnuBxwmuepeBWlTGnDX7a87T7+sIx+RGZO84RrfH6sSIlc2u3rSvA
R4bXb8sV0yp9TogTLEi180YOQ9tXwuS8eXBfJieBkruugAvNbEcwogcLc5I99DS3
a1kiE7zmNAPfAEmuY0+ASS/o//dXGH9mbq7HECXYxkiJzgXr46Uau6OE3ZhkvG1O
KFGF1MpFX3DNqd6g3zOA9hD1lIih5mgWKKi/8ysrG9IvLIUnJe1Gjy0gRPOP/DIB
W8piRWJF0EOkBooMRQaqf5RDx23XoGk12gRTlZc6WxdK5hh6AnizHF/H9JAGcdJ0
/trTZoEi5kaL+j7u8voImoF8nl8FjoAt3hLd1YebFSMiDDsqg9w7wjzzBWPmvKyM
mXqAw6U6XcBlYq4b3m0fKw5Vrhj2iGH0ygm+zxmwVPp+VSlTZXgNebZTyCz5lTad
dzNX2B0K3evLQpuK1+Ivvo9sGF6WZQ6TAZBS1cSQvWV2Q1zKJZcrNCvTbecu3k7d
jWsPtVSRQ6fwNzsL4/V+No3uGmip5UfVoxccu3/OS82gMbHreWT87EHpRLVnwQtf
/78NmwIPudZFOm3k8LLrOagIQI+tT1r/pB2hvjW2TWhFVH697bY5BWg/NFTONlnj
3Z8CNLrwpJ10TT7EpArIam+4oxncoVfF/lX0KvGfOdQUPL/tU8T8US6LYSkeR3TY
3ImW4Qep+ZoYw9zhqfdL4TDodW1E5LBWVIFxmQ6ieiktYQAD6y1oFfxvb8Rkd9kF
AXnqpRrmra/XYgz98/MEktXGDglCzNtDJbrtdcHiQGG6lDjZkoTOfz6c+IcFCy1c
BGArvRsiV+vJ6rjZPxRpGty0VjRegNMaHgkgUcgDTHjKx+7r5p2Uz8MCUzR2OifM
CMUVTfpayGWRgwFtmmTpm8vVTAsc5vTewOJlMejf/AzVFeybJvC/JbXSi/wo7rwO
dAtUR05R63qHzdKPKqasu9HeZ901mEwWJPc8q4BZe98S2Pm5PNXR5R9yjtGhQFfJ
FFHa2ae7iyhCo/t7BP+oHMBT+cCecHpr1fiDHjCszNoQ6mW06GQZV7j2BOLWlDlP
f6oSggPqMmaBp6I7OOaZ9PZrs0sYnvkhQboSCLWx296/rmoRrBZSSsrR8BAEY+tR
ilCWh1vQcG00penSvL8rXORZXkwCFlIbgrFy9YrOyZHzKTXj7/2miS32oir14ZHw
JRNB/40AG7Wv+JJo9bu/dzGAsUqdg6lpBKrVPKK8x10bMNtLVAxXcW2uIiyI0zyi
gTqIH3zYGPKb9rENSUJJpGPtPDQMPjv3zUi+6MZTV2LZhX7WdRh+bGOPZJFjbIjx
JaQ2n7bUjh5sgvB0hbyUe5YKu28ydAJ327s8S6Tj274NFa6RYGNfnTGnU38lhd5K
uU04I6WlVMV+2uTdTH2CFGwvyPCwsUvM7mwYNRTgqkRa236eJC++yr1qgoQjpqU8
yMRtHs+jMwG3S0HGYB0OB55XibNXbaubprghba4gvtbvdABn0rcM4n7AbReTUnFl
JegZrHrLh95AnB++7xN/B67gZtNaB4S+axofZhHz7Zj6/44a/GU4GeDPx4Izf6Kc
1AOhxscvWthuVNrfsZTmbg3Sd1iXAWU38IgxQ7U+GBX54iguMEPHKL5uqNvgpHSt
iUyiUV1P4tYTNCsNTN5MGDvIEoHzE8yzL5kfvHGstVHYEOADzpNv+gm1x3eUfDsk
Bq/r+n7p1mr0pa3Iwn43+a41gySoKwoGgqbYIXRyXwQA2pYACjOuBsNtHGPXKWk+
1Enz3WDWgtyWy3u+YpnnftIOtIT7SonYu4ma/Q7L3KKtpW/Cd1wxZk/MUoxAZSUv
3ooRy5YJ/rJ8JpRc0SKG6ba/pATZlOu3hrUotdlIS8JMm8mUzU5BUm+aMXHP04zP
fLUrRddDVveMh/RZOpuc/3/TdEEOTfMzXlXCo7NTB/fWimqYUzQ3aMhi0R89xRT5
pnACs5OHwPnU3nn3ps5Pm6DWq+Ja4o1lqYfN2gF2+srhSRqXNU1wGGZI+NB7q8yq
x222ET0GQEqkcOpTEhqyrg+lnupAsxHIYLe/NPn1m+o5kMG+KNtUalz3stbmOEqB
2J5m8sAfKu4XfIWoPNs+DyK9z7ov0YB6Ej/V5mq5nMJS+s5lA4N4NOdHuXgBIIXk
YdRoEErLaedWx+8Le/r+6HZwl5GCHnjYrmQztYUt1lV2dkWlMt/arNcSbXEzBoJR
V5hnenZghHg5tX5iVlfJwJ+ZZoVljnsigy5+lw+SHVOl87bFhuvwbeEmS19WSpYP
7sA5WEwZ+jfORnHuAk/5Ov/Gbb6p9ArNOw91bmfOTSyv6PNR3Q2dNOj350lWxRix
GqKjmLWfbqrMunopDu+bdq9LTyhCdAf2htFcG8ej0VvSYn7Du8geT2zf/m7ydeea
tZ9ldggtKYnX6HDKpi8MVrlnY/i7nkw2A1Fn6be8usnT9NZ00nCJWdcc1rCXpNMQ
5VcTCaXxe7gOpuFH33q5drgJmv3IVAnP/dWq9Shf5Rpg9cMGuHXTKTvy7eSOingT
T6eQKQRUvPcfkGKceBVNnU8iHyxe9vLGNjETell2VN3sj4sjFGVDUdRl2wijqNlz
9hF0pVuENQx3lChGTSGrHg==
`protect END_PROTECTED
