`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DkoNwqNSQFSi/GOQlde6zYbCTe2I5mtVzhj+SwyK18h/b+RSZu0AY/HMpPfwz8YO
QIykuO+5rokchn3Nkt7uHTur4QaWxz41D5nPoaGRkK6AJEan5+79Qy3yh4a9QfdQ
x5ninBvtVE6wOMzBZvdQB1EjA1bcYkuxsmipH01LBK9n+R/MvJN9ZWRHi2mxl8QO
MZkG7BgSNfyg5Hr20L15wWLfIjCyRSvC5eo4SUuGeEuAA5hoYIltH5aOxnL4q4lo
jZZ5XAVBzlaf0Nj8VDqYCbnm/cb075D6OzoD82RRq+9YsSIMfi9qYCPxqmB733oV
UrKNTooILf761YZAne0H/a9pPTRnlD6FMSrAIZA+kCImxuU0WN+s/crZiASQykJJ
jaMlSKG9dMZhRyC2FbMQuezLD4hBBayWjTO4SEoa8jlKMI/w2jeiTRIvN7vaY3xM
RsAEpakV85VIjXQxDwVydIk6sNOzIM4CoRC6U6O+Yu5wq8FQLoyTUpdP+PWJ8pPp
BiOUq6+KOIMdC6UhkZwOSOcdnkTz7EmGTKs/QilMRYO/QJOlJ+PXRn/oUJvycgUm
Z+A1nJys6ysAJvDZd47Hnoa3BJtYTyc4ahVlNI1ZkkQ=
`protect END_PROTECTED
