`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OY+N7md6RG4IThHRQ8pxu9w4PQJH+ipmDbOrrPSURcPmvIAhJD1TUbx2b+68MjPk
cTVOt5HSmzLePztZHVBdNAvIJTW992PQkDyxVvwPnB/hg6ccBHHeAyli1Bs9V+xF
OjgKIJRA7qeZ75KvhYyCH43KrOYqtBulZwAq+oYC0/K37NgVojgaVmIRkay1Otis
dDcOGo7gEO5v5jpZ44CnY0BE7GS+BquLsFRZK+hsDl8Km4OU1C9ANMmotqOd7Iw3
YHlrfsv0AbWCm10uM+DV86+UV5kWWna0+a32aZZablh9kXtyHha0ooP0rJ0vK3eA
QkmIXSckps0moq01oxPfCcsFyEWiNjJ94TeLZ7h4JCVrgV1+EP+x9hCUjYZQclrA
aqsACq6X9hGB4E8BQUw7dZnnLmD4Qz3QBqFVmfvxkhOTkL25aoJHNxVqUWtzyyTB
BTw9G7l36N+RDz55D8NUpYv7JSxHV+IsXSW9uun+emXxlU6F3L6HSXlYQ3oxHIbV
W4ie/aCrqc3yTykNb3zgumPJfY7B4tvy+MWHThTVBJh39CIRmEUmD3TDTwnYccbd
ecKQ7mVX0MYjCTzic5scIfUyCM4T1dbaIgrT6ui6kek+a1PjAHZoYEmFHZnE1GNf
RiFA5o6zixPXazlphD1MQ+NIoRguNQLM+fST8y0niRkfKNtBa33ZmEoS0uO1DhLf
UJadnqT7bn2c03mkjR7Mn7b5STNLRAqpJo/mq4kGUR8IWvtjpMvvbOHewyf31P6A
QroUDK7vLR5EwrausfpkJhh86ASadcQYtGieH2xaKDyTKBqf8MqmKRkc523tm53Y
cc7C5HLfuoyRnB8zxPxHEgGv12lTTmzjnqDEGlrqo/v87wH8uYVAaT/3B8iuZ09E
eji627Hh1xz1qdoWdMY3ZRoNlyNdQGGdES8YuG6Zy2U2FGcyF3FG427SSp5SdHLc
7fxpxTJdNJ+TovZIolXfdzRY9WXeaCELjLxNva5c/qrU2hhEIZaIBB4gS7AwrhY4
e3rmCWQB7z+AxvwRgBpz3dVNjpz6LqHtahJxMPb7ETDblT0QGIchXUXk5a1xhgpb
W0FkQK8DYDnZhdI/OHVaa8l7sJktq8YiVGRQ/uuIcgKQujirxMjJN2frYdLibb1V
3sg37LhJWz1pCg9NHlDlpmWf+VHRHDIPG+yKxEtpPyiNy7rJtEPAsWL6pefwFEcO
p9Z+nljYuK5UySIJm6+PRcgS5LSfGxt1mZ1K8bxlQFkVjPcm0HeaWCQ9hqcm9LHZ
Xo2KbxI6uZgYQIaqitcLgOs8XmhJieXirV7Obg0mrXfoqhtMot293K0XoId4jLRB
Ll1WAjCQQiiVpGpEk5gTxtzKwj4H25hrlkG7jqjtu/YonojZrupTZnUHalg4y4xj
YDJVmAt9B5c0SGUunKM15ZJbxTZuMVSs3/vPwcC5vJcryC8T3FyrsmE63vdGYepr
eKzcj1Vj2gX1D+7eNdnAdfywmXaJHz4VqkcQKdwfmPLc1zrxqWXmsnKo6yFKoqf9
EwEs92fs4AMbOhagiQVHGf95rbSUxCvGx5iDz6e04zX54132gzLuRL5F6GatLv+6
nx0QkOZ5pAWYANTnAhZXMJBLcKTWM61FxL+/ndjOj7MM2YD/E/z1ejSgnAAWR91V
VqE1hkQ+q2XzlOtVOOX8okgjI2ubw4nmsO4p02+ybg0OLfF0uVA/KNdXaA8nhBp7
I/hwTacy86KMCgiNcjFdj9eyNF3cDkN6gPvV8Y5XmZuO9aHzmCAKBlrJAfPNN5jW
h+js0i2yFYOhWPFzxXXNINAytUyFswvPMg5KDkB/AfuZ9xieSvbCHZr9hiWHd6mv
HilU9qqkiOME8usLgXpXZwmIrcFHL/cVR1/QBgMURYd0v6JeS9++WLTgfih1tvBJ
uKR5QetFUE2F6AwlJt1/sxeIiY6tL4GyiJYTymydPbRqllv79JtmAak63HGBlY4p
GGyW7ONF6TuoMaWo++/bs+5HLLyksiTM1fwSx1iivdQGP/i9kgy2U1v6294XQIbR
FN5lZVxhXoIzSSR0wUclUiHUvzHh226UiMl78DxYNlOcPuDAdiq7cnXwsI0g70Qv
zvIw+zMQLK4k3K3gIWIDvVf/8PEiktncDJPcKsawRQuO2yKjqtSv7C7Zmy1pibiG
0+A8f9EbG9Kgjet9YEp37TzYs1yLbkh+2g0SZg1kEukRmCZZt1CF1clE7vvIRAyS
mQ3iWZGQu0bH2BEci5P0YqrnOy7bb6PEM2BzW6allblxRqRCyQX3+sDbtCxdUHWy
7yBnfxJy4CgQf9Hxi2GSKG1nBqVjYF2DroTi71ssO1EJl0A9rplkp+JR4rkw3gbE
JWgCillzq1rsvzMQ7tI1IZsmo/0hpjf1gq7TMaqlS5Lo3DbZEcTnfzyLliwpArNZ
ov4bT9y4c2VinqOD8pbf11QOpOgWC5EBfABzYa45GZqqbkTYFPVhGIbU5H+Y309h
RIxR92/aVeR213k6ISRl78/G03AssZc6T1L5JiypPrEhwitrixEBDYV5Ep3tuFj7
a4w3HsuBAPbDwT/w9U3JpKz10c+whRh1Vc7I9RYkl/t/T5SY6f8wEd85BV5h0nY3
3eEaiDiwx6NSi5rQ4apdYacA4bQ8qRvOgxYXkQiK5MI+3bXPh4xTI9cmnIelrBo4
DsWNGHwYFHV19ExpIy/FjeB1Wur+VEK7i+1JDLQMV1jB8RESNNJtltciC6J0itLa
PFsbn2xQkf8kbb8kc3pbPX5Sx/VilX+4GJMfTqkiAcVAm3jlRKBkzJGY09rWa+Av
YvpwlhNi/eDHFt/DowV7CQ9BACV48+GpSXB6T+vSjm3GMtSGBcGz5HYSzMZKmUFA
FDq27eoksKXnu6hki/3OvxobC3d5wa+8pcRGhaLJKhRQNArSCY55mPjeozmL8mD8
87knHtmmuxcI2wQPjghmcoBjGdE7Bx2bHFf31Fv3YDb7uYYmQy5emGbS5SlnAM44
ZqrIqhRzciF+OqsmrCxERf/pu5w+ka9GgFQyIy7cu7gtCQOiy76W6OL07Jie0gnq
lmZfj1TzVMezBeugBSUJXAsPkiOjW9eu+F1o3cFFgp+hfHXPToQq58Bqzr0jokq7
MPcE0sizKJWfC+D6nJ3Dbq7QAQwaFzCpNeFZC2rfpZfO26+4Mx1QG3kmzxqmTbSh
SP1qYjkXNPYdwBMz5Nv2AZWmgiTj7kDklMsSQFtPk1Lq+FVGVXKZEsBLpy2Wbb2A
1kZ9hDyzTYDE8YjvDBxTIjDraKXQuNWXwp9nZyrqC8XM/W9GS/QNJPRhAnRTutXu
pkhx1KG83vLUQYgv0YnbbmUPsdo2T0DinTNkJe4MqQhlfMr/x8GsME/1yiuZbI4A
pS857Kbr1gNQAxtJpdb/1BCWjiaCN62WS85Q3qREBBzYqYcEBYz3V/FLo9sK1oc3
1KPEv/IN7PjtRYbEKzxSqYekd1mBHHNMlAQtHMnic4G2hwVjeDj5tH3CmLMyn0of
p7E7/nmHHx3EKI8KYxeiQQoP4gVrJKm0OeSi5SmXygjoNCtzJjTypcvse1Hm60+h
KyLts0lVbxO8oYTCMuRbDifkK3x3CHzb3TlRE9ezwzX7WwmA5MZG6547CmsuntEY
PD9zkVkz5ukry5Xsf7eEIES9k9V/zniBihDz4hqn2W42jqOhLdGcP4tWwsOcWQmK
tg2ofLAoUSu4tUBlssf69OiPV4mraYhOGmNJzMAh1aHrxwAiumzpOyw6+JRcf/7C
RDeTHqGwI7gc/y+Og4OjbnbD+MI1M1+3BwgneTmmRMkWYYdnLvUqheDovj7cwmTU
YSi5XcbyOUPI+jkNurwtOQcpdegNnCfTSvItxzbuOMxrb0RmkKXGGIMVcUw+atq8
HCRwmhv4L3kKPtxZslgV3CbVvynUazqlzvGXCLA31mFnPTJsMXHVIVJUctNPpilN
efl4yDMvx2mBPp9sGxfoihOwYCR3wlmo2jC9x3OPZc2ZXvrYenufM3HJySvpz0Ed
bwhQ8ozByE8NfZojU4/Eegu2vGjZoXF4zdcUr+eGFGM7WkT471whOQP2Vm8RIWZl
9/fyH7xJ45WgOuOKWj3lPuJdr7VE4viDrG7eNc3Y2bD0GYUfgZxuURMdmkzzt5bJ
RCWdqt8FNvDr6bM9JEOm3cPqhWII3+IA92bNPY4Dl1jqI+A8WDH35XaCLuX927sD
NzuPWgGVx8HB6MoVZeHjjs4/coVWetiTyf0WZCuUkeTjJtUYLUzGjfbwpo65teuo
Xzhmwbx/HzNnczs7sWwjwmJ01hwgQIkq923H5SnyqzmTL58yBmwSZKfPdwJsNveb
ibJJ2JUlq6JKs1UfXCIWSXQ/ZEWP3QvNFlWqdG6BD32WkIPcibszKnG8eKdUVuj/
jUJItfEER4ujPFsQNgEt2KMceqNUIWsJ0ZRfwg2qhJ4wG1mr3ShyYqe4AxkxgBHb
Cg0Ii/xLjKqFpCfvb7/fi4N22zvSYYQTYemdJCLxg1ERavo3+WxPst8DbPDk/G/M
BY4qMTtGgy+3dZsY9ni99jRvJECUMuVy4oNNDd+CXRhO9LNslnWstQ/Y8lDictDa
0dXjxRSpvwTSiQ7HYa/jlShOvoluty3XpGyI58k4JMcrQ/C7nZs6WaoufA+cCf6S
5GoN38g8x32l5xtbNjeCdXju7o9B6o8hzrkEdj5OFESMMsT8wT+MSvsiORMRTrbp
HtFAduJpzmAALWgU/H9SP6SpAAvXdIcbfKTUAHV4bNjV9RGqIVUKoCQi0qaIKduT
ybDnSUnoQw9Cl0uGL4tG1SlU3b1tnXufjDg7Ry7knvtkDGQzjTT2t33SPhcbJs1Q
3qi5YGRih4rUZAaTV0Ft4NKQdz+w7NihdE9WSSVP/2BJOHVGMUeULcON/HUPFCuj
dBoK0pcUWy+5w0O/kT47VULBYe07nLuqEXii4S/4HQriYYFuB8sv5mjO8Qy91yVj
aerqO2KDj+LK1goYNPVF25sGpY5beOW29ixKPQ3iTpyY7cEPzzpzWTV1PjN3Dz5L
Oftq4LmnrGzEgPZIm3+EEU/19kv27tb4yoOisfIR9uGGlHQPMZXd9mA2xfLz+v6L
1HDV+hqODAfxrCt8ByDwg8Fud1YFlc6pkbAL5BdeH46scVf0jspkJdeywznF2GG/
JBsHpmQ8DQzYcHFVoQjhS39+eDgIiN1r1jv2taYDDtkEjFZp8HoyP3mOaR8ys+j7
zGcGJUtNvii1YQ7CJhHgcsH8GZzWMp3RcsY+OMYBx928a/oEtU0E9ForBFIc1f2z
rKRbKRZVBV3XjuRg7noQTG/cEoxgwSGPbdloRb4GRXF2GFrqA4vDdfJ2fsliWo7e
3Tl53uxV8R4ic/GfzFqqViQ27TB32BauYtAvaczrKtdkoCLjd0WeWa433RWyi7xY
Hr7SdZo2mYvP0K7U/CReUdq4TrFeDGAzlcVbgt+pjh5T7DKBjSeSLicQa7bMBL9E
DFrkeUxxeLwWylYcIu/ToUVnRvE3IALmwTTpidE4YnckJiJalG83CAPidtPupKfv
lQoiV3zFIv5vQ4yA+O5QoWg4pP/cNdlVuMHAqVx+sanVyLxXCc2hYTImBTuMvR1k
h/vZH8MVAH8a1npbEgff8NdncaAYkba5VDJbWmIwL/1EZFMiXbtj23xcfyGu6N/U
nU62AHoVbYj3RYITz2z7QZXG+cNUvjAqDk4/LEpBmPyOd5YZGvVivk5wryjeqkBN
VcxWlmc/0Z5KZGdXfAdq7m3YP0JNvJHfymRxsoE0nwzBo/CauGuinHJUhqKwtBRZ
gtHupVWnlUJMAPxkIDKvatBLVjA0QQT8/OmKuaVunXGpSb1L26otu2eAoksTocqO
0VE5Vi6Tn+dFYNmOU/xfnxyjcFrYFnJfB9F6bWwroAtlrTAuRUZLWgCp2nsAVw++
BF6e8wJVT+5NMBDuBAmKSJZ/p/pqfe437VCwweXvmAzU/NzaWt+tfd/uztaBOmoV
IU4YSib2HefqUPGTBezEi9kOTZR+2VtwAYy6HlJ8cq0ZEQDZv8xuE2414lFLPHi5
GlFLZ4W6mQ0IvaISZkDfddqG9AVtYCz12dF1f1Eue7xEUVM4Lg3IXbP+fXEpu21E
UF4eyYjrN34lYn2GNZJu2Wl4+x0KrXpoUUnlsNWDK0sUAafLXmI/YChyG4IvQ1xL
2Smc9fuA9uQzDA3nxtUQPz+SEewJSK7dF+TuqlrYsC4DMRLGquuARHAfvkY5S5j/
eD7b+KbZad11IB3milekPMgKNeqwYw0tuS/Nh1V9qI1IlIKZAn3h7gRvAkIjesSE
K/oTJdCN9z+Y3/OIhX2aA5Hv3l52gC7tvQpN4qiI/0B3bsersNQQ7v8IoR9YXXhN
PharHVHgZFcieBaviBeSl6yoIHsTvmGYDrzQbalyFhPxpl2vBVLkCLCZtHySx0BB
bq2ok4Zdy1Lj7E1CXUfKw5HO+2C6l43vD6sW9R9mrodKOqti0IAoFOeUcNCahBsS
UqLtNw0Aqjf6eHEWjGy/VwAC04L0N98Uo13BKg+K1T43JHR49WJbbM5B8gg5gxnh
PeKjg/H6cLiQCnLG0hVRpZsfJCnFetn7sHil09vpTa4NzHuLfydEF6vinxn7elC/
LFNAKf2jwInl8dBTCnXFPsmYOsQG+aSdUJNpTvlekR709LdqaLtIWBn4skqGfuE0
A0EDJHttRTt+y+G5890EcTeiqwNCljnZm9W1wBHdZR6mMOcmHUUSuHCINFehGIRA
SmcDsQIhyPFHNQYX5de5m3Or0pNhwBjaDuWXV8n9TK7XQW0kMIoaRzdPrpy5/Rjm
mfl0T+ikcBc8+fTt7jgD/FDjwU1AR+KB6UelwmrZCjHg3R01rJa9hrYBcWu1VjIw
ZWIVlEwzoXzS5S0Pb2zJ6At5bPzuxc949bVkbinOVa6AzlW5LjCzkuBKCJJ0SV06
R+KG1geCL3IL42opL5pQzxO+mYyG0zBtljAN6XQqFeUQrDxsAkbDYcKaOY5Ptx8c
lLV8eBoc0zToNPmaFev4Wx2jAXkngB6By8eE29wtbYJo3qOVB0yrPt3MT/qFGiFA
DBOQYnPp5ItCHdefRdJzHXTSe9N8IE07kPj9dbXF5ZfSL5kJv+UblVa6lDRmEP0G
9elnn/s8J6CaMJcKGc9KoqFaS3EtqVXMa0PkFioG0MunnM0CTAkmmJBxeWY1yj6R
PpTrdMkqgMGAyiXLfWI5bDRzyWt/sQDiERLkNzk8GMuT0765rtknNMevBRPqY1z7
1cXQkbDFl2aaKF7QDgymmcZIt4A3ANdPt2e8nOeV3gXGACNgy3GXWphu4Kt5Ej+m
BtJhqZ+V3SnuPwNG/AImaZIlLHfemUp1kM0QdJmg79zSAPGz2c68mMgwAb9Ehe7G
96w1nIQ427oqsboMM7Vh5f8qsjThxRwl4eeSu+cOBmSiwSuzMV6ZNLd9IdQaLpV+
z5HiaTTCvO1ln9HlTZlB9Q69HzU5wfbD7SyCL0hXNkspgwqCHfq2k8IPvVhSJH+q
HR8L5HJRvTtun0AWLFrZOK7Awm/N17Zwdxz8DBflkkGxVcsoaB9wdyXmu1X6T3CL
UOyAwMx5dXV6f1dyb1zBw/8GZeJ1RIiBE1H7prxz3SsDUTAeNXZY59y3ZSs2ilOg
x/kXCFNRsc4ZP7mLGdbJxLTNHHOjne2RThD026dnKRiUo6uiiKwONixg4WYXSGpI
wx6luPdoTlg3pkUWle4dJ16b+kQXvL540UM/csvqWevil+3gMem4whfZy146pRHt
IWv/CrBonXKFq/SjRCw/QVTBoOm9hyk55QilYTwT77v0iyw3wao0aJmAfh/9Mh+b
OgL8mfDHjCcGECAvDIzVHb0T2nhTiSQwXR9zhvxJJH0EdnJi/lF5B4DIUf95+oY+
9YIsQxEvCVyYhLnWSg0rjxIISyzT0oZairwmb3DLJRaMznR5S7NFFpeNMNaYABuf
uRAfaYj+V956l39XUHNS9ZR/F+jmqNB+FNHLi6D7n7AFEZrh2ie2UCZmGfA/IOqZ
osFwwg4ET+x80qVE5qPNPA+erfbUAz7txO2OWqihW64BZ0mgPlqu1bRfM/iv1czz
legitwfjc30/ORKyrq0X11SZvpDrNfODJxFuDHNOaLckefeoPJ7I4R9hHb5aBlaL
CAXxi0Q5NHoH1fVXLbvkwpMkT5mXSbVOgA20CDK8zdjEpQ1ALzgRtQqJRb7kuLr1
W+AxA/4jJ3VIqE7tjyXVBYoCj1pQvZ+DpXN5gTa/yz8QShKIs5f+hWrPlj3D+0U7
2ZnbGp8HZmQdpXwv4CrsOGAI9oIc9GVUd5oUOegniplF+PdNLKvKmtJPaXnPn+g1
Xr/qqIiE5PdQG2rKCg8N//9uGhE4q7S4wIxmYctU1WM4sXnRHudTLfymEF94Opb4
ArbkTW8D2NSPYBfTg8nk0fTuBsbuh0dm7mDGD2WnUT1fSJObZCd928nVwCvEh1Sq
Bv8N3sUhOVRBhqGxpHjDLRO9IQ6vIWtcMRma0T0OcdC7XoG86hVcNDRlUbc5dPtc
j+CeNhAKzCOGNy4tV4maHptK6B4yw1BSDnoM9X4In1KkHyt3vKi7gZqUUpfE6g6Y
2bsgR/458Dme+jV8wNS4fcWlu4OFSvzIqriizpTVGae1SB/V/JYDFjsT+Z6kxm4Z
WRS166ZoHPyD69MgsEVscgVvm08cH+EXYXo3Cofbj8LNTVV1/yzcsUFUpwtGIJCe
mXZ8seYLyFcTDkJM7rxDpCZd+8v3vD/y4ZP5Z0oFSBeBEcYzWpujqiELrm7+C5r5
np3sAh1Hd9Sr/hh8+VpDoMJbZqfhvA7GWriXeEY4asI7q7rHDJvpmP/gFmMX6MtL
uY3GZV/xTMLxbkrDLhdEHgItTGBsPjbgp8zIV0YSTG63pYEg3zC/QuD0TZOlRDQN
KAQccBD7Fmh2GxG7YqpNlciGVjCshGvpwCbTcX3W18hexAInp5a7z2dX+vmxpHRR
qFjm2zmKVAiFP1oPR5LeBw==
`protect END_PROTECTED
