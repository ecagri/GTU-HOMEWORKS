`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q2pGkiI+3elSGeqWSwvFt8I0rHioPMQM2Wj6bgZq1edZi9strCXo4oFoA00rusOu
04T7hFFm6Y58xSkC5nw9UMg/qwyuysjNMjOf2AduJXalSgZVKXnDVqkmqBzFVB47
04lNrzShGycn/MtHbRXd8IzT6Q7mn5pN6k9NqJFrXXCqRfAYhEHwtFGUKohSWMNu
7RRg8bxco4aAXbgyLWiaBxNRVUYfJ4dD6L5MieL6jMt5iWggdjoHaMmaKz4HfV+X
wKnwA3Uj6kss8VNky9/c0Q8WozGAzgjdGzJFD8GiaRepgulZyLbXNMKq4o1hVdpO
xpeHCSSoL0qJY1p70HoWy1NvdT4GWyT2tsXgjtSAi+TnPNDd+0KH7qZd8bdZn7PD
4/HcmfEn1HmYgTHDyMRHsWMyEd2u2l2eYQCg9FJ+R+L03mDEtfQmeigQcq2u4QgO
QqTKIBH7SHqkhsxS6FNm5o6Bo5xfdmfIMdlXWAzQjH+ilPQy7EpenfWp7Kx5g/XR
0T2DciEcVFVV+lhCiToIXwOqHmscKSGU1FJJVZZts7ufOnks84bIzxweVs76XGaD
YKlYJF0Mi0v0UaIzgdk7bvpaGDnlUMz9tCV4qoHWvPogYXOswhrN2XBfrpbn3bIQ
IV2+B6zgIRPoB0koXzZfAocMAL6SjLp2qDQjzt6s3Arm4t3AsnxllQKUtJGWszsT
/o14ahjFYIJDZ6/IqN4nuHAq2QpJLdL3YzDLha6qNPGFktD2FTPHKi0HytDNKTty
deFPXMyXxl8h+F1ursrshJMf+eMiDehSIfyAI4JaI02kOVJl89dglHbBhvfurkfp
KHxyW/cDCl1b6rVjtN0z8N4XQ+NmyeHymTXTuObkiVdUHxclPdzS9RGIGf8TtRsa
NwREeus/0CjAkYAA4g0T0a0CG251tvVYU5AmEgJswci29VCrzSKOzISKCRRoVWJe
yhl8EaCpQPhZOW1DEHXrJvYlVle8vEuSKLZCiyfq8/UGcM7JnKjNG6T/z9mQNBTq
CwTTBtp+JRI7EyCqgs34QI9ItVFuCPr8HeiPWxHntU+YTjhpNwVEEchhDXy3pUy6
Rbn35cxBu0vf4gzfSlHC4CoNQI66J9/x9NCGYHnIBpyV6PuHVUE1vy9T2MmRr/pI
g1zylOsS9YKV1ovW/nq+U/2Wu6N/6Ftqh+u+3rTTmUYhu75KiXDt4/lCveL7Nrrx
JrAlO01fWC1OQtZ1WiyiqfC8zGeobG/cHDXkOjWQMfsu1cTQRJoVIYTi4tsISJwi
dP0Fk2VAHBJwBLSRqATKOvS4mPech0SKyn+BeaHSI1kCRerTMztF/T7khtaAuvzu
qDHGfSgjkf7hD+ChA2G8FIPxcsZeuH4iNHSqYCkwyohjy1wAUkRlj1C9p/cExcdx
EeAkuoznmR027o/w3vA8nLxk+g1+3lMoXfDQ0cXjN7ke9abIzOyo7fmL4ZdXohle
slYjWQEr0u4fJV0LGpdH1CMQ7VhZyrCbtDv44WEK8hxdSxXzkGiZtyUszPw9A/Xf
b2W+iEHkRD7y7vZBZsaekjC2+hCapVau8FPE2Xnuv+wgmpPUvgS45JvfwYmhS4uo
/4x+k12ATvsBunbAa8F0Rk2E6/1dNhbZP026FQs4kKnI0WKaKbliPNeNs3iMV8GV
e14i42Lhb6VFUKlMScsg9ByF04ZVAw3EWNM/T0+ZbAurwdSmHJj6KoDf1/aj55xC
l+HKkv2nLO+MWhQ1iVRSkZPuThZEujQMf1WRVsZVLFjgPjlh8zD/xVE0mVy9Id2/
bpvnjkEmnAPpNsVhnmTQZzlOml1KFep0jOS2uucVNoT/nnUJ4Kkvv3ggLWIW11x2
lCswXj1FgoyXFXZycHEpcnFW4OV3KEXOCdFDDWWjBA50UAYdstyv1JF8JdtGPvnx
gumRFHFwpgYAaFxszj0M1WnWEz19BuqWUiBe91GZvEip1yhMvi2+cn/vrkl2idNO
QsRTHJ8+lSQ3jX/DoNDlETCOlGLOwqNuUdIyScYVTTcmgbGa0Az6R/s2UyBjMJ1+
pD7HhuB04s7NjRg97cfsxDiYV0dzKdmtlv/bwkbcgZKmaQX4232tgjbCCvgTJkxk
a0ni3l+kfSEBMwia92PiyWtqkOV5qPv6G0zImpHJdtm3ZdLIsZGezKcISJuFHglx
TDcHDgVE/0mssF6Tb/fWRxosdChuUcdUykX6g7u8SltFwEsINyJswBfsB3m395e2
g+lbw+xal42ATXu1YEQv3r6kGp3AHRPEW6lDOj4wdLsNG700loqELV2vl7qlsW+S
mYIXSSby0wmS4623fezsNWgMpAgTXm02NO6l1+/9bpNw/mpQ/+05yxap+QZqiGzg
FeROL1+HNrkp4/fkMgQtXQk/AwvHkTktuJ8t/MFDYN7N/KiadCGIK7ucqIzzeTYy
OYfhVfNE/AtudofKWO+JclbUOwPqr6sIk9zfEWo5yKnMp84IEv8d5sbRWP42fGbY
bWL8IdrhG5SDAvVdXXkCPh0kYfX6F9U6UNmmKJnClXEVcwwdV1x+ZCPeUKdhwuWI
uUOQQRdAoBkpJeA/aYG5ScAtBoThaQJhmabv9o74XBKEKNmFrbDOgLP/aomZLKHh
3P18Nu+pRKnsZfaNHmngZ8/DuSrbtGJv/JwRYDzb2wVGG6QWGhPHEQCJQQtyAjjG
v5n774rUdGDTHJoqhIIATRbzhz2ii+yvObw2NNXYvWiGNuih5qWc4knCpGc4kYq3
f43iEvDCexKCcAreh6dZXMABfw+q2yAqYNqga2t00/QGqbOv7QQ+mHXDGxGVSiJm
uGZEkMfjo00ASScF+m5WTq8Gy0nuA3j154/FTyFL0uCXsOzpE89AgWxCQinoAoED
wUJWCZ+fFmYs7eErBOeTvjCeZdm7FVC7NqAYmGNx95TpukV5FGhEGyUr4QRcJcie
nlu+LpdPQzfjtgVgphxss+ZxZ9arwFz/rzdFCMxHgCE9QWDI0mrr/h23ftyrP1tq
e79JFX3KQNXjAX7rias2tFvJF9z+MPfICSFEKAaQaYZxtXY+wOONopEufQwCNioX
Rx2pJlrCQku+xK/nbKHscx/kSOoEk5Hi0kGDPiXWvyQRxAX+1c6YKJeb3Yw1GG36
LjiY+v49qtym82sukAm4hmhGYbnMucRV+Ts/QFbqjibHdTlRbVvnHosaNFyC6LOh
wm3UVbfxNHZriZqdgU5BAgwSRvleMq7mVZLpu5EPqFEaEVAP11ufOVdlp+nEIXPx
kVzcULJjKJclBjCkaRIrq5efgGmtsxR6Ry9leRq19FmT+BZsqd6K8x09BucxhtIm
Fh6df34frBHYluHNtcAbvj5eIBU27Z+xTB7sAmwWWEoLfXarALOOooQozSAmHRX8
ZbyjbUok1T5pwuXEtO8dDvsSTwy9zo9VWIQbWsNLHt+A0cWywcSWHHdEZ2mhIS0h
6+qg314tuH5QwgsDHnM6L5MVcxSLNvxga7SIvOObWzthZV4OZapLy4sUAY4YRO/L
PfUhJgvnFu7bNfYSq+5Keq+W2ppDOaPVuGJ33vvjJ/PoOiBb6K6BrZ0nF33iVpW2
aUkyPn9Q2zxBGC1RkYBmlwh2ZhRbs1qkkpo6Ri36If+0o7SJfqO0bc/rBrF72bWM
L//2+cgjCHqepfMqs1/1qTkFYkmbewZnA8fmqhL1uIshA8kit/mxvfCNP7rgRmdP
QeY7u/alcAwOiDBAOzbmUGvQ9QDqYEhMoH/4Cy9MzsEVorw1Jd2nQGl3XF2hZY0v
++kzCUdwF14arVGemGLKBO+OLcOBRCL0KgjiJ/jsVXgA6AhG4fyZp3mw80dWNxmq
0CnoMFm5tChpYqGMyPvjDxQsRDu2aLf0GxI07+pUFvzxo6YU21oSwQEFwkNn6Giu
zj4oK9xSZwijKt/Z9UdSxNFOolxaGmppWGpevNkC57+VXCyffqwqVzQg/1WSgAbd
oaUKwdjmSdCZzX2ebgHm9mCNrmuBKuOSbEY3qhC2k93iJBhAoONHFlFL7aY63xml
o0dkiEOhmCYS5RDOxwAAfEBmJJzN3Hen+7ID55gidvf2f3M4O5NfcXVVxKrZk38B
XrNVScJNVDcPUThUK7W9dPx86e9A3vo6dlBQ9JPgOiEwHoZDXD9g6ml+E1QHvdCe
CzIq+07n5IL/JBxU3NrY5515dSdZ9U+xjagT4p7IM67HjfeMTLQtwghFgSM6e2/t
rBoMKEyKHYuMdgtc4PR0CUIxWnjPewOcHRQF7J2eOPbMlXdTERX92KUmps/7Ov21
BLF/OncH2k7kaj/XSsf0TF+0PlJ6FpNqnCQr4+MfZ3Pso6sgjFjB622bEG9dqsC9
sYwkjJgZ1EUMpREqUQK1W2PnRRR5UFPVRsJjn0n2i06W0/4hYMXF2FZnJNbFYiyJ
uXuG1zZ7XLDQV3AyseQtX0NdyYtS3m2+V4Fdrv+uO6/mEQuz9B6gwsxl0Q2O2TCt
mlBepjn+ksJpsJLoeJNhbHSQD/pjewZQYqy04nazhuVqqjou8oNtpmdrCXcrWOr1
See9+aiHSw4M8NeWUhRl8eDXPENoV4zth2piqc36gHUiW5CjQvadKrLdKV0juHQT
GNtiwA18zOBOqlI8eEIUDNINb6/tOrYBLccGQoPfRAxF70X37gG4RgiYErSsc7vS
TXYYkE7Z6l0/JBqTzW5yQQS9Ty20BgyUgaaFViHw0mnfKSpL0LFCC27BBRR7jm8C
2e5LGb5UIbjpZXJMpkYWFY1Mp27uKLd4jDqWtpNHewaQY4eBBN33jPY1txzpC0ZH
o9jnaaahUMX7GWhYH7vmlV7ofiJflAwuHHwHQuAErGb9ECNsmS7vcWgfrh07bKBb
2ojUs6nYzmClTQCSv6rqbEV0ObIF1v8qfYS0aFBphbYYnfWV6/+WeJI7jTShxqtv
qoIWQj15usPeN/YqfZHQd+hXgof43edxtrDGboV03u7RonPLKY7xB+b5B2v4crXI
dgCJpRcrWuiMpTmLkUYDACXnXVWKcOFRot3PdC6Qox73RkJsyY8FePagYF3lenPh
U25MnYHTfc64/aPaTQmfhd5IAohKw4PY19wouhi/yydcF03djIIyoEppkvs14hyH
ybJPMvNKR0urFgqQQgudGFkeMLyaEo/I8xzFdaVOSFT1xMgWTIt83bKfMnGntPYA
3jTTKBMCDHmcfUXK7sfg8nwR54+oZQhDIAKPDst1gyfz5JZFT//rPvvCsXlAWL6+
1mKdqJ9/bJD06FDQi4FcNMFCEVQxiMG0+e4c0sppqkR2m42KNm+jW+geXGdvLR66
pYK7eussZpMBoerEZJ5b0l8KySjblFy9PS53GvN3G7Id7309zcM46MkSo2D3nT2B
kZXvwFKH4eQdFJmt3m5sEFbDYgkFxyPS7Ryw3w40F6p1VCoAC8C/hV7LSmYU9zqX
HZcQ+0gAOxiEGQl216GFxwJllN43rjB240UWcSV4USP0Moc2GBg1YEGTr+/Sktau
ItI8+/8U4Bne+0Ju56AEaDkszN6Sk6kef+II6QvJUgMCPbXpMy9mTjFqzW2W35ba
SmTF6gCugEQq5mgYkXTt5W+2wg02GjcAXL7lTEkupaLKNl8rL2Tv4e1Hkiys/0S5
izEwo3yB/OlFzE/oKmVj8CMwUVHdbh5De0gUNNJzM/xFY0RtlMExuSka/uRuzkCI
dI9hZ2WhQC/oYZlH/uUTWjeSRhk8822jkjxXSnyXAREOzYO9oXtF1EeefD+a2Ssl
psZWsHGT0TqJRREGHKrz8XKoL3ydookfbcPAJPWO5E8kzSAzYDpH1d8390IHa866
ppiVnPAjiamZG2Pilp5yZ2FhCoVSbSWRu0vT9z5BPFq+9PJOOkCu9eNPc12WWcBL
vDqlEGs/MXbtWU1XQAIpuk1GCs8/Ripcigsj2ItonFB8TNIIk/5SnT6j6LkwUImC
f51tnakHAOTnE+d4Zc3+Nnu3X90OcC05WLaYK4VIjXGUWRn7dqIH18O3MXvK5bN7
dfhWe7vYgbQkkxdRmLqlrh598HOI8DPREisR3t7Y+FLdz0wbw3q4VLd6FensnZ5x
EHn4ggPWPcSdSiTMh3Qd3YNrDj9vAqS/f/MhWzXKTvsCMSAqDEAsNg87QLH92W8X
lei1FOD+nNH7DpeQ011KG2Xd+koKyxkC8GTjo0mPeCL23mnc/6H5P3cM79deV9TX
wHto4CwBRLnpiuKQSIEkDdaK72FqgJLf+JqUDsaQL2ojdi2Ue8LpHhR8f4ccz96M
u/3OIq2xmfhiAmS+ViYnsM9HROqBWRmGGTVYYZFFVGKFBGmPxJREoP2KNM9EfRJ5
iwZf+TuztGzW0ldVQy68y+fYxROxEvgqJHDQAHRNjR5Vg4lGJs78m8+sZs00rlJn
frqCQdz2L6+B3mKy2vuTsu/I7rkW18zjDOrK8VUH+wU9zZ2tfpQ2WVxmGPj/uVXG
ccr1pGqWg+WqtWc67R9pW9trEnl2nikUyDGRjYZ4lVcB8Giae5S7l6xf0O0hnwIE
8H79qCdzlB/HYrn5SM8M2bSYR6DLBJKqvx1Q2CY/oGvoNFoj69RJ3DdwN4Nk3WaT
Lui3TsnHtMXyz/jfL5KfemGXOBCRRt4UiupEf5du0NrHbzs7lOBrMbLefyRt0Ava
Gq/HpYarcXnhynR47rYJoX/i4gRngY4YsTfkJ4G/PR+4kNIIYYmBhFmYncO6Omkf
Vqu7+7nFX0vQnCov1dIrtKCzIIkwD9CaVz73TmwvCp7Za/LQU4kD12NQRQIWgEIY
diCWyjpcj99UBP6dGnFuiFdjMDfZ4IDAM1uaxtONllSoScuR0deZv5UCnjq50a8+
YuV5PqHcIqlMNrWXgY+16DRBzunnUQXCp7i7tKEPQmuPJssZ7g66Cg1K6SwlCpY/
tc52qYwnHHkZNggFXaguTGJ87yClTC34zyAetYy5f1+KH7NPRY31T0g9L5Kde/3u
FRiok5YMrtRxS7ngxJ1BdHyVfB5j7P9Oujp6NTgaBQOm0sS/8v6kdT/kPc4Wfty2
DpcoOWtYwPKFrVKuCA+Lpl5Am8QeEhzWR0bZCbARH3U/fbb3ox5irmPKlA3LrWHP
sgKda3jgJaIXV4yv677XcxCFHCkaQVOtwE9fl0irojFHuhfEcTuKopzlaBDyFoFB
RgjBW2T+Hq9bZOKIW7OCDZ064VgWbMaetHLG2CykllTsEQfQbTBdX4nYBDMXwz8h
g+IgE66XOAc5tqObK1ZGCIBmde7r06JU7GxfQTT7k+PSjZaHbrbvfm+zD5ISOoEK
kGP5PAgWct9+Y7zCkUFXexwKTBi1B36zpIgB9JBxnYDMYYycxTJP+U1pqc4VaFMb
TihSLd+e9kpyhVFeDdsfYD34iXUHkHEvWwDZy2+F4evkt7x1MZTL24BE7FpT1tJS
wNLyAuvdN0GCNzEhEVbRPhkBAyTjupLqBBFQrN10L3liaHvSn6/Yu3XDZAZXdKbK
yAgZ6zqiH8KCElDbz7Jm4OGeTmCFOCY1XnrusWbxJ3Wro5+0+Mhpp6anKvcnY4GV
6KtEus7qD0iMLEbvPPEEc0VXs6gQyybtVz7m/b608Cilv5u9U3zFh4JqjKtvl8FS
OkHrkPrBsAnhOfiKv05hzoyigqFQzfJUdZNGJDM2llhOtfxxH7crVUr9+5g6gpc5
cNixygTiFwELrWCl3fdlUIa1PwkA5Me3ODtaYdnwM1q54wmttWIZKNdq+9V3/5Lx
jbZfajjIWHRmIPbckJXTOVK+BcmpC661GY8U5H12WsmBhHOvaNqpzC6n6td9siGk
fa7khkzZmL2rTvqLooKgvPin2eXOscl0WuhXThhM5c7DKjjzRjrDbQDtz96WcZx7
IjhRT4V5QxBfQNC6/sMHwnUKg/VEnsaiV5dOZpvvTYIYPx8fDeDRTlvvHiy+Poiw
TBuhpB8FFYrq5Lg8t3UQLfWuwP3J1k3Uv+mhSyoGZEJ3FVwzX5H06ZNoKb5vjSnp
6h/sqO9RUUwJ+W4RhZi4BQR/1Nl7xztnUJ7bHrI8MSp2DTequOAAFOGU6e18KgvD
OpICMJdAMDaZfqjN2l/Jou5YWKroiW929HUO/omAiDernL6yZ/0V6QbqFkg9ql03
cMgz6FXWgphFVAzldef7Lb6HniMzJMwmDPgjIezbvTMVjQuCCVlHOfX2NFypYwsP
uN2YdkZjOdKGQlZmJWD2J9AfPMDciNGE/uaO1uLD8prSCf18xkvfmTkCnaXs4goZ
HlH5ndI/oQwt8BJr+J0/7qtkSObrhPjjU37MZiaz4uDaSdZSMS4VJKe5MMNy4+71
xuKgdT7hwYSMN/wMIkSYQqA/xj+tBWX/9Wzyb4WnhUa85gvCFP2UYySM2Kd3eahG
vMHFlo2B9599pH3zTEgu5vutwGlAIUptgZ95pC7e/GJumj0xM9rIVfaFejo4gNko
Pd50aH28VLIydY1hE6Xmuh8RwRBf5Tzpw70wiKEQW2/0HGOcnKv0vWNCQuWCYejm
X8o/EttquWADlax5Am5ov22/BonJ50XJoCqWQ8Alrs5KACdxxjeR96uAgT/swbk1
h9HYCbrQBdrXWZ+tutO+eHYTHp5cGwwR9WApvt7LpyWR1/0wiF+Gj+rWcX8a8dyy
8e3szffLfhYf2VOjxIK4gK8K8DYEgEcz8cPs3vgHVVLl9aN2D+H2kwWDmeLSLHjr
BNnyaWG2PQlu7pUUtoQ+ow6rylp8lXd4mrfQ5sudW4KrSqa/qDKLliyD9ELLBI5e
tMIpbSciDlm8klKABcVhcqF/t2+uKHiSSmE6flOe/Br71vrN/YxRmysOSwkAFDvE
wDE5lya9838640q0k+Kvt/NiKDZBkEfoCqOo8i87ISM53/DVyH41IiZScoQqyn7F
v1d+WeFjYtIfuJoP4Y4QG4d/iERJ18q5FoopJhqhhDxIWiEOWtZjxhSwjbAKy7+7
5/xEdNk652pQL1n4tmHp8v7KXL8BcH2D4KTFcf9PtAogSWipbXI1rOov24YzOrRC
4qcwnPcQ2l+QkCUA5x8KesX72h8ZBuMTMiqdkdxaLUwOk0Z33V9qy8iqR5fR4pn4
dgHt4mYQV/lJS2gbbxHdVl8y+w6yMX2bKFRluiyEZw25mQxl0HidunmDLT+opXR0
Db4Br6ZLlnRY7/xsGIRDvS+NDnd+elRMOoFo2mEaOfFUyIfr7/N7Yu262E/6Acz6
vH6pSs6wfUFyYQg5BUk3dnUDFTm3Wry79O5NymZvkqizTdy905MGWVOx0RzCxJlc
Gi4uokkQ4exGnzJ9EAmMfKkWQg8HZ1oQOKXeXIj/lFYxAi7MdtZqkZHpp81NEwEU
9uE3FusFAlBAh4SO8y6fknCmW8OOgtO/tjj3E6WP0EIvOum/IslQ6Vwv/AsvQlPj
YOoBXlXGYuzpcvkNE1yp7S1rvKjo/LzoV4Idj90mS7DHw4a8/YEGW2zUVXKF4fPl
VmNHpw0rSz6cXHqpNVmp1t1B0Tg71BvqB+2+bDoAzm20rDuJ+LMqe4sLsaJrfhHT
URPTYVFBTFdLkZf+Yz2LiPY6jqtCY/Of+qypmDctb4KAC8l0nwqIOUcAbZm/0+0b
EKUQ6R6zd17UzUTWz72dFTU6FrgyFb7q/3+/I8B+CfTnCP4truZWNloZZx5r3FAY
zFnIp6cB5EQejS0ureZfjyu8IC9Wr1lrhdwlLh4K0+qFa3ehERq3KFb2TcTpA0zJ
rnk2kdvVspTrIoiwXF7cyzUywJlsRbUICGUtjoxGuVzqWJrA63l1dhyftRw5IU19
N6jI/UyAq5lYSu1CV8IuLcOpU3IpnMn2jQQxlH734LiIP7VsFmfuCqk5vjdBhWFS
5uyc3w0lUCVPtLeeWtCk52bOvH178+IJQeE2M4q+6Keah/4teBim6CL+WeKkI9YM
D8ZBpkFN0Gwqp+Xq7JrsVDRsiZX7SybwCp2YjMdiP/d8jMIFOP93+ggPiL7yrGf5
CYnVEjYVd31AS7WrymYtDeUjjXNPWUzxd6UhcWYsSpovZD6YRVYhIAlYZLIkJTFX
QzuUdxTrX3NP44+BOFwub14eyacW1kDniJ0hyzfrrnlgsPj+vf4PGpG61FoXnDTC
EJcSwYIZZyF5iHQAXrKIz+dQeof30QKvpZjxDzRF2NFUNY/ffhC/xaOQV/VX/Z4/
yiHxB9hvOi0hgezmYbjfTweNcbtSaoRlRl/WqIUOVRHZ/XLMmwlt1DfZU9qZdWwR
qzUxKh7oek3oKoL0nRenEc6nMJoBrMLYhNTRmSMkvsid7C8sQAODEUx+zsZMOU/S
sJpdUK7/Lf8EqltXDDqIF27RrQuq2kZ3D02UlJDLuCV1oxZqYMcOqO4jtdpqJgma
3CcS1YGur7Xejeai77h77OIKHDyVP7W8P6VGLL9zHZ+0cO58BQP1IFwsDBUXaZGN
k1nG7cZ61opfgRBE/A+s6g2QXDiQH56TmtOFLcFkKjfrYHLAaw+fTdRf/MY7rpHD
XwfCnAQ+9MbD//dJ/0Ao4V6XRuyAzJMK8q6//Ovb3JeLiVqHuHW7A/tMIgE19XSH
MaqK+Mh9Sg6hQjwgkn5n5dnk1e/LQzK1dbIJTwtvDW52urIh3u0FBd2xKVBB1Xvz
KbvY6sbSiwg2lKkbuanW1ifyikQeRo7rSaXC3C4om8LY4iIjHxJSMr2SO42ry7NX
cAG+NG2sTMz7tsM2ILz28MPICbcSX6iaIodtSWTc/706/r2nhVdK4mRG9YiSvGc8
AcTqj5Eof0eQr2dGTLnPEKmOYStcAsrfrRQrGU0b3BXrgVE8PTZm+tTomT9cjW9B
jlGkJephVDgLay4JrXNqZQo+Y7yVYgHEycPkMsUXaOMRS+FjqQB5F9WznJUTrrlJ
PGd/EZfN4hlCZk64fs+WpKNa964/Qo3LwC9US9KLbgqGtxdmJ3yJNYQ+Ii/ArnJb
6rOIjUlqLCgJayGdzsFGifkJTDtXqp9cSmPgdnxqn3P7fXweV29D5RXG7pK40uAh
6yA1N+0SnPzgNXELSTfa0tmmMSL/6Jj2FKBTb6AfQgx/VY+bBkTzZ0k56q+uYy5E
uBfN6JuJe8TkmxrCvgreFH4evG5mnsna5OVc2Fh+jwB/1oCmjp6GeigEHwnce6NF
UO5tSpQgkQIe281IB6KlCI6djeF3P29KS/LsCPVPDhnYUs31bEAeQUdVZgf/xLbf
ef72CMLyPCCWuMIhWAGddHjDgVDzFqE4EC7vPVDll1ODf1f0gw7qhyhVPjjU9Hvs
qIqvVGN+QCJrH+Zaptti5u3m8tVW+Pbqn2A88n1Kado5Wm53NcpGaw6rZfe1PmPT
bj5iCFJzN4Rbgwo3PoOt35qxL8MgDKH5wK9KDKEc/2v5PhN/bf4az97n4gL/1bQ9
K613+h2K+6HUVAZHds/HFC7sHGSNqV8gIe0IOq4zUb4S+QnxNuflA66lDWkUTn6w
rEfNWBD09LcjsS+USvIHczS8i8iC7P+n8QZ0IbdBWAdA43MOpJ3Bt9GSwQLp2vyM
QOBPMfkjK2lByqywM8r7W+mzRMG7nJQUtHt7RVb25a90bnVl1kcUkXN6emFgWldf
1z2lTVMZ9wrKDg6NX5B52Jvk9XcP1q7vfstbrezRK5CMUuQhT9KHZG2l9q4LpWd3
oyQamD8FN+Sl9ld3I19/KURAQl3dnr+nS3PJpwwpx4LlI+k9QBvDe4IpUDGL/ZG6
sdDkZjaKoUpC6eKXFIDWmCXj9SaU/gJ5Y/PTrEkKTOBNgqr+xGqt//RF1uGQsB/C
q4c4mLeZyrbVdATO+Ij7xg3dUf+Ldc6knyBluZ7DF5dcFnT+9nGwW+yyC4HNl4Ez
MZxZUid+AIH9v+jlYFsMs9geN4WgIFNxV2cv3N2vbCXpOMeKGmZU2ZDb5MB0DmED
OeTc96t4Dx/14DbD3TFyoIQvCwWt8XxRDPd1DH3GorWiT8OR/jo7AcG7XCcoLmQ4
AIqkmjNoU75QDe2ifhpkUQ8pHNKA4r7twXjbFEyU6dsM3ejd8D0eEhSn2+ZKH+bF
wOZ25lONYdxdOdCFsiynsCGKRE8rsmsUl5d8KeyaHeV89yJKMxN7eEFmlLrV04mh
3vS7ZulhX8FgAxz1ZzgYVfyQeeTHIre3Cg0/JSl/ciz6ORzwDNZ1SHPXxIJaJytZ
GyhdryMzZFrI4C4DGMy/tcIzoHhxkp08nH2dpbNTq/RtkUyiiC7kW8iOE2R874lZ
BnEpduf/Rxd1RGymMN5TBcooSIxd95I83SWH7XpBJ19mbHi92GDBFNBqkeIAnfjO
JdrK++wdn9pHEkDhCNF1AHWdABFWUAQPgVtgxgfJp5l0rnF2ymGmLhnOpy1+gBif
m4+CBOIX8vK5MILqcVSOQsOMQC4CzjGe/v7Q/XiX7vRZu+grCBhG7WieE0+80Zsz
mQOzxi6W97gXnPC8CywmwXCrSD1Nae6HX6x8fFDZqKzcurWZ0TJx6ueRZO2fHgaz
cHIID+gQD4hNjOoQmjr52o/Ca+exPHgX7kN/vL/Z4I7VIDbQ0J4rtNVU1xBeXVHW
Ryrvn266EeLYV7FXTjYIa5z+wzdDVP1Gj3W+0JuJsphIRAJcH8r4WoyPniF9u01D
fu1ufAbj10VbfZQR8up1VfWMGi9nTAjzSTmxQZmS/LUIa4v2p4gWwRpvjFI/q4IU
g1fDroBnEgcpPvp8ghjyj5pkbCSRxNL7ClDc7wXoBiufzPbGbIyw/6XLFYas4ica
T+yTtrQ4lVQNhzqGdVBlBWFOnG+1adaTBXuXEhC6jLMWP6HDW5PzEZn7vjMIr/Pk
zx8crWMoY6jCU+tArdKRxroZnaUbN7O5KI2ZkKwwRN4l20m/wqhZJKW5ggWSaebX
Tsq5L1cv5t4+Fbiito6T7izQ3f4wlI+W7S1pi308xy0sFUWKK0ZypUWDm2RTL/p8
szVZWnbhkJRUFoqH0lo3m5jffG+PQcm3By4+d4T7OeppKCEWzEvRgpHWJJYHCJ5/
jeUXn+wP0RNxiaLlpazT2gv/BnUTzeX639gL6eA/X+DaFMSfSTUqUh8KCtvFCzlC
k20PaSpCMpuBQ+orQ1ebuEN2LNlv59TcBNrYw2uSdocoqd6o2Qov29YxhtCBXLWo
LTfqlva7VorkQOatiwdh3IwgeJ0rieVs6znTcrUzsiWZzncsWtJ4yjpQhZcXXVo2
dBghUyl5WrZQdw4WkVK+TJ2cgKm5Fc7BByAZv9Q94fLwvHW1q3G/cq+pMv7BMBbc
QM8cw6vEMd9Z7nrstlPQbjIoYPmbMw+H7W9bAouVGEO6hVwtKloK8esyTUMg0cRl
Jpu1mhJZ+ymfnGhkJWb2QdLN2kepcIosW6oDFV+rBdASMF/tayio/hW3adTbsoQ5
B6Nyw4bbm5XYB2p5BJLULvaxA8WTJoPWmjWDan7QCpBXlXlvbh0t5ExRqE90Cbn5
e6rre29NrpwQjW69wMlAn2Y1ndbSakV5JKUrq5o1+vsEK4r+iRSUrhZR6xqpNH4v
BTHHgAVEPPkNl1tJNEvpnCm370NotfaIT6wH4mc1Me3GVukChHKsMrRpUny36wgt
L3UiiydL1dJFJnnXZGNHiKLAUhDaVUe1fwdLoELK8BI5EAYn791KMs6VFQ/KostF
tymyU+sJBCglSzcDpAt3VhDpt7JDEPzQW9CU48HHdXowxoaaZqiV68PwOG59uZIY
KkHm6nDe4/00mFfxRmZe7A0fJAt1f2646LAiVmoBEID5nFAsa1vCU3FEWAsV2Khv
/4agMA+2eqc4HPt7WJY24I88/k23F1lCpYzqtPN34rwdVGBP2W3jxdEn3KFeaqHN
NQxzcpU7UaQsD/4aLQxhN5QduI1XtlBh4wjPJPg2jW1kvo5wJsJhbThRjLe0vCwn
GU89oZPtulYNI7QU3eu4/kmed6oJG0ZCBbztkU3yAwAjZwgSX0Zp7IatcnPQ/8Zq
36xy111UGs9ovfdAjyDhHo6BItaSiit6J78b3YNjHzJ1AxGn3Qn+NLXM8KKIo6Qo
Ni1RIBVbncdw1HqKD5xs053eJfEMPr8f5uOoKb7nvIm1fPNVLUng5/G4EmpUJNRB
J8hH77bPYcPkzOOswpknTH6VY8mmTQNMRIIdURYffNzRAVLXYBrOPOP1nNUjvcoY
JJMRrNQKspVr+oQ0ONxaHAIYRgwRmScgNTLcU27FfOze3FUTUGnEu/DDXE+LCFSw
q3h44cue2hherQQ0l6jfyRHD7QjFXsR3eEZcl8vowB3OOCJhmeTSTDdGfGK7d+FX
lWIehqw9CP8QIiFp37lR0s/MdQcOzb938CGERgKCY0bN+xzkXed2S21uw/X3kCrj
SigR+Xgtv0r8EUv7oX2cE+J2rFRONMb9caiq0/Oz1vdFp4q6WfiDnmNSATJJUgPe
JAmdVkZLsFvmhGDHQCgcu6gSNZqnuZyxQwSf/N0ueP+J17aGWrh4RjW2wkXN6shK
QDvNdjIsfb0MzyyBLy1brV9mAlP5qEXVUPoF31rbRDK/HVNYY1mDDeBnkCDVKRaw
FsKjg7rWnq/qFwtxlSzOxD1rMctEp/wd4EGFSUOKp8wf5pzNmMJmphVfpINbAjFJ
+W0uF9cQIxvKv6g8gd+GVOLrBEwJnLKEo2/izxvYrCO47aLCOee+xY1ec5ifAcfL
lQic7kMSG8YqeYX0ilGF4AsVHKXZH2WUcRyJh5HYCfdnNtNmBnd878GM0SH9x77L
/3r/nYqkRdMDATenInzkIL6O74kwYxTEPJEuNSy1eABk6gtyPeXJWPjpChIBNQxE
PPQpt+SpbTi+fdPBBtZuVg==
`protect END_PROTECTED
