`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q7UPAl/XMroI+pS97rdnNnyv2vs9rUerYcFavfejwkrFJqlCoAw96KMjkb2yI9ii
GeAStDfhCwI/KP0W0i4dtqqsHzuNxza0i9IoVwVmGlCVqcO5+cjbrcbPVw9svlCH
nF69iz1Nr3CowBPVd7GEIl3UKzqayDzbgxi+TtBXBSCs2uTDhDDOnrw7tVY4DyT1
lR5oRGY2AJmQVoAFWOZNkn4/IKMT8tDQCkR9muGaMgD1u/YMFX3Z5M41lZfuaCNt
xnQCz2h++H6xSE/5ogjvyt8w/DL8G515duLeshLiXuAi0y0o776h6tIq9KLs/cii
Pn98OBApjbe8EXPcqrSNMHbQlko8WSBJWmxT3+5FvzhicmjaBZocnvSLM7NQ8w2e
Lh+8nKAznL2fxTGigYhQhuVMxvv+P+kAdvBT97fFlZx+pu1+ZaavHurRX74C1HCp
roybxTfMZJGyD1dbjntw3TAmBYKoYQtKTLTWWPfsMZf0W+puGT8QsXTn9LfObEw6
85+iAaZ7JN63Y3L34h7W0GWoIor8ceYn2K6mX/E42bQ87Pn8tXMgl4OeCpuo52vD
4+95FwnZuzb1Y+R3gL/tIyHhb7OUDKpWqtksaIXh/lJAn7LSaUxZsXLmFUL3sB6m
axq+g9mx7dpIXoN5t0h9A/Au0Bsm+0M9T85sHzCGDlC5nK7CSjXo6fxQj73FMK6N
UNY54Ws5pabB2YuJbqrPYOUst7SX0xG+iMY4Qg9kkKEXmZWPuSzahfE1YkUOk8bZ
nN3tsOyyhnZSZzuFcR6gy5nZvKoAzV8rBxi1xItpWzc9mLoian66Thj7uKqWo/n1
eQo/7dhL6TToiLBgRke3LLp8k507H/SRVWkm7Lwtz6KRicuiMaGRUlsLQQ0AREp1
SiKc82tTqDtywEZ18uI/Fje8NIa7SuwDbce8P7WgyPYJC1z3FGDK1sn7Caa3cWkE
XH96yU6uMQyD0j5/OzicGTSiVCnjwJzc2sjCd9WP1LRgTLKKh/QgamvDajPtratY
k/aKHWTigDcaOPPbxOSVS0qlBOcOUTamINTProrhiVCu7w5TvIx5881ekGvaZDk7
SO2MlMUS3QO2OwjmoAVCRYQs/NxHrcgBXGAuvwB1tN9769OThkwpkiDVCqQhbsBq
WXyRHau4ME9G5sBAHNHircS2k4qqnw8LBvKjX5j6URhtJtQwGBEgUTRn1dxyW3Y3
pLkdpd9YM0RqI2PmBLAYFJfcUQxcCHQRxMSqCHzrV4ZgLG5c+BnibxI5BX2SNeeJ
AJCZmyJBNtQ6B11WN7H+hNiYteDh55L0ykT7IFosmMtUs4HSvxjAKbQsMN/uCyWf
K9mAB2iyn3QeWqzIkCNXHQaAq5j/ysU8dSLUy8PV3h1wXEoPBoI5wrRZzXMUZfAp
zFaK0hrlQttuF3nOpiyBD/w6OSg5OPSSKN0htLyNJ+d1Dc1XGiQztfA+L+0pJawM
RDKcDprxYYnqAsF0HJTBNnJir2IY0dRuctrG3gteNOCpsb0eUvASShoBxpCzjJYI
CW83erPcVS+IlJdHvz5SHE0Em9pVr1Z4eFfWTkFFShX6bOVYbAxrVCP7jf6Kf7Ki
58YlQ4vJ7u2jD6976cpjnLxcKRslPLoV7T/jNotLvrxaKtPVLcHvsz+A2JyMFRvr
hK1OIujvvYE0SDwN+36/b8tCbVSY74LZDmqnj7cFU0GWfH3KB1IxRZ/YVVrlVpTO
hSxbIwVSXjgSosQnZLKMoy86xtVZ9XhSrfhSg/G3bN/twWy/M++auwHzluBop6PK
R7nULmg4RTTpkZJQg90fvLQKxzHebjlQxFKBhv1MlfmcK637E0qPsVRmJkZi44BN
BS8GTpMd2l32QkD7Fj84QaS5Feng10tZKJCelcshy6+LO2S8u+yiZL+nGzT55vod
tQj4ML+ZTsDNydLpTPMwxtYniC0YGsolLzU222WzHsD8LUvPvc67f1++ala6mJWB
M63HzKEwu5BwDyCWEW4N3CUzmJugH6ve5fQriBZCsaKPwBEVQeRxEyKbinw2E5/F
+kwjKropWx/mgxMMF+iQ1yfPi8dPCLrNWseyPYNW3fNwBmV4wbbGgYvY62+YKnQk
PMjZCshI+uKqb8D/g6EwVQm5IjwrQPAxzvaimHuYAQowHSktHfX3lnzNm2x8MrDR
fDp4jQxU3CCKy2Rra+qX4rw8myMqcoVXs5g+u7V+W8X9DOdWqmoAas/bxgfHZU/o
AfLScWOS4bhyNeD0X2al2bqloITunvSPUjU8J+xQShVYefOF8zGwVIy4nnYiVlK8
iYXkEfJaPon4XTqnVJp28fGVm1D8llD5NJDGph9PEYBB3BKjXKDZWk2XmQ+aDlgR
/J62v8Y0NsDrHkEM7vtuBcTxvEzCoCtJkehlyltw0U77xo7GrZ2/G9odZ03Atk8K
QvADpV8h6wKK9rMmFhDzeFGCunt6d1O09d9Pe4Vm0yzBkKriiQ9ocUEo4QJN29JB
32K6wf4GMODplHEt4C7J/o99bNuK1vJSwj2gZshjJVBBoC9xtMJ49lnNM/9cDpTy
cWPHiltLSbIeFcv/Dv8W6KQHjnYH6IuWsLkF6Ydc58FSbhr0/C488ZefZRMqgYWt
Y+QXlDr4b+dxr1q3C7ZUuoNIw5TWsvvOrXAaP8NaJS1KeELYYhIU7AeLdqTbaBmf
Qxx3NzL6NfTatOgpuE1xg+tbjnl412zXyHDQuGYKh6UkvxcQmzUaIgDPRxIHCsUg
JhQtMXf8RMZlQyLaQ+iUOPYum2t6dbil851n3PHEuzL/8x94HQ6U32KaX7WidCPx
x9OAo4ll5vw7Co7ZcZANQqxUS4us4B40Zd1cCBw0RU/fbQs3F5/aSGAUTP3lWxdW
DCraKjkvxHUO6negVUOiuw1VTWvo8NCdF7rXb8bPwBPwQjGT1RUQoRpRnVN9Gn7k
Zob6cL8KbC6a75sr2JxAPpyMWorQMRHqwW6kY7QR2RKb/lI1O0Jy0UjsP9OioExI
UkGs43/ZptftLpgjdQNu3Rrmh229LC4OLXI3vYZaBu5DernLZBOTFiSwCBB69aqo
dY9SJxTYB/qLm5+mVxJq0vE1MFD81zYLMy5rEl69wKXhPJKeny+64eaaNOq5KjWm
wcNXxeSx5t/XioXkiQpglrQcMOu6mgqnk0RGsHqYeQv9wKsCHEnLoajAZEEA8EBi
24vibfnU36HLxPr9psHPW5bFX9s0PuBz0bLafApSM5EVjOp24oZbQhAASPQPH5Ul
G3/DcfcnVdGN5l+hyMglP02dsX0w7hDMlCqUoWSye3a4m37EcDzrwwiSQjhBbKqF
5gKfTT6C5TqP7aIMztICMm8u7QaIuFfd8LDjiwPMooVJEsLUEVq3IfgZe6xR3Eiz
GdPWQG7vywXPRw9/ecVbzftBIUUZMWjpVngq9U4WZ8M11oOZPBi108ANwClvIK7Z
TcBnAib2twdyNEy2YlI6PBmHpNrAlIID1Qu6aMONLm6GJNAud0CRPdGUr0bt/mA7
WOtWPt7ksL9TuvwIfRut5qmKkvRrM/hYhyChoQInnqWbqdQhdga/3MSc6uOJYh+s
hzPYlBrfWvC6T70BuJ5O7IvKgUzgV9goTWpRU5IFL381OA7MMfUlKqxXWZDrMSNW
0Gt2CcnYTYTCpk0jESjqWolSnCQpM0Kwb6CG/6z6poDXPbMI7LpeHTjP9up9nZrl
mPJKUGO/s1kIfeJy+jcj+coOWVcJP/XDilZ7b3U1SFRHNJKEiekWfxjQgVwhDtia
IM1849wkgl1M3d9j8088mO1OAbBV0UjOEXp4KU1dhjD9sebXBGXcCmMS9TgVGJN9
N5A6LGv5ANjL4nNpfI+FO4PBv7/sYXGPUecQCwPpaq1eTj2VPztnggpvPSrReZ9R
gpDnQe3pd82fJA+WUsOHZoo7K+Witdt59oMO7GTj4EA4XBjB/sgSs1ihx99lbmqo
1RX/2QIDvSGubdx+oHgXqDbh4JZP8R9YsI8gRBIZRxTiWxVXdy0OlvR6VftE2Kza
fQ/ly/4Y+sA0xHLGW2I2SULTljMmhWYYjB3a0xTrDV/aWELzT3DZYslQWCP9xDYp
3vTnEKmwRg8ePeVzi/qTC6Zk9IHeShPROj/ia/YQzzTFHrcjsy4a6vzWnTybamSy
jDDNJQw8gg0V3hhNtT6IokTP28JxJiVKo59OO+PcYO0z/fNllymC4mnzrCi/jxx4
BUFslXBzWq7eAWP5radYeOQB2Kqb3hFAGIOu2h8jHSZOSAaVxpaQ3154875rHjK6
GdOHtt7vyZIhygXuRZiio5XsEr/r5w1MqSBrRWqq06/+qLijqMGd47NR2SJ74L+X
j+vJbJPNCGwjNLBvMrVYsnvmtGZxftkqM0h9QBiWtHEQWSzoh450iomcGDPVCDFI
6ojG1N+CQi05VIxKDyOVb7ZLfavK1SpHR3hD1DsTVzbNCp0Dvu6hLFA4vzXgT4RW
2XB02JIab6qJEIM4TKccUuHKrRRvozwrMmV7GkLsfR5joYqmo16ysPxNOJMC+ljQ
JiNfC1FGyDYGKQdCkaDbbJDisozJ9Hcqvz/UlEI4K5n5cQCJExnohbcsvdye2UIR
UibU0WwqYxkQMIm0b6FLvAlDHk8vP31G7EMZSXEOYLsdADpMJpoAySY3G8ISnL3Q
TLJoeTiLYDk7xHX+ymDygBQgstQ56RpIxizCxv+dfF4rA05djT5T5tXCGCx7QRa3
UyRefX2PTBwKV6OYzdn4FoGy7AOKMW6uU0RcMidiWZIoHS23J/XUGI9FUhu8VM6T
f6cwbZkQg9/nOV+T42t/W8GnUgX0f/iNCNVPMSpAmK2b0AgxmthV/Sv6xtwCxIjc
bGzkne3O0qLi5ioSrs55vVgHsfXNE9M/a0YsUzYe63jp4B6GJx5GhqdBZv4xlpZZ
aGoDlvLAXDaLNh+PIWHrGyIZuFcl0vuKs+amSp3olDKfjUhgigWdW9fC59atQF56
LFVe477CYqUecdy8TYszgUcGOheWScp+QIQj0Hljr/wn7sYrm5sSq16z1MVjeXA5
CaoZXbmsRkqmF/Tn1dhCSPmP3hZufGAVZST0HstXqxMQdiYJvasV67orEuB6Qhgq
ubYx+MeKDu6Bxs0HgCXCrT7Rj9gUHAW7vA9ebXwTPJWyVMbG7e8/GBnyRUhW6sQu
s1ZTi3XolPYyntt4Sb8v5X5PgmcuUcg08nPGpSwRLqXifa+/1PROb2Tpe8aWn5pG
FQUcPcX+8HZU8WFX7B6huYMuFEdSA3Uf3+lHsWWJUW1gapwvcb/4pg/BVi9VkLr7
DUWgMFqXp0G3WGcvSiSUKLEXNg0ikcA0tBIonmaWnSRW9a31UMT0o+1w2j9GQe6a
n0NxtHwNQ8MLlIgEf9vR4IXPxxbx27S9Q8KvQ5jPZmFGK/OemIo+bF8+KH2RRvYP
fzbe/t9bHggLTt3PBQJnJ2XjKWt1rUk35bSorqPa1gZqhn03DDgqAYSz6fAfRw4E
fpUDxAaU5EUm7jn4l7/om40QkN8NjS9TtKAdt5PvE52yWEUZw85+Ybgv5k7Q/Guz
33WTGvkW7FTcDvWW/VCbCkg9yQT+QlZe76QJr9obp6BLY62SxfRdErBWvuJMZ2yz
oxP5VyB6Xie6gFiejEHsuPLPGj8QdQiJBbmPBuyvf1/FICtQfvtRdp2XShVV5Zn0
ACChKn5kxGtBHKWj7mgigeCpmhj4/dnDlik8iqyuQq6Rpq9HmweDfQ8vptCL2Teq
jQcH+mrZpihmn+nkIPEjqmVPd+y3QPmtd8IzI7vZ+h3YLwlfU8aguXpOpNQgzpOV
3sLA7Kpqf+n3D3Jb3d+EZaiqYkZ3PcXclKIdL6un8+hN2c42ju04ZNcXWx78xod2
tfyNYsSScM3xLQpFQh3kpOp0ojN1DvwrLVekP4KfBTlO2RMKAiXYeccYIWTmvpUa
X19ZVmbCgwjT+3s2I7ZhGPqcApgpRcjx4J0HL25GGmiaGw5uhu1gh30sWqCMd8vg
LQUMLGfStxw1MJkYUpJybhTJLHRZwCUHAFpqdtifpZGhJkj0e/LTM+o1Za51QEPX
3wP4OHVc/g0wWohAp5ccje3MBpY4/btcVehrX7CwpA2cA7QjjMRqLRRnhznE4xNO
RrdPsd58B8fy6KkimJk3225jiYwkirSXWAVC0LOhWw5XY7o5oDOlmpZ8I8ahka8l
4DdBoAbagLB4ENgpJPgLfZ5sFxw84s3SdKIfkkVXFGyFC1k23eC9UDkrwx686Fdm
gN49ih9EfljpGwnweFUsFjQnysGac9Lxwg0j18eVggiCVHdb2LP9VE6QfRcTu6F3
14zifCSS9s1itT126ktmENObOnKMSCuQ4R6omRh5SR6DzKMxxS8Msv3VO+jpqKPf
oF6JLfLxPj/J+s30rHUSGgvsA5kSKxZS3zoccV7xNkELv8EM1mdXdUhIwuiElB52
glevtFSgRX+qUDQmbxBel/qnLy0cLWAqmJ88J6ZrJp8Nm9CeBAiIGjD9y48vcYoc
cL4pTuS2c3AlrGSLxUfOaGxFXfgXEgz/iNACfAjc2945qvf9zuzPdPWHAQNlMmUd
f6Ec33cTYG2cj/9qR9TR8o1qou+nQu7kG/IxOECvdcImsVMJaMSZuTDY6r2Ct71+
5BPURKXGaAKizwiht8OjwDTS/E7xmu3xqq9et/IfP/6Xf2WxuOPDoSIXhf6QPJh2
WzDlbBXgjgCqfhw67DBBx2IjLOx5frD4lZqQz7kLubx3MmOQkNhthVGeiutS4t6M
bJzKSovwSazKUkRo/vQW3EoDFo0c2qkFPoaWnfpIlM/7uszP06TWFJhOGrYEk+cT
uCuVxZg9MPDyL6pDhtfCREPV8OYD2aq1mOdEW26yx6Z24Dcea3KsAYb87zxpOVqr
TKK/MTvvBQNmaTyNK7uWg2xhigFGAUGaDbo/dCcXYxWmzA29Rk0bgKfYgFQgGYi6
o7XEBGs5Wu25HjXoYMEM1aEMMAt2YrsQJJGmV0PxY7ZzR8pCYpZiWh+BS62yIPd6
zAerSdP0dGHYgZUNsglEuTJTnE69viGzWow18fS8lXMePH48/JaFnYLPsWNcrO1m
jfMYnBYVl1ISctdbZdMLxhziFiuI1bGrNa1fI2Mm4hAx5SfG+Um+G+MBYpDjw+WA
/pqENaJ89YiCCH1j/71RV4OQ7xxmW3lE3JXZy7+dJyrAfdnlO9G8phMiXDWabU2t
/sD79zVz3T+gv5R0kJjMnd0u6kMVRJPIcljIng3LyOcgzuSMKem3fRYmlv5YM+ZX
vaDJ7whHO3XfD5wWapUvLuicoznEhsD0h1dxXEU8UqhL+m4FXY1Z0Ot76tDt8+lZ
YADxMuCPy4KF/xbt5kS/BQswiqeg38Bv5LtYYnlg+NmWCOAq4EWaOXE/ODg6v3xi
Ak3jTFtNjgQZciAJp3HzxVlL10ojs3NqLCl/Buz1RrwozSHp+7kYzJrhpfU93cgs
r45uHFsXcT/KEzSfDAuoFXPGVNRtthNP0k0pPsWwd/TarnHGXwn3TVFKH545odpK
5fOaoCvteO7jEbhnmXLQHt88UdzGri9bJ1jRRugN8K1dD7cOCal2jE/zvbY1lQyB
dCxbUeeAFuTyJsx1oGRp0eN9+gcQIl02KyFEY3YQ2gc8A2mwCnf2TiXfmDm24NGy
wDHNCD9s9EaoG/oFgjpmhDF8hAS3+OtZK9iEjfdY6l3qEcgPlWgETtJdKcjDbf/o
S0R1npK1XvHWw+VuSiGoF754ecNQmUJYoT0c8xQwhP/ms48BZqDmtdL6I4LCrOuk
PbJ4vZcGbi6OoaUimOETstR3SqUMvq7Jro9bNsR9jyo=
`protect END_PROTECTED
