`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0dChTww1OQQZlgm4tT1iX+BfFQMSTXzS5wArBkJnBcB7imDwcNuT7l3V/Tx6yIsv
xcSEFTuU2NKh6DSDpRT7tAOoL/Vgg/8pb/w2kVAQAiSAcwr7+wAgNJ1HSQ+oGOJc
+TI4iUPalIHaxzXRCqDZPQOhdPUpLnDhl9RoD8/DophIE2PSHDntXF012N+sAUU4
6GRS9e7L+/Dl6BXkzjvPcmhvqDli+z6hsrHnuc6iJzI3V/BwqaBQ5tcE79sbnRUv
WIe5V3FBsuekom+hnt/VhRei9VQK9pn7ioU6nlb6s2HJ/pHmRO940S9BocXg5lz0
FiEF8C9s5IMK3T0gjtONAbbic4+8LOO8MOPqFmiA4hz88753t1qYU4Q8DlwOfMRM
FByJ2GtYBG9CmurBfVamCrqjnY6Ve/cdqyS9mHTgHK36mHNw5IjQBjfTC/PgYmGO
0lsPxRNXlb5VwJOfGKzIze6LzcSYOY+0rbmQLtYjxNYR/S/RkxbbN6sEmLv2fN6g
gSMq9lctmtoseW8HOnSrENkWizEY/cS8qulK73j8hWeWDj2EOTGu+Nusji8LEUMZ
XM77dtX94IF27jwOIGRq+8+vX7CUCCCm69a+gnetdQmYy7NIEVlrkpj5ed1vTy3w
EhCvvXMZ0t0cXLIeIDxkoUJxCp17DmBjZT5cnoojiP15FcuMiPWb3b8XcOxQ19yr
QHxZXGjI6m6D+6F3QojoQNoTJu0etVHVEsd/EblJw1KHZyXRCrZwHZkTIy6ixCqe
q5GDavq7huZuZ6KO6AoHjqj3P+YkogYn2XJHua/GxVv8lIyrlg36HvBD5JfhMa+2
aVW87tscNxG7PvNwpuwm9CIwqUNDlfy9yboQ+/aGlZmkQoQQN5/x4U5HlgppzZVv
zwOQJoyQA/mJfk2sprNAtHVsI87w+aPH+8slYTQaFcSpbSRAA7Kaf/vIpQBlggEy
Y7bTmbvLS/85xUYO2Eb5tg==
`protect END_PROTECTED
