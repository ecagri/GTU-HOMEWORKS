`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pB4ti0hoC8GG/+p9CYcgc6pOe7cg/dw1rbSEBg4nN+ZP//awTFga8Kaa2CrIrhFi
mqNgkx/V/sizotUNvvCxU3RflUXCOIw2XK6KhSkOyOjCSmYp8mlwAvXknZNKnlEn
56fCcGUag5Kx/iN+QXZ1jU173S++kdTZGDvrleeLNT5YcbY7tAyG3NZYwrrQuxGv
iuB3YXx7DqoVaMctkDrpqm59pFGRYO3hOYhJLSDKrVB8sD74Eodg2cZ3/x72/0E2
Eqcl0OSos0GBXv9Dsfw2vcwX3UEnSf0wOTdkvGdKS9OTaPCmofj8+F2WFSlBGdAK
LBYozt931dg9U8eN6GQ+Jl4CAvUXrWsBjYvKqNf6b/1RSgaIkIqgJGsHhRBnqw+5
PXM/vxVTxAXIWS053j2QCr/Dpq6kjB2X14IXMSCJqTdGWmk0E9OiVKcvxKKu5ow5
MZMhkqwcImyVaqFkA62gPgVlE/jHYzHHJFbwbfLq/E1SkMhcw6CQVamCK5kSZZTl
wGRpAfaA76HiFk+oGZdorvGXvlAsxr6qnwfmhbtc8RDiHEujdIFct9Qs9aeV5csa
ziV+eHZK+YVpDIDOWZ54x9KusPUgjkfmn8AZSUk7JDAc3mmNieYTRLVPYc4mP1v2
G6Nv+LPVwbqzp8MqhdTweC2E/uEiewqqbVnTcCEjhQKT7E86a7KR3BZbU7b94B10
kbsfJzLrvvRtmXjCkitnr2vEW9PcBRRun7uAhL/4ZeTOD3AFgDxqiIoojJkUmhDN
1JbUUy2NwFvBuXYEMtk8pwaVD+2DGMOwePeo42xkXUTZRqJVlDQhUg8ouWlOesU9
wcce9Mfrgu6ZcLL4LUUeLjcDoSdueHQyuIQ/mXQfWJ3xw15uG8udL9mVOyKNAqDg
SCEweIkdFWSu5PWv9cEA3oV38ETDa1cB+UZR8ei6R83TbmkylCcOzrE+CT9h2cgC
LQPY01yDAjLBy8J9msbmyBOy0CSKboqUpafK2odPolZ1vLu8wlIoq8akMKIxJygv
GjI1v3ZtPo9iF+C/UfXeZmP6eYT7rjKUFzfs4hr3SzQ=
`protect END_PROTECTED
