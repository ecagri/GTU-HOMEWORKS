`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+LYnsZyC6Sfktz9AZyl4jCvjJuH2SUNQYNOHTLaAjbUj+zbFJSc4/GRfmLevV3Y5
AP2MFRgC5lmFTuZ05ZO5dLwaNssU+P2OhgL/3Ksst7x/4jo+Ls5XpQymTbuR23P3
86psSqa+Hu8GfeoBGkkn8rJkFK4KexjXWVvWE8A6KEsj+7y8DPtbdPNHL1CquDAa
lNIqCZnOabRuKiC1DzaLC1BnQv5Ylsyp7h3J9n+0KiTXTolSV6r/51r3OsJ7Hhvi
qAS/ZX5tFhtmQYLedSIY44aPGelXJMkdtisow2yGnJLvQkrkHC73lsKV2rlMy+N4
7aA0DCXBESeHEn3HImBa0H1zM6G5UfS05LZrqlo+lPfPVJiurV5SRdczVkD/BCKC
wt8+g5/KRMVdBmDs6GzRkO+wZXq/nREksD8abev9kWCw/dAd5DLbO/XevWhAM9jr
PcBIRQDYTE8JzJOV1rd5CiQpgF1D/VWqUzTNFL2nNFq2+hA9N1Bt/I8I+94Vq2J9
OVXVS2uAv8CahbJJJe62/A==
`protect END_PROTECTED
