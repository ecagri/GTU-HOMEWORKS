`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EGblruw3P7BsHsp8u/BADNTGoBMSNONBnVUz7JlCENjXuAfKbzKy1zGlucIhM2te
gaEMPeN537Y8qO2NSyBu8QhMRKVSdboaWYNBxrgNMjvk94vo9Fp70VEbW4V1wHtF
wkge1PtQh6mxd7kfy/lQdyBbWD0XYR/BBRmvzeB1AWoaKJj6yYUzPvnBmGkPrTSk
Zpz0cbpR4b1E4w2QCSqabK5kZgyqu664zTDNvkQZcKRawMk2p9QerWUtDyQXfLwT
UzoiVFQcUs2y7RVzNH5isk3JFH5yrigCjRp92aYWUr25yBp40FP27zz0ht+wpnSh
Y09QvB+z3j+Gb2qg8/6yu6X1Tv6J1FASspOH3HvumVzWEmtF8QkZSFXmqKbsOJzw
Qem+FD7+KR3bqAWzNcIxZjUzyBX/8LwA+CxspWyrdn613OVO7NHDahFuLgzPDWbu
oS1sWrHN/LWXUQaP9+atguY4kzK8glH1FLwRoK7HknQPzDV/G5w+iMveFxA/13gc
rLx0nPLv9KHqIooHI+MruWMBYSO0pOsMFUt8C+XDQEXBnVEuEvBUhbyzp5v/ehI7
fXpGKshd6E81hdjAX3hUTYR7Or76J+3PN6Oyk+B+7OEmMJCqGpvPnH5O6VcYnTVT
/VULPo/sfwChdYd2woOhlMG5kERodIEr1QWWcpD4Bg5DF787bpJBCoePRauiPzq7
CyNNqakSwQCIPgsku0F2jKfh/e7FgqN1VEEA3yGQr1mt0YDtcu2bQfQK2hPQMZkU
pHMruOGmMC//Dz82xUhUEGDu4wAXNcY4BTk47G1m2yJgTiBCqdFAU0Mns7H52Wfu
kcUm+3tUFtKaRo81DhMXNFfFKwnnaY5OOgS9rkvEG0Jj0yq1CKrB1Qw7pRsJAeMt
CedY8c4Q+E/KJCV3JIALtcVBx9qpCFvsdt8N+dJAcrmqJp9GDZ7TvrGAgXUTz5m9
pSMcvGqD3C9+RSvHlGQue/iZqzmBuBdgaP5u1hh5SHr30kvX6RGNGRX6iE8sntjr
Fbg+VCRxD/I9vWShqnLDlun+kv0NAR1GdXyv+52sS17JobhQrn1aQOVU5JsQEusx
4skw2fvJpjJK8EhsRiVlxakQ4XWocsRxDgRF+I6CEEokLvkWum6Snd8X8o8RTjZm
I2oXQPDrxIscQJN3YoD+DA667yiAeOMqgeaGcfUCzGlu5lh3W2TEOjJBnQWqI54G
q+0wRNJirZJWsKswn2Py2jqF9QhXuWBU5arNQ3Qu03uyrp6ltsdBYs3rJresivTB
kMB8yYQvhSk/f4biSEYFeI1F7aN82udC99knLFrMLwSNUZat6/XHR67QWD+5Mtuq
TsIuOmgviWQ7BeGWCik0j1TukRns7nYok+dGfJwsdhQjkaSYi36k+Fb/0H+rZ1rs
+01y913Hxb8LJBjvk3Ida4Z1l3ViunPfffrZf7RWN1ppU2c2yHbOy4wyW+3ZAr4w
KTZTxUDLHOqaX0xXz4KP1aKXXY8VIjSGRFRJxZxJiJsoA9RNDEEDED8eUWHAvoKB
UOAjSWsUHL+V1MnZOPJOGvXMFOvEf1YZ/cpe9XB/obKyJFfSXa8BW7bkBXHLLOzS
UMyA+M6xzLd7/k8+DjnvjP8BhmsEKBTLF8HWCZsWg6UiDVaaJ8O9S+5YzT/PvsM4
BPKKuFXtHWQoeRH8feXfTXKxyyIh/sPH1BT12qCAFqMra0mi/udswhkvCt4J7jHS
CJzbJTWObC4ZVBwH9viJ6+fiWzevSWJQXRql3uHGZrKsgBddBVi988DzO334oZoB
kGU+VGXDWrhtSzyjVjExiMjJavi07ccQTR27yqlSi6BBkLfHzWiSCKkgJQN5N7Ql
QhzoAXDeMp6G9Pi5DQlXH51sYAniUuUjLiK5LURjnRi9vAsZJBWSTFzrllSA++ql
+UL0Ur30x4i679durHxOv/bBJc1ZnhtUMqBWSzHKM6VkSdrUKHC9KXnD85gEppAI
l0cgtO7Wo5d+0gKPUBE7Z2SvmW1GcXXbc2hcun/7DiLxQo5LKfREKSD37qrBXth0
iWNu8WfCY5c+Pu4IWMFztshHI+ZtFCXItP1BqxrkGYdaI1N8AwrCtpMQqc7T66wT
lBVpWMkiM4xGiZzZMT4/cCwgIX0nEf6XvT8FR/2TKwPFkaJuSdPlapQpIuUtUpIi
wJu0o+QziUnCSsmAJDDW6I8YI5lS2T1v1yttDQ9ajb6a8AQ5XXydiuTBKslxhJec
2YC4ShtyVLa3wwDYe9+KvA0OxoCW0b7gxpvB/Lu1BOTLjaHSuzgPxMqALHqXuCPY
AxCBMziL2NV1/SVkiFO22kcddtK6oHTXRYbXkbnwpyXTQvdzLPSFggDDL5P0L7aF
ZTMmUimvr0ZMz0OUEqu4C8irWVr638ZFpxP5H+cVMAGPktsOW3lwP7if0X9wi9lk
fUSmxRJ5bhxXvAAOFh2gtzZDsICZJt5b9oec47H4VmycGOMzgUiFo/GBMsfGo1A4
4pO/4t+Gyi/4dzqYcZ5yBwIfV3aL6xokKuJo3uFOb8+vll8qom+9UbUN7a2H2dpf
zh4AzmnImwrFA9w9hYHsUC6WLZEnNhSVVUZx2yii/Rfo2o7QOzmOEs0Fo7KlVmsi
f7dLEBadlBIm0TCUTQYkwNMwctOvalhDBFBxd+dYmJBzGlvOutBOGnEKbcpxuKug
`protect END_PROTECTED
