`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hg7icWKMcNRwiVtRWSa9NuPsvC427LrLfDraK2jK9ZrdB22w6xgkx2eY1wiciY+Q
hms9mzDRCDXqZNoAQErSchF8jLxeTaF+TfsB7L+JE9kzJYPYNwRS6y4ds3VzVCYb
k2Yp4SPtmbl2Yydm73rzFw4DAwV5V8e9zrel4OKx+vLT0seYrflo8Y8yF5t0/xbK
XO/3o6FGDMaCk0sglElRmkgHIZf7/Itctvvb/l7VvsTqHMHlyTRH0BMc4V8YnpY3
0dM5h+or82loKlg6UwqhPsNIc3i5KLarhQsCVikzny2wCvFPfPPNV7MIaMAJWVRC
C3uxb38yvWrHbfKWCEhlisWj1e6HTY1RxDJzL3IXMQbwVt5n+UnzkdEP/L6/jXMv
cXg4UYI1O0FQ0zo7YroOGb1UgvhbD2DX1Binty/G61GqE3ai+hKKAZF6xxwufnZD
xBDDpXSMDFAOAtk6zMZpI3T06Oi+Yl3h6ltRdUYCDTgyuYZ0NDTJCUgTzAp+BMC1
BZ6/4X+Ae+VtZJ3qZlZZuCdI9ry1v4AMe0ECOqRkA/wHEv2hbPn5BDe2TbWuCKhL
Iw1Lx+OthR4xk97r9BStkfNRL3QbWZOQUYq/rKN4/84V0+4tvDnsg9WIqll1Xxp0
pgiu1IEfq+b47Ri4awlCrzllQfXSkfnVqGBmak3zlujN4WKJhvIV77NYkFxaMtwS
ppU1jHwa0itsjfI4MiG9dVdtlTXGRUQDv43knJLRM6nWLS9eHuMrjYF2GcbkTuIE
FHRfG2UEKcuLoAs8l285eNQ9sLmlH0lBQ0XQi4D1TyZxFLH6F1EJgCvflwFKfuum
OSww10DKkIKeBUZX6Y3dVKU0xohrr4Na8d31xJyqYNWseWNkm+5y3eQJ23T1aoxn
GEy9rBSmrsBfdEdBE4hy3KO4tqUFYPuQXrUvtW2bBCXsSXr0QZZf6JdSHFrFWA26
kOo1ZyNRRi0RzVMmhpjdSBfi0G5IpQgMRTQwu4xQEHAiTNecxGkfPZAulKIVTpLC
Pv3lHlP2ujCxXISOUxLFglhxae+pMqSLNo892WzaahDnX+MlHuKkXQKi50VI7PSB
X6kpCdRturkvTRfU+CoZgHajVdWFnuSrtnsfDsonk9D6nm6MksnULLMTMfel7NKL
mt5JxNqVEA8w1gBeosoiSzqfn1S0KZzHmDJj/QVY3HfPeZvHRVaSotgCFOAjt7kK
t5/3+Z2pJH8MLwbrB1ilRKQSOcoT+u9qfNL6z0Q+JuUjj2eVVghyDHEni3r/tYq4
9xFYeYJLVaeAtHfhFAfcfEIY1T+fcLhLjoXxomB8iI5N8QX1lrQkpKuek4VpLPZR
8bY33I99mz1jWLM/3k5COlQ93hIG/DCOAINdu4k1qYAc0sfz3wte2CZymG9wG0YQ
32/KpQdkZAV6/WSu/i8UnznEHs0t2wv59iDiTE4YzYA+QFinIGgRaR4K8PtQxE0h
K0YV15g9V3IyAKyHgq0uyRunw+sg9QgoCmjdk1gnWhFs4KhaqGWRzylwbJ9NhQOD
U1gVhjVgQkDDQuRgvtYzvd57kej9jQj82adVTHsWWCMuBPrnUkZRo3mQnj3RUZx+
uHV8eOX0JX4XXiAgX4vWD2a5oa7Dk+8svRfi/ajakilWc8Yppdvz8f9TI+9GBUxF
xOeAJcQQoMilDbw0mDYjPozh52vSJbmOHzOl1U6THRSf2jEHuawb5P+kCsDGne/I
AjMbIec6h0BD9yjUjE0RntchwffJgbN76P+Y/LE6zwr09E1ZfpA64tLhZRUKTC9Q
0ZASgK/Q2Lsb5UDeKBLOfbVOfwDlRaokrXEQYbeubLIfD49daltcXV4IttNxDQ3t
6gMfUEwCCkbIGw/+vZt1gJwlDYbGq7NjQVkpqaZIa9wh+SMPPfupAKMDDQrz86cY
D/CamwDjzJFrw1j0OugFboy0YzpcM3grxH+J3nkohmw41fvidtQWmxoXoAm+Fhjk
Ng2vb3UdNzaPspMd9aL5bideo5hz/LJyxvn9eshdZNbaMIMBC2QxVpv12J4kxiTJ
78roRXPovK1YfKAey3F8f+9zwW39YWtLw4WX5QkmBDoA89uaPVuSKbEGLPUfXs1n
xtJZWsehiyuNyrlUXqMmVUntr5JANTlLJF2t945XxMrxXMQLgSpU+mvjuhUD/oEi
hOzZIK78bkGmqqIRwmy+Yl9ZSkAsBtgExPd9J/W3PkSjKVcCxYnC0K952+vjlne2
gKcBfkDAn0xxwVmydaD0NBkorN3d7c46opp27BcqYzuqdSQrYYNVM22JDrnNayQF
d/WThQrmKmCSBijYZd8ABQMSTk6EdnBOqp4Gl/SxWdMLL/p8tpsbW4jpzLjFCD7O
+RL/t/aEM15qlsBORBIst9o6ug+ah1j3MTcyDeNNzQCeC9mx4klzZVxEeKwA+wUm
CGn+33eM05Iy/WhXTrQOHhiuLbHjBLJQHSRBwjpxIGNmSndF1pxuLTLMMKGk7dBU
hIC55qcKYMUMBKjOmL+5Jy+osJEieaOoJvTNbQGz66xNdrmc9YIVznwo9l3k2mSG
KhZnZNeE6lvvnte9PrZbFHXMS6btyUdPsg+uRpKqbsWroKLX3jhQULInThs+F/0C
MmrcufssAcGxhLeBaYX1vpy/lNkHLjR/AUbOdQuAJg0ujaepO4O+oHP4f6W2Bvyi
IFmZgpjzCTJtNHbY3BsmyZT0zUKvMYhh27CdbDRqbafjp5crDvVC4uyjE/Ghs9Jq
8UX9aOhMdeC8FT7ItuupNK6YGSkpKdPVslQ2r0q5T3r5HjxZOgBHFDnYi8qygAru
eZK6ofCHPwONztXQ7RSkbWRuhXtnugiupjyLno5Ud2EoGyy+e+8Z0OSh/BRsJcwc
ZIpE5q7QvoCvl2qIBAL99GASJk5RHIB47W3o/jdNFKLfCZ45XggU+nHlcBQ9AMQT
DAYtO88zyqd6c4xHVm4ENbk70in+ryt8lYRknWFT1aX5+geyhrHr5squ9hkunKgQ
nvxbrEvj4xVzu17hjoyZV4i2nLb8Qe1GUmQq7mSlYo4SY/lxqO4BOkiOMGhxGW9j
vKKVnSp4LA+CLV6xBrszcbtDwTOcP9FKt3xjXcvGwbDiL3K4HndiK4ZYNZKZaaMy
1jyuz/qfKh2N0yPOkbpDhFhiWTpaBB7MbiVIa3rTgV+OzOdTWAok4mjmbs51ASP5
v+ScF2FPx6DTxWP/lj+9p4jYYaYCuC3TS0SfEAFVRd+pWYmeDDNBZQyYG3utG1/x
qaIxiUHTMXRQLd2Bpi3TxpxibaGi9uLbkqRZhglGooGN8X4FVSzCPPxoP1i9G62A
9lnuWZP+jO3+m7zR+hyF70VHxuDcL98BJeBdm+igSZBHcmQoDLZYVeh8NhMPPs/I
b71I/LQhm3CBj5Xda7rHRPc5gUOnFl2uyth/hCIlGwMaL0GfiTdWm0mTIAGq9B8A
zcffb4tLczNSwSwhqc7k7vX/RJoxOGd0tq/uzfrVAyg2kmeBsGkiS9onvt6oCIes
4qlO73eSiOT+IhKSf86mMdoiIqHZttSl+VLaWqa3z8DCtkBliADweJ4LfPcEaa5e
3yHMdOk4RiSSM4qwsJ6mPYCjXrtI+xxTPA4ZJiZkfLR5Qohkqcf8jveacHgvkT0t
H6oFYhV7ik/+VFlo7BurfSM6uO81iQCmuzRnn6dHzcXRVPEMftPA8dW0/cL55nCg
7lVNb3A3vMOLlJLYo5wa21WUO7jAZfOP0M++6smOPE6WvGPD7SOnFNHO6pChUj8G
FsjNMmVloWJbHs/DWgUEPas6uniuBFuutOUWscaxoHog7huCqaoi504csz7EpJ4Y
5WYDG8Byhv8kEsmPw0qyjqc5XZhoMEmCbXfKx60tDnM3BjJsgNGQCXR1gbfXHqOo
7HM/s/O+Wj2IG5hG+B4qvk/QCCX1lCPcEAHt2IKWm5SQor6vNxHK7H+ZSUpknreh
psTOGQK55pbrZfK+ON70cDhZ9MH64ypS9GJ8VlsAdJpL0oGDznjSs8G1eSybvBmn
Kr9G450/1y3kWIfNZCsbC/U6q63Uv7uaqxhPFecmwV74ZNoCaHR68BDJ6RG+apvU
JWFrhPYOmcwzu4MiduRu+X/6irdbtJgfk/+j4mC3NOzIK2itTz5kIGqW/F4joOvQ
AcVJ3rYESr27yhbvCFV5NPo30XOnKPHskJHmcpMpkc464E7RJS6mX8+tQizV6zjR
z1nlEf3a3wcNPCvLUKtcKcFh6+X8IUUtfCKvPPKzpoYHXGrnoplbvTjyqHydOQVv
i0zArQabjjxaJ6VGQfEpXwcSmJwXB6oilND7wpzFeM6aAz1bhJhSnCgiUTvQEIIn
y7hJyJHejqcNL6QpZk0+RC02hYgCi9Cc8KGZkrmYTckLfXkuEhvMt8V+zx0+Z4dF
iDO/OVEzBxO0uQmxcLJO21jd39KThDLORC3zquohZViZQBC1xaCI69aNnceuyAxB
cbiGDupGywltD1CxM8vAgqo1AN1q6WPpsRY2bTWEsBv+dFNYP2h/EJMfkpPXSwJV
xmG7ksbM0ANslsliOrS1kT37M4y3SxRoHXOrpGPkFPygI3+ppyQeT2SHQTFLlYj5
mp7QLP2rlcsFzWgSsqNlSwx6kxFgN/kgze13CzzNCBC+pf8VTrNUc32O26TB84Q9
zWy6abKv6pIGEl+Dq97vxwg38FAp5w5jo92H8ADmEFv8XWdeURjIsxd8ZxHe2JRJ
u+3Uh0L04hzOvjvHvcprTADE6YMf52DvdftiYL9chqLEeIqy9ece3NKHlmElaVqU
Ejff+l9psUum5ayk3nJVL10u7sGGYOVPyXzbuURZaqPl8x1lQvunNt533vTzjAaq
6XHEaC86LdEQsAHuKZhTfW3Lu2YOejCaNlbczv4+kf373LeShqKjsd7QygKWPrCg
/wHZzzWsEsvhv9GWHY4hFKZHHz1mhC5Gv0SLbqKEsqYBR0ePNN/txK75fmA2I4rh
To9/BwHTrLavsob+F5NguwTKv3Hu7h1LPysRqkSjIkCKNmn6PsIa2UgGviiCsxm0
/s1dVdFVm/TBa6yFVAFwTOJD7WETic3YiukhrPD5kb88ZkGns3e9geMZDGtjvVp5
lkC8rUiS2knOTyDXw8Y4ZlWMEkX7nlfdFzcLA++EVVK6dDz8K6vHF+QIVNaFRHId
TnTt3xne4XqwUXX3LnZOBGl43YJvSggOqD1/nzkq2FtUNAZ+LPqgXmnkTKpJGLit
OLH4tsZ38C4qStt2+XT8bupZlNT+OZ+ok65eNHbs0JPZV0y42dgB7OOKWe4o5JWT
goYUR3wpX0iaxIrAj+tJsfMjpbE4AVIPUOj1lQ6D2YLaqFMuaOn4Qj4lWcc8LtRn
SV5wTYe0sPq8ugSo/bIA25YDU3RemtZux/8dC6CjVf5F72w3RjUtDYkIFfRjZRKS
KUSlKUmtxyPT1Gv5fUqa/vV4kDVlx7TTkvUNEZQQ/+IYpkw2sFIoVRBPgfR1HNk8
+OqhJvrDdMunQUyBRwxeAezRdaNA1617/MSnglADEawG6UQiu65U+9oB7P6TDCYk
99esG+efgo6fqveyYESDumeoGgkCqK79YlhjJz9P/+4Hyl5q6cx8Z8dJCWxpieU4
BicIj8L8VYLOfhL9twLQ4BNMc98idzNCdM7o0/321d0bYdDXZJ9OxRfZ0IMeeTmp
M6GQpyJiwys5r4VniaRUJR2yUSLqOtGTxa2GkpIHeRLh04z3d9LGdQHbkgHWAbKs
kfKbNEP51RCXqBNSPcD3zJikdk/3FFYa7dNaFSys2WtjVTVYqkN0NcYn2FS3L4Lp
KCL947q5fGm/SYMr7/yDg4SWmicb0apeTeCxPSqBF00=
`protect END_PROTECTED
