`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bSXPrT43XT/5EjGDOX/LWyD5lB9MHh0M9PFF7C6Q6ClF0Ca6W/506uMrdl9uXm72
2eKtWVkh76yOyY0KFfCr40BRcgpv2rRKhj6lOyP6SZ7jjfAQDi7XdO9CmPAadB+u
QKRf9MFGulyPxTYhsA+RC8zit+uFKGzO6yxyotv+WIgUjYlJjEATtoNZL3DcggA9
tje3ICYTcYD5W09OX9ETstLm+4wg53UsAu2meLbbzHd73aEBB0zJvu6Y/77L/sIL
k0q9X8/Oah3DkHH9HZXLAxtP4Z0RaIrLt9EfpIjwLoyHBs9NS9mlUVjBq02kdArA
qu5mu9vgzC2nA0wB7/KW3kyRrS8kIjodnJf2HyzpOXLa7x0vzkqbYkXxpPWSN/NO
2aAKbb0C0SYsNBWJRrhcA7vMnDWw6uOKDhuOp/kGFCuRHH47vPp6/5yKnG/EJeKG
ib2z0aN2QN01FkjyA5JYWOZzzzSse34U8AiAY+L/VayIk6hpfWMJVi9uzkRBDGJR
xMODRghLGFDJzsAJFR3+PAXsbVRqNQY1gbiMorryhOeJjAFBzCf15l+dmE5WiPAS
LEHAXmPbQcj/GIBdMfnuEUnslwkrL7vJGgxJr9DWYqOBKIZIULWCQQsaG9OYDTe6
yzw5eXjjsKca9yPCceMqBwD6gPrs14QxYPJhcZ7+mPanaVif3lnQslwXbRH1h6qh
2J75SGqZmxzNGKUt7mi/AEG7EgolEzT9WDDcteWjQbMXPydunxaiGtJYHZ2kubMf
osJzV0AmfExMIu3wuPMrcCJmbppARRcXeP5Hugl6oLmvtgzyQAGCe4cvNPS9xX/k
/T4WQHjH8Z86Te6034jLNcNki6J0anBAmc4HH02FqthnIMWxvSEICyGXGk97zfOO
4LNxBJO4AE8kLnFgyE+laaMKa/Ppue1QJqbAiqE78MlX00VkYSobmsYdk381DSf0
IKIDA4ZJLRIQ2lmzCfnZIRlSoUxEu1hsWSZlkGEXScHapdcLwps5WuWl3ug0SrVz
cQD0Vt2q++7cBpNIem7hkPVvkHLTNn0pk8hRsZ9RGHaHC+8xNEQzWbHXIybZzCog
TWH4Muntezobx4iqYDxuKU1TpA7KgdDrKgfkCn2tKBVMD+49fSjQuW9kY9LNOAvg
Q6kSE3/DNIjCZmaj7m1ocYTQyTR/8Q7ghWWTRJ2HWsxagcxQ+IpLa4XcSY4UyDuR
KbnXtHAS4fFJlTfrktgj+p2S6BlUi8kcsd2mBc4NnCVdV1f5+INpFkj+tbKfR8CE
Nt2i2b+fYAz1naAXeNjAQQF+OXRCTr19wVTpyz9lSdVEXr0wRnrcqPTFV7s9r0Ax
DnSiFfr6cI4hj07g/pLQEDLies9cf3hTJxtJ+qfDW19RGlDoQm7/j/h970HCFbQ6
ESuCvdu2wlDbvr+buod7GoGfYCFd4Jymp42+wDOdYIXkJx2iAHPKRzqQFDlriFrM
iNInxQVUHtpHmH6D2OVrQJwT7G53jGCUAN8UsP6cL3KvjTYFLZlAWspIf/YE6nF4
Awwl4MYetjqhKX6RfAC/+xHgF92+1LjEgAs8fm0akj+uzJmxawB5TpNPqxUamvzP
ASdiU2Ao4a3CrkyUhW16BLTIj64F+G8QcOjrGL1JpmQWbrQtHbWq+oSw49dkPrrV
lc1ulZvdn5356OcS2R1amWAMGhBqLUM+GRL8X0BEDGM/tgTTMoWaSM6ThsrPmFKZ
fkk+3IbAriq35YehgpxXDczQ8DWynuiOq5hWSptcDxu7DIKUmO3yqgtFzgRQC7Gz
APE4itQH4MGZx7en6khPMjfmEpDSGMVMIj2bP6FydEnvI1oh9H7TC28QK8GuzfSH
Gmq0OCBWa3NKzP6PARv+sMGk0dVb7LAHtm1yhLkx5rfhz6QABuZe+GKa/EdgaEK3
ZY+iLcBItaEcJOloZUVGdaOeKJwEHe0/1AhV9RN8dFDrBE0M7l0BWuhFsnwB5Wfi
oFHsjOjTWPbB8m2BHO16XuBlsWcd4xE7rmBP4cqsnRVOmfhdl9RFMwmdySFSYxgX
zhRtESnZSbN0LGQpce7W6TsJCG6cYmZzLsL/V8nbpmAFh15h20p3pBhezIUhQJpS
whWgNcnlOwalShCBA2W6dAsjshrmaG+S8YfiU1W7QN0DG8AARZyRqUhHODRF50Rj
bwUEGK6qUc4YZr7B4Nzxoar5O3TJVaKBlMfWAijvnn6nsH9NIioYgN+PNThMuxiJ
miXgKJsfkOAYxdiu5RxAcJH4HK5VtkaAXAkKxAC9DJkTKw8R3OD4uTTA45r8TAfv
T01pRh+rMp5Q9fha9vpywM5ovhM8aU4dA1NJ4p/GuCHhQAtf7/w2cqudpuEkIM1E
rc9mNBhe6WI8xbDXnE8zVlLxdxQL+IwBecEuY1ZX1NgLj8aUS/qOBDNgVnOacPeV
R7zVYCBhSJF4/WKlRYLKkUYI73SQLDU0wmxHwls/oUHNV6hNgvI3NNCythHYE20o
pBL+PqbiAhLA9+tTmK/I9v9PVgmj4ixg9u7kylhpEEkVCcwvWpo9q0OX3tz89hPD
4A07nfK0EVT+AhDA+UUPlc0FxGAsGfwFAm2IgO1PFoFRsZyMlXkM3M9E5R5iYTws
aFnjeRDhti/KIUFLzwRuhDsxbLmnl7vOgY3Bwe6NbVjh18OqKXR489c1lyefoaC+
KfUn4Ktg7nqicxtR8BddRDD6+3CwLfn6YJYvqsSQnjHAeuxDD9X6ADkfc+CaK5BL
GFFT6zYSaFyWPR9bKbTU+svfnXYwas7ItRIAUzhPwrnFTY7DfxqV2iyZksaGz0DI
lhu4ZOEug8EOZRnEvTLKjTZFKNgZSkY5Cb4F5qZaBHnPNcq7mKOXMJaOFlFFHenS
34W0re3XVxzof/Whn8M3O2ecPrjxygAoOUGUlzxSfzZkXZWdrjVq9ew5EJY1bDAR
eKkuHQVwzc1RzLe1zsCF7wCrjT7S8NccHrNpVxvzN1wptyJA6m5KQAhKysM4RPSA
sx1dX2YgXYo4FfnXmgqr/5ck7dGrKco3Hx60rXYJx3+uLdDsMAWXtPEoXTQSIuqQ
Auy0iIVxIoIFiLrEveWIKp1hd2V+hvhDuDoB5fDG9Ncejwqw+wwVfwER4mi2CKz2
9iEXFiFc5m/fJoXZ5yShTCgtwOiVVNgcKHTB9ruagZBIugOerYtQNiKCdbJ5IbvP
l58YajEHKfGMOnMsa0T0ldXKFSDWGmmlZMUquJhWcsCUweCpg4uEcsvlI+s1aGlu
8M0qg4OgEz1pq42yDYyK6+SBa6Hdt0u0Qop/elo49BnkCd0xqJ3L1qR/oeK0sbBT
4qPrM0Bf/ZU3tX/ZXBq9m2zmcAeOcGsP/CQQtp8qcZopcsgQak7HYsSCBfjzMi3/
eGp98q6E7NmuMcTwatgsZYyJapwbPVgZwA6zkUbX1QfMoTc39/MP88EVGa+tVWqy
uRjLDAlcEvsEVr+z1/phHekgi2qLwhzmThLUGDR6ScM7lKQmNISQaD5f3C6vm4n+
rgz8qYHjDvuMZOedPHVUBlrTuRPCOlH4oOfdWydIjOwwNLAAu6IsJFHho+x2Wi0t
REmJ4uVCpVusgr2EGz+SnIT4D3ec3MIp5UGFazcQJiqlUiOlS7WwMhwEVqc9nv+1
+8w/Te9t6Pybc6t6FvibgOQBt7DBKxGoMIhvDncz+cDdw84h71fWiFFg0k/R5leU
iZocU+vDVHOHdEzKGjAyIEdlKsI5sT3kJP7ESJUVpQASFsgqkMo6WjuJ0cnnT7Pz
fRZLvc01CPtjFI2LQo0ClNGMaV2p3Y+IPAdRnOxjjnYTE9b3/W9jntW82A3rbAGw
2Q9BrDy5B/Q6fLAztq0i00iutwpuGXN/9swIkbOblo8/3p0+6CjqDeTDPvUZoN4P
AY2UQdxrOnXpOFYk1+XHjZH+0gVgfVuCmOeaRF9YtElh4ycweClrYOZKQ0QwL7Qm
D+NbfDWFtWRHEkpGCnzh+8Ms86g/ShgcwwaYqFB2Szzgu5JLtSrN+DOIaOZShRlY
ZluoxEzKiloC1hoihYQpF9488px/OvBW1Ao0hKCoCjJJglSLCBvkuOJpNo9vQQAo
Abz9dqRQ1OjBDbRD68eBZnEkUGQtoK7Ul6HR16f9lAv+tXLh+zyTVHxnd4HlzJES
UmjcoxwQFe/CzM7WbHGx4XR5cHIhyDMFyOjopoAFGOvLDSRgJjMy3fQBCjM/Qry/
8FGPI9M4LzlIG6rAb6XnQnEhHcNvZ5j5PyyeNje9qCSpsGQ33NWHYrPDZwDtc5TI
pPYE9KVn/HDPFjw5leH4E/CJAGO+AocnKcwouhOc1E7nm3r7BBigo203oIrqfI+B
vC/ra00uHezgdgvod4ml7rIoRMpE9pVne9txa3oEJLoglCXpprP/G1fFTJNpwQhM
QEgS2DCHMCjvUrVsD/RX6SKXyimuyFFW+kJZmMOupmnQtBlpxe3TrwrKqX2J/41R
XwllN3EHOErs95UhO5icW19fJ8H4gYOxqMIDR4vLCGT1QTbVNZnY3/E7xvS/E4Yc
9zASudUrFPBXiHmkjeYGRE5NLAObhh3i88JJnL19JkVLSRxf/kufc2nw8a4yAErl
USPBJfjyk5CsuvAWELT3zpMCVc74mZMJkDLJuQ5larhhl2DrRpzScwkbQQjIUlr2
E66VlVWggGMD4rtFzB8AU4DAnoRcvtQ/WEl+auTlR7uogEewAmMhZTCnOeyznnbI
DwpyOAoD5qhWZZIUvZICTjs85Sea2pYxXm/ZxdQ9apFLIW0Vty9A4v9agHDhzP0t
X89ilCuvbvHPwNmudsUF6S8VPi4hfciqkcOg+H2g5XuMmtzik5qqJleHbJsy+t5v
/wGVByXipFY023gxjtttQDEMVdDIbY3QGIH3N99ZoNI8KJlBPd+O4BoUuKeD/WHf
1f1jI2Bxf42h07rFQPxh9leZKjIL2hYK9zmEnX2N3eKZB0Bvux5D8LJ4fr59IAqS
Wr32S6pEkW8gRTglPt4vTLOTEnh53U+w53awST3PEYUWYVfLPHwa+3MIYdc113Vn
2BctIhnaqLAsy8M3f7Fwp6VDQ8b1LxGcVqJvSKuPxzdARpHNQqhSnDRgWhfvbjcw
52mbzcvl0cT2pxu9odAk208TpqRqh862OxZioJLmdbZpo5OannLiFGYEYtvFW9tJ
ZlBYwU39OCPUoB5LKP4uIFreR4cqTqyNf1FqkuTo4nVKYm55fxHKHjyoDdp9vUhd
KZp96XMELyroTA8I+PzrIgYGTwg3ftrkq2KwdsDKSQb9mtlvX+v2qZBhxod5mjKv
lS9EdO0rKx2P1XtjGxDc3/Wvl30wV42Vyh2vk2Vxl2PiisbXq+cJdzSKHG3H0o0s
jmi0/+MKx32Eh1BvgSZUyjyolLJEQk4m7E1vaIkoVniNwshKJT2XSYWToCdyuRY/
89zM652tDD2CcDRpsnRbFA2PYbXW7zrheX+IJVFhCcLyxsPlo3QIjUuTFcwSA4Fb
0MGkReaKUBIbNRS63K8ImPyWBUZLU9Ao1WNtqXq4CqMSnJKXfdvHHYMLi8OL9u45
j2G/KlwiSMuvHYsoNx07hnP487BSwohbIb19hF5OVpL96hPXe2l5+6R3VdkMfSEk
ToGGZA3xs4zFp5Ek/ax75vFRwWdFsF0IQviFOwO76/9fNyWVVrBSJLHXt4EodcEY
5W4fG6LJqra8go8n+HdAShwL3C+3ck5OtutLMCq7jasnl3aNW6hjdI44nuset43B
+xBcATN8EAtBFXzWsz+pEt6ltvh326zy4lMe/pxtboOFDXU8Vo2BZWQOR2OO0JA4
GamRU1BoC8/OTcIlAi+HaBC9xg0RxifYsim0ZcF1/N0AeZLcqgbx47GXnsuz5lm7
GnK4wUTA1bJ9OuI5SI+4I15wgudsYmzz/s7daRMSopORhd7lFxb6vhNJfHFsRWIw
7TrgfRRRpO76ZePd/ehMz1pi00tpkKZ2q5AoT3jJq0C8PkD7/TbWGAxDpCQj7hYI
8jgn5zWlN9OuJ4KbFt+B8H1l196GLBufO4jYh3mrLqeW8KKI+BuHxWE7jz5dl/Km
r7xJZojJSe91PfZysEAuI0LwsuIsOfAafSkoTub9R+JNK6H7N/PW6IBo+/+i8tMT
ClA7pkOIej655srkOx0plf+nCM+f4TE7NQ4LkLqhvll/1fwjtZ+f0MAEls14UtTC
Q3J6grxdLGdxFtkHACPMmFbtdOf27n8UkDm7JOXGNW9YGcJGdFMd8aL5q5kQzdl0
8ZCA8oIgZ0zRJOSNPzL/MtisIYUMHPFNK3ORBJSYzN9zlfdFi7sbWNfwrGZgw1Ap
AWVYdRWBfV6Vw/CJCZEBReHo3BclksbQBsJxo39x7ZkmZzIuHWbQgDgMAGypIuim
BDMZs8NdfRGDP6Nd6guf4C8XTRqpajEp+qp1GSUkcVnNHpR8w6pR4E0dJETPZ6s2
jcXL3kTERqXX3kEcGcw+mPq9wjF06QRCGmSTTR7nR7S6VfomLe1GR6+0xDnXvEkU
PB9cz70/MHTrHhssnRs8W1wCwLEtEgI+KpKC8Bnb9Ub03fpSX+mjkSyuTfmqfdUN
35am+BuN4ZGJzst6vkfZspoIlA8z7WjtsGC7Z/qv/FZfqOPnAXbLZSRSMIv8nIS4
ibj/O8OwZwojCQ9FtJOPX/kYbX13Un3Gr3QT7/FvFcLo/R8JzQu/eyEqN4cbFNba
a2SoQtWodFYPESj/emTkAYHwl9OiJrj3rPAeiaeaqcBWJAeMU8tV+DBHQzUXCvfR
VSLPxJrYNQN7C9QiMH0r9wVKqx9dl9T9NG/WIDficW1TLaMFKR0lUNaD3AzvFuUw
+KOoVfoS5UT2lXM6Qgmq/0o19s/kSGKEt7EjFBChD+p1gaYZglY7EWXvpeQxPwpv
LZJc2033hBk8JLknLawAiRqwO7hQhrAMxKg8m4HcmIiPtsHnwxGX4HZ/RZLaCr7O
3v2GMvsO6kO1rgNmB36S7ScFVZLw1RXkBf1303jZaFO62SLgCf2W5qB9GHqhvYLA
IJ377tf7WpfNz79EvjFjn6LsR7MLdPgnjeZVjz3h21AMYRgUJdl5KOfnjH+6Pl9u
FnlOqDRWfWm2vJClHgX81RmjBYIy5hGAtshCAN2ZfPoBXPdJOkTYNDxw9zd4iIX+
bFcX6cahHFzItIbcngzxVDiO7t/g204ggSCBXDE+CkgXaPFIGC2A7B/H67tj+Qfa
tfL3Bca7o1lfJicLnOufBuuy/sUlOn1Q8BBUbHzt3f1SpukOvxAEN4vKn8SA8XAO
M7lK8LehCTtoyqRzrxViaBc3FWxlKO9b5CvQs27FArUkYktMMqNru3igk/MxJuYK
ZI8/gjf3Ng3QJWPqj1Qd4pGt5GY21chpaz6pOQgeXITA2HHc8dLXNXkuO21xx8tq
oAnUdZG42fkdxoAg+0QsBp+d4kWgzVRGyl8Q4C9Vw+gwcnp9G3ZuGAMBH7sdOVUL
Msu5vQt+PrU6TheqOUwD5BxhfnmHVs6oHRJOjgwXFP/Fa3fUBfMjRTOkhKda56bt
vv3Mh4PEVVzjecTkwkpYab49E5+VkEu9P8b55K5I9ea11wrp2BniHKbuLzCVQF/w
jL/UU5v/1wRtXOYd2SpEHKpQnq4323MUTfAB5qoo3RRCULuxikmaxPdLfGngJ0/E
LlyrZh/a2csLmGInGo2+YK3vfDW+ueAyUNw6dC3I5vM2zr8lrs7AI4l2a3fur2mD
RRWMcLDNV2f1IvGp1ChqbR+MjloT6MkLU4U13QcLFP9kQUAt9gPKFBrwPQRKOvm/
gxkRtPrO847FGkcR+3ZT3Gd4y+CRUOQBPfF1i0njLoFzuNBAkpCxKZbtDWEMD9+Z
+b4iEsq6EREOzGzvHwU8lnHOALC4n4S7/nFXbRgS/L+vCGIIFZ/wYnkYxaugWMwZ
n5hnGogCH3r6v57NfzLCKa7kBK5tr0qLcuqJ370esYlxPlnTCXKJc7Mq0N43BMB5
nkFcP2Q4wwLcXPvlgWdhYY5bAgZ7Z81g0DgnJ+ZBiNNi4DAX0pJtV9e1LE5w5hzk
lrpLoMqprubszc8gVAOrROodEkjc4dw/MqvYe+pvH98aIFuDJsoBWor39WrSIsfK
1k8OwUKVin97tqq96syQGUt2W4ybQHUBPUtRQpuZ/oiMKh+65NsrBeYefzUVJ3rE
2YaEpb2erI3U5apj/npTSgZkj1ZXzLZTguTP9gdfyiQ=
`protect END_PROTECTED
