`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rwV5AdD0NM7ji09ZETEYEsGQTPeUvhR5O/noxzCz8Pc7V139MXrZbtMMBiPIQfQQ
PjwPlds+kk2n6Wc8MXT5tWOvUMMY9c9JN7cDge1jh41P92UR7ZD/YKXf8hhOyq8B
KATnBym6TyhjhtU//1+iChgTmsuYcGip4Vc7GzSaoYo5yKizMUdzJ+VzQWDPmkbG
/QX/aqaGJgknQGMeilpV/Iq8S/xIgtjVd6oQkdDRWqpkGIfPc0ckvbs5UQkdlhut
syvYksgYRYVRg/8SNdAGfv5zFqxGjoqtf5OooIgK79aQaxjvgPAEbMg4KdjJpQ3m
tpxnfCjDBxECCscAJ/gV7jFO0CwYsQ95qawzqX4dbf/14nkT0y8hQvn6tCJnw5V9
wSjYJHtt3v/NvU5UvHtm/X/2hnXZlJC3nxNBrF+asu4t0jcgra1Cv2nbmwInFKK6
WCA7X2EBBRpjUbiuYljyJIPW+JfwnFpGVV45MTbf7/0=
`protect END_PROTECTED
