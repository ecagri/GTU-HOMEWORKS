`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r1DB2MIYyL8rdWDmp0xKEhqnqQCVKQOhrpLpzcYl/F8c4q8zKd2ZwudswW5KeBnQ
lySdWbQ8T1b8FIYInWAS/ZNma5WV6zGXwxYw/Rc2R4VxLk6MdTU/3hQXdVFG5pbh
njdoELSxp8qJVwTU6oiF36T6oWLsLbLhpOwEmUtDQET1tcgSRSjYUyxPGj9E6vaj
UlhI9asfi81jhcczHmUbUDKmdV9gTN3dQ8MuwfbyGRJxqUOgawF4ddOQ6E7Ezgkj
hvWI963jKU16Yx1YS/xT2QK8uZbzrQiK2eH8ZI83GWg9YKg0uzPxu6WHM5ZbVTC0
cuCki7q8iNf6VLFx4DY37vEQG87E6ZSLJQiI3m2LugDSs80u7z2A+8sCoNOjajWG
piy453N6bQ5nyxFzyAkGAsTcLCxLOh5R+HcT5AOacSRa3aBnUh2jGY0gT+zWpEjv
Wqrgqsti7NVY3A70E/P2uVWYRNMwjk+hNUCELD2e2nQ5RrIhZNuuludjxVB317Pg
sU0zysZQJ9gfjqcAyhImimqNqqwI9UOYfJ8C1Vc1oWsg6kM7PpC7aRRn4zdkWjWT
ZMGaVHQASXEs2u9Bk5ydm82cYykuvEk7oUgZE47JVVn571CH1FFeoZ5MiXa/VTaF
5ephIoIw+Z8ajeuJqeC0JBQLrfAu8Lg9T5Gbk6vFAaWYqlOkfzDBeswMLgTZcB2M
WplU7PeFfRkRkO52Vlkkg+RRXCNSb3UrWhmvfp0Jo42BWA1wBxmue3CB7cUM+HQH
8hjsWPBJVlofWBzHiBqvr3r+JukN3PC/L7T4dhQATZwT04SzbbFlTxsYdIBQuToF
hSoy63j0CV2icPEN63A3E6zCTj089zlZ7NfLGLWVu5W2xm4rlXH/RSFM2IcNj9yS
d4+lY1Yq+zO/QROuGHjYwiBN48tuJ4e0qkFwr5X869xwgS0wu885aSTkOCZkOA13
Wo2glYySBxVRTdsuhg5pDqi+3WSBLv4WbIa4iYzsfrVVtf6iPA3nvb/QHFN/1EBK
6a+cbzyPc5g6R59KH7OyL8mJskhVCovFFBgW9xVxIwLw6B6qKhvG9VMkr2U3kCw2
9Rz18+WlxT+hi1aizA/cuZcrW3XDP6xO1YvNDDICzcAg04dX6H6MZr2tB49shwGM
ij3gK0jFGsZfLNK3RR4CBq5bf+cwAMxrFKHxmw7fV5tsCQ9GCumvgXFC5WYRxGQr
rThZnvgIgyCwCNJhqJBy9LOXyzvUwe0As3pjnX+huMs5GWIaG5zopa72CoPuH7Sx
n7l6b/k4uf8C0+sHgcencNJsnXfX61zGEOEAkrPemCpJUV/EJxS6h5tJiE2qV7PC
g0g4jxnZHYAZu0F9bF0RjHOOBty608Gnl75Q4KsWxqF1QNl89WHOauelGvmk8dF4
XsFyzT/Yo52MexCfroqTZQ9aVLAAqo3XtlZzRlWBSTi2eTvWa7Tyw/8fQcyOG1ah
5qPJALPYK79Ydk4MLE0wRkP9JR6DlYXI/QjQSwEbvGIuXOa0wHtTN/4miLtBEHPz
c0NtqT6lMW87we4Am9XaQ6ddDctEh8hBlnF1wYjrm8oYBI/zjNt+rGGoNp6XAMuN
WtcyFD4urkx5LoeTD39c2oxaDqRMbeLXBCsNBTQa3f2SKwOuH5WvMCb3KSWcBPEJ
1IoZqnrSfIuPH+RLg0uRMXrw2jUQT/mVWfHT2fBMTMfhjHE7ZuyuFQksY5nageqw
KEkCj5UBouh9DFCwXvXoRwfWyn6cuQ8yWaJMLXGoWwwLBjXD2u78pKOhHmnbnk8j
b9EVotJp+ZxSLKomRtzQIdnfC25Ku1/8tIpNZV4GuADSv0Vz4/rfVS0SqQtxi8KP
qRuz57pZHrq5BeL3eN4mDwEH4hNXZiFkkU4wi905XW+XJAXE//f395CklAgA+GAg
XEnobfFOuJUMXuHnGJf7sN8t41KzcO1QNV+uhX1BdwlN54ibamJRwgJi/nlGI38P
4c7D4SXVo4PaTVVPnN4wGqFJOPJnyCtOVhcy2Z93188kRFwFBo4VpRq2y+X74yi+
2MsNBVQyE1MvC9Llqmw3UnQozLGHPKgtdlxpwuwmz/sMyGax14eoUUZgEFFjbNQj
mp3sXLnP2B/8w4ARrmci3xd+TDu4N0EzJDhRi0Plqve6t+qgAK2VkegumI4nWf91
5vRGr689JqO5G8z+thhCzn980fvdlWT5nAnyBCIckGphjZ7UBNi4djeldfjm71ys
XENHKJ0hVVxZd9MD+R/DK3HBhWqQy4F9BOrLtZ4R9+FTB3WUx/TODRv9oV1bNen9
Z3rsALbqzKiXnKMsGUwMy9j8AftDKShY7XRriiibsuZSYE/dzQgfBAAVK22WKyBp
xVCOGm14R1nqQwO800IjBfyIQ+TSOLXvn/QvPiKFmLOKaFpSrcJRnE38zgNKDmeg
VxVYu35alfYxM5QFgPrDixL89UBOiiiyPui855Uh6yzSac/oA3RPmIaFQ+tRtlvI
8qx2VOuIro47ENaiJ6UdqyD22LGGPACcxeS7eQVaBfy2iAaRhkc75fv1idE6DYXr
IkVjs3jZjx6Yk73T9Bg1MW1eOxy8IGFiGfzmgNXJ6TvgsRm+XmMLRaG1BAame8iu
LPvjsjUtuFvw/2B8r9t/a8xI3w/5iaogEXs2qs9UDon1h/0ykzQVP/8d2IARZ4ZX
d41mzavktUjIvvGAKGgCHtae/uRXk1mpgySITF4svL7I8Pv5BeYm5d/nurEbiryL
6QoR7WIO59A2jT3dNLP3bsFRjKeaWmVcaLe6h4NT1wZjox/SSvz9PKYFEC+EIJTO
MW3NV+/zA3M1+HqHzLKVzVymjqtGYL83oLpdd/NogtYDH2Z7qfhSUt5SAyUpF8BQ
1VxXDAIaQvlMhYxktiCBcYP77adaSerNiMMC37rvwIt/AXkiw6giwZ/er355Rpnx
5AMMoNHOvMISLSvt+k9je71u2OE/w5aZlerbRzIbPKnu7ApLF57II2lLKflc72uO
j+O2GKaft0LVuqBfNhBQVo5gITRAGzP75puHNS/4u3rj2pRzSywb2OEmPfUg49Vn
J9n72AOclrVQb3igKcV2maV9MDy89RfV+J8fwsr8WwJxsfAOodN4GowyWuIXcZvl
+npiDOTUuY+W3VLwEc6Tytq+2tMr27K30fN+mkxYWuPIRDUhf+/srKLJXA9WCY9d
JTt3R/kJkaxOaTQYA0WMC15DjpQMatlwSLGXn9hcHVePPMoOhCBK2mMN1A6YAP1B
c9j0UjUlR/Cr5fAQZb0nK/b6R1gSsFigQy6+cv9roA31C6a4r2uWcmynR/8tJbiI
Rx2/olxA6f6vXftEkU2yUWWfUZLuEssaKjNEQLcIsjJs3KUbJ5fny8dEOFNOHFUq
CGK4i5mCwmL8iUW2xG/knR0pjzPGv8calSAUANZGRcSd0qFKJtyc7QKFQ+PWk/sM
jT6XtRFoxuKGakcTq/epVJMf9wG6qE/PT4aBM9iXaUNNTwBIIc9VAVDZ5yc2QbCk
3+X3EJ410qYqvvKt8Hg2Q83aiHkrGEvrZcehNiW5NxZ4oIsW4ryO/bsgsPi6njAx
08KDiuDX4Po3xSSZegfWdzdODJ1UxId76R+A+jJH8CX11J1SPihxg0OjvMAwueCw
kxNMK+GZYLc2bjgNzNDjDH2Qx9JtE1LqWuRiGOGMgCYpf8m+mcv0n/QH+yRuYGBy
x8KkV+BpHIxEjF7oy0rFH8NgGpe8+J19a/Hu8KbQG5FU5iI3oKCwN1i43Tddpkzu
M49Is++pZpxfwkx4+sNAKYbRSCPyOzgY4M+aIdBD3mt4j2A/NWaoPV3lGnWa/r0d
02BKaPT0drmnp3kQr3THghicShmwCeJFVm06C0NRTJQsvEImNqQi+EujjFst/CVp
RGdm06cw+AaW8J/1uBKfaApwrLEakBC474/cq5p5dvD57jPBAHkssgd8p9aSutqp
wuGRz/fjApqpMeE7TCfIYQYN32MbscIDq7TRld2NnUeWhIsqYIRmyOYtX2f+7k9/
McBKJwPPdzCps54rlhy5CQd5sNSB//hZoylqGs2tPJBEPp8n/xCZ8YOV+EM2rrZe
TiQCqO29tGOlV0dzdEetPLwnMgyiLezGc4uoDFto6IEeJ+LBJSKO0K9TdTPWRyXi
sgLT4tJj3MHDp694N+rwi1jniKkmtUtbXl7vi87KZEduxgOq+kSMCZtYh1qHhZ7g
VMBAifRRn5ieB30j7WrxNOTA449gJk32dQp9ErxnGg+elxAFBoTyDSbTuvgMR6Wq
C+KZMMhsVgza2huEGdPcx0w+O0MeUmt3KR7KUpYtnIPzTk1g0fH4Ut22zBS89beg
XnGRbN4W+OaSfZ3ZBdQLZoEzeq6ojElmnkr1XqvbegPu7O1JnOd0EeDswMuZ5OT+
hUGfUOh8uyIGXecvHehiIHev+QoiZzP5OHFQ3h704wEXHjtTph2v+MCxTCNvVxvF
YnY2ZjVGx3htQtSB8jO9TpAYQ+oG3YOVx5GlDz20wLfkPPzkyLLlIxwpq5GLXqOq
4HZXu/w6fCMS6EtFM/YWOVEfpjJv2fCOghcXEeKVbZbr89cnjLRu9eTvtx8Kbw05
DFW5CAOf0AgNdLis8mHvGeKGd1JlWF2t214vFC/QPe0pviU4cAK9302AanpwE4Cf
k3X4my5XXkWvAj3v1JDTKiNF9Xw9PpmqeuujfE6vV0M=
`protect END_PROTECTED
