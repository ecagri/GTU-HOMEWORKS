`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uxFTwPgjopx8jv6GuMVZosEOyfQXZmguvuwGiCplbAgN6Z3l5eu41wgN1xhXg9mU
50YZFMzOuBRlLoaOd1tdr/ppozLlhnNWrc82cZaK1GWqrW4tyMAuzsiy33/VJs2I
50h/FpFS0UgSc177Tpnup20ykrvphTUHXvRRed+plHrQVsPdc18p0IsbJZ8O8JS0
+ktxEikwdSrFVAdvFPq6RyHYp0aw4fpkagUwZMB+ah0CHYfW+Fb3FPCtreu6S4QK
7OTgMo/OrJine626JgwPQyhA9BoYfOTPemNLQ6QisJhB/gzJD8TXvtJY/KkYvqu6
CNhzbIhtgcnhv+5lDCI+pTg6v3PWgDTkpJAn5ftwKm/eu9phRs34kQFqJn2vqM3f
C7TLyJi1Eo0HedPvVZbblXKQKlK5flPrgKlR0S8Ub/KUKQ2Z7L6d481CECTDqsH4
lyhmrfNWk96rjoWoaxKbKcFASZeDm6ODq0TkxAVSAvIHjKFW7g2duKylnTc1/UOS
JgefxPukCTFA43zmKM0SBed5/KHe+uSBtDgIZD4oYJQyYcNZ5x/wkwIbOPnQcSw/
Dj6B79bTw5Un8g7LW4U+bFjQpV0kyRlxWjVOyJZ0KgBM/D5hPZJIz4dk9ZNpRK2Y
U9SsQeDKjovj3LcqKyFspgI3ZD+kNyEIbU9mEnZ2lElnB0GcQkrsKurakzTsAvDA
jBVoA7in00xbWcfIbjvZ+LN8/FslvmjC1xv98ty6snwQ0f443iAL+lvsHpTr0NqW
5cps+e+/uNyiBCx1t0nP7qZLRuEluMzdOOBYi/ea+sy3EDnSzqif4KmmNjDfBBMm
u856yVl7ALH6H0kZoWJobg==
`protect END_PROTECTED
