`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z5y258E1i16EBIBplO4nVqdTNQAOwmZzeOHq5CLhFSp8PQaIJ1q84Qf9aTXpKTde
vQ7d7N5St5HPYQluNo0I5ssXN07aescyx62JQxCeZi2dVGD3P/UMh9gY4ZFutV43
bfPjfylq4aCp6BcYHxy/oF7DnfUWzmfObusxCZB3ID1ZRJABS7Rtp92bmhgmiom4
M+tbTGv50Rx8+FGWSJiI7WcRn1+nyE5sP3EVSk27TH3PXrN/T7TfWUmS3IJ30eWm
ff86YtqxsGB3X7Qi/Yp31EejGlA/g4FLjS6PNg6NQihB5KRJ8Hi+tmRtvbVOneFu
U289T5QpQwkfSm8Lao6cZZt/t7IHzYwt7GBuuA86STOx93lihoQ8U+jDwg+W9/8v
AyW9EPgBK9m71KbAwPclqPM+1knWPsuuaKOhqnMiGPnMpUM7KJNfm30cnXfjDoMM
QJEshNdNos6+CQvQVLQyYo8cdsVtyyB0t5KuYO+VSP/fghWdE9IwVtOniIrdp/zj
1XTSYrCHiVV2dHWKgrnjhfpKQ2THo6ZP5Y8Gi6hDn2mYxxLF87zMCtks96N8aUcQ
DE7GyMu+9kTGBxGfKhyNBt+7ulNtZieRo+OdL7fZINaWSL6Bh2kONVujvsIPtHdc
0HeXZAmZjTWnwsKDrX96b8P8dZ7vBN68CucF4WASURwNbD1fztSO1q6a9iQmRk9P
BZJzV4nvDCY4J+ZCkChcBX064u94Vo5UUoiofwgNTz+dRmjQCmN+v4yKOOauRKSv
R3J25Y4fvYSx2sVoCIJgsHNo6yzLRUo5coCe10vX/dCjlhKm4rEOBIvQ0XZcahel
`protect END_PROTECTED
