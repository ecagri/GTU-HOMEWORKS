`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZPOfOn2clLsGHxRN/2u8khw3VP5rHlFM6WGGLUtiChQ3D40zyciahdhDwoaqEeaP
QJrPsPMzzpbcni1MU+rs6ohT5AHMu0xggKUJNxtKN0hZJXlI//Fc/7IYiq04M3iH
yHCNbDoi0Zj44UseCpyCv6E4JWfXNq5MG+AdaFMwj156VzRQm9B3Ap2u5AtcKnFU
dBhq23ikSzfcDyMhhqt6oZNHzZtcxU2SxJd3ECqSiggKkxraWVmDpKv6YRhB1MO1
B2RBVmUClXFxhgQJWn8c4229ttzOAnHChEFvBl2L6+i/bKufyT+srBY+UsXsKgSv
peJZDWMh3lQI6cisQiuimWWKag/1zg45zgSOqZX3E5+QEMzAPdZBnFWDftkZ5MnA
gwD0k4E44U77OkxiKgPZayOnbbzr4czv4QDYoGDkwQjiahoEKjNc/wE70JCqW/f5
yakhz2tsL3Ct0zo8lW6cDMqd13MlgLBsAupH/7ZtY/gsieTM7UTam+gvKCMMo9wO
Hie4zHBFGMN+L+ewgmxy/xU3zDYUMFtOWVrkpH9vO+ANr+FWUyR4vcUHQUlabwmf
LMqLJdpx1W5R9ZIWeya6bXPa+WlrdZzgHMpZ7dhC5vgU/e5ltbgqU1lI+9Hxv3hz
Yh2SCkcObDvFTGGhtxd8egXoxxUquu+3h32xxbHb8ilLjM/eIG5g9iYJH7JB3vff
CcGb0QCQeiovEaJ7cj+0jjpOqm3lN0Wr4sIw28YFxJ6/NOCcL0winAUXJmmuHiRA
jeOEtafLeOnjyaGh/fbsn9It5Ls+aztq+L8w2Af4u2RmzY8LygJMBsU1uQLircIG
VPB4knTD0Z20tstuAEgdtCiXxBYQrx7X0xeY5mZecxN8nMbMAF0YZDQpVte8X+Pj
+yYgSLVVsOwf11Fyzvua6tiwVS1ZBAEkf2RuyYgHovDnL06vD219WtNm6Tv4ti5I
l0qG/ePKo54rC38Cblw7Ea4K6/oN/XzKJeFTkkWJF35pgONM/oalG8ftqe6NWdqL
b7z6dyieVr18R219hgzvjWEUPIIH6ZCWkla7EhfDBoOjfiEv4w3fHSMx7/GgMSL5
YLSPJfGzo3CwonDVi3XI9xcj3z+c7wT6LclEDLl3TZYV/nn+64iycuQbIwA5dCYW
8KiEDlDYVtF9MOP5HVXbwdVnlFzCzISsIvn3KNiMy95c+rkp6VKP1ZYjQ54Z4pui
EZiZDaICl91cWqrWe8gxM1Yg4asrSHz0tO2CWKo1r7Ul8Wyg1odRwHW/Brz9jDJs
SIdmQUDT7VXw4nt7M9Af12C1sTsGBE77WOFEBT9WSnxVMtiIDUq5+sMGJn4HZTTd
r2SkGNwYLJU6fJB0eoUu92CwQwzYbsCUgZiV5rxOkhtP2ZadL/6D6HV6WqfsnlH/
vWCa/Vm3n7/eemmU1R9R+evzLNZlyoFeQIOrddFdQPgidx80wSzJROGgZoExONV0
mZ2w302viwH975m/i3TGIB19zeq9p3gAYqNSq6TTde/Oluk09aJ5n6cfgLo2Zm1Z
ZnyXey217xu0Sj3p7Njh350rBNoP2fEBtV83Mesb89o5rHhSIMYE/AXIvnxcEYXm
hXIc14mcjG0fBznScCBxChQBo3jw/vPyeB4MT2haKSc6TILV16mGQaqnlp6RweYD
yrPHQIgeHPZ7r7+Fr13M/Aa5FYJS0KdaCJlVEf5uD0wood63uLkWzi51vzV+Zjjf
nZUYfcK7HiGAcKUqdaBrAg==
`protect END_PROTECTED
