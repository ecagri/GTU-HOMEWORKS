`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pyd8RCZZDEW3V/ju4Hha5aE7qa1L9QdbzNeRTNH4VAM4EGRpafFBMNeI7i52xz5N
AvAv59KCHtoObDP/YAKPl6dvz0vTZ/sl82DXTG4ESv50IBv2CeRQFtJ0YfN1gxs/
73/Wu3D4UuvR+W7A7wBNpkGJyUamXzLlAT2sIqjuG4ydJo8e6+MRNCQ8SA1HY4fj
4WHBkWP+3mUY4lwlUw3d3ZWspwt7R1nIZZsWYgCz9qVvnlEUKGrDjS/c8zlbzLXw
RfVHKuRWun/gmLLAyUo/QvvBMKMJpH2FLktUmG2iuXNrmLwj24YGYjLkCJ5zDqxO
ojaZYtBy8v0wd2gl3XZAU2SKoqkdVpQxDgyNp7KzS7Jg7dXIzg72oFLuS+x7+PRK
bPa5b8zyqlvf8saIWkya8QuPzmAfB0sEbYDg/GOXYhSiNSWAAxhAV+iIDvwWvBjS
ATU3VvlSEldhIX1G/caFgyH8lUM9pwFh1jYSpPwTYHynGaeG2p1nmq6abmKROzwM
sxrQmA9QpaXGRPuY1lNxjOEmIUw5TUs1/A+GFG6PvwiN4GjtXkgEeTuuFDqZwo3D
fDCbIFjDYsiVLcoJlojFjj4L/Z29RsMdYZsQ4k6hNG7ubz/4wccu6jaRKi7j4vtp
X4JhbzW30q7VCHIyPgBUJ76zAlHZ3pt3Ey6G0PO/vGqxqPfEDRkJEBJQJTYJJ3GK
CuHJ3NtiYvac5EEIuqQPkCBJbvoRV4z7Rxv4boWrG8zRxs5zcl+MzrG2sAZYniDQ
u7ShJSTVF5pCGLf3/A1QenljpSXyMLeki08AAPOpjfQP4qN9k9nx3/9nPM4ATDJl
BQWvZ1FSHAknaRMBDx0l5umgqUWlPviGZbqFGElZZpO7oeUd03ymLuB0aqqhbxSe
N+5z8QiKE8JmqRyWfSZtS27NGzVYMFZGvntmSDC0Et7mdiAXcRboF+vsrmhP8UNg
5Y6bpsBSCAtg3SDCh7W8l3doKc5XqOOCGiGCLuJjxTFLiKxJOdvzxE5AQ7V+ZLlP
Q7ValkfY0CxE7UbdfyKWFjTJjXr8NevRVknYo2yVHCfmQJZlYOektRwqhx4kxeiZ
CPTE1OhwWJZBSEKDA+R6c1upZ8bmLGgn7KvbF1l+WoepOi3xmMQqw0Uv8+hE/2o+
iDYPtP4wJZxaSim47fCxdEbc52mW7G5pLXv6AbwMRE0a0auZrLLGjokVvlYXFjd8
MOLglwEelcUGYYoTLonUxBGkgMa750ZEocC4aok77foHDbfLmU8I3Fy5LkeKGlH2
nJ3X4V6s/IfHZCQqsAjxnktjLaJ+8WDxONereaLkEmoiV9llakxwGa+BlANiX+Ju
k9+mma3Utj6ft1ujiRO/9ggEp/aUYx8KQKmZ11L+Sm9hce64hznQjhpw+0GE2ckP
sc1SJAtOJ1Vn8Qa0As7hKIJ+oS94fiEUkQSxoiyHRCYZ/pVScmobWcIx+Pic7Yqj
/G9LHVyLqUJU5NRMor3QgONk0GPQXw0GGi0MA13+/ZAx6Y8EQ5Jt482pC00rg9it
jdiiF+f5WuoMDhjaY/vh7RprhzjdFUzSa3QHU1CdS9RVE4cHK96tlzKq6fpsAYx5
LO5AcXwHqSyyr2kJIXO7Wz7UOXTumo/+Q1sxLtdGu5eUrUXheDuX48W86HYHP8FG
ydtkRAbp/VHaltrpn5569gIz79rjJTCaNopcwD7qgX0DeYuoOKFhijaNcfWY3PVR
2gRcv463bOI6+6ty1/ldw3ezhQmzEGwyzx4YaDvLZRbNsTNc6DuO6y4dnVB1BriK
jLyl718pS5HUVkTiyhQfZhTRTA04+cucquYPlBuPJzabSDsrHn+y4i3XGx+zOtuc
+AE//L5xQ8zafyvhFJxjU/M7RtEbX2/vW40233NRDxMXiLxfmijQ4xDdvsaZ6yPL
wMuMLdhcuXXO8scM3lVbOE5DLrspX2TC3+TclEfFeLOkN3n9FlwaqVrkRp0oxES+
oz2uDVNogf3RO30N7giamY0DvUhHpLs2xbMLOAvYflxdUbyTH3wDu75cB2sdS3iJ
bkifkwI10/YeqtoiVdMzTad3SSeMF8gRmC1mKfDjEdEIbjZv6IOio9AmKm8/bC6g
jvS4m2YY+EhR0nWlQxXF4pm/mfxFV5BRoRZKMLffgixx7TqI5uY9Ab2+9nwLx3lA
rcw5K2u9AIyKAGs0OEdDf8zXEqy3ig1UOyAGT4NhJrz7PfWMDvw1Lq9PNv8q0eIt
gI8eUp4M1QRm/+0rOLWFjp+707heluxnJB+ezlvqi7k/Gb1X9fgXfl0GchSkHbTZ
TkEB9nM8FBp0lCvfitOxumGgYgOzJcW4aFDXUSYFyJHJpG21BlWBu6nLl5KkeNeV
hQBUkH88IV11ea9RRsz+NtarFOcAIJWWiR8MbsdXrmGUDbSSbd8LG+c2KUcrVhsA
7xIFvO3ptVXtJ1ct7c1ocvCItLkKZ8YtJQcyC+GwmMXr+bEvzwj7vu5YkRZeaKAc
nVjmqmkXFlaV3GIVkp4bPOeq0Kkmh1ja08aSuDPRDyRNqszqwd6sEf98zSVK+/p5
jsuMMK9nRvYJrdK7b6ktr2wFMHhb6OQAqkqI83ZOiFA9wZNvTV+/in5DKu35IYfc
InYXYObB+hUid6dtMIGcacSKrpoyeRp6CcrTKeOtOtk8xzLjctq7Kybj/huLJbrj
GJW+xykm3qzw/OUHWX2XEVY5XU/CeGRe5hfy40UVkr2W7PT/mh660ibXdyPth5+n
bT9UmzIRczHsVIOISaXqg4LA0s3al5qfKaw5geN3AnD++VGaCMggDHvs/Oz4Xl4W
XAGWxT5O07GP9XtJcsfeDWRfjRdAHpn8iHuRhO6veB+iYPa1BchfYjPmx+mW4PTP
6/3SCwbbElEcyLJFH5xi5ncTv8pJb7kzkNsQo44tCdB+vixynErownpzZ9YKAZ5a
pfMd8or3exFYZZRG+adrZGc1x0e7r2rm2hikIomc4o4qjKZ5yF8CaMImobhDJgaQ
mjKbIoJ+mgfpho8K2k3ztXQwNYq/jvs/6GHMCWnq7M80uEmSzwoj4PF+0R7P9uJa
trk3V214b5JFPcgACQTvZwP8wg1CwG+ZufNTtrAO3TJqcZbo9XUlttaaiiecl8Jk
OC3aoU7m7GeG+7FSUhH1a7hAv9X6kB5hbcwA3O3unhYWEuMUbhemC1ZXtlLyUP7n
XWf1Ok2Orxqida8LiNQlUOHKaU1Rb7WoJFXt3y/doaypqJb8KOxus2T7IU4V7aob
VOHK730lb5Lgb5Vqtv2IX3TBCEHjAsVhLFrqO7QQt8oDQVbflZejePa5Y9rwKVH7
vYxvSszbSczVDaaC/MwI6/xqQQBgFaoVgjvKD4yHUM/cFWLbqcV3fLKFkR6t3Wze
vng+ZI/n3BOniYUzWwuqBjOCNn90JAoNxGfeSd5JJGOul8ClXKxCEBz+9LoJ20mA
Sp3qDrjU7XGbPXIlhqNI5Bptf0p5lWZZLGE37uy2B06Df0SrLjZ/uqUEgLQ72XKO
2MjIMv7hLl3XzmlGDLiP8qIzV57CnzSG/3qYkqxgh0GZrvlSOUS+gmK1Xz0IAgSx
HzcvOnQqk04M9KkOt09BUQcziBJUiNa9+4kZ29G9xkwVSEiXBOcJO6TQfes0NIJX
JYtoZenofUMofhfUyuyOksgueqKagrZEXKL16YnUdadsiT24gFH8VJfJfmyh0NsR
pxYTcGCoNNK9z4OIJaNUebEk0bWQDFAzko5cat3IWly/2ra5UO64CQ6YJVLsJJFQ
38Fku/2WRCsejYsFiWrEPlN1zIdyiPk/D5VvnqlmYa34gH33/nSe34a2EqcBV+UP
QPQjs8jvwnbcpn64um72yuPr/T1/zdAUjTzolIYw4GjBvCprxhgfUiEJQypZJOfn
T9Hsrlg/rgnp6M4etMrIVqtOVpyy+V298Te4ihQ1QFqpa/+l9OmSQmrK3zIUmEH8
gTmk/8ZVkOA0W7xEcASOk2sd+et1zZQOTyHYrTnrQUIjDeEVt3PuBVhmTCJl4UZ/
04ZZWqWByO3PgdIV09CQ0epXNAW4c46tPrvvA2+AiGZCxtlv1CJ8aVWsdbJuBHyP
1dEjz3hsww/6IqE7rXGc+3Zi79Tml8QR+PLad5L3SZzK1fIO7IVUFK44Bm/YDi6P
9h9ZB79SjCqdRBlPTh2QtyZGrasqjtSXHLl/7Qu1sJHWVdbrK4ByldYdYkQy+Use
VW6tA2gDDstEWOVT9nZOsNKkzCWd389UO/bNI/JW9Ijd7yA62iePWUQXysefgMgT
yp2oc0yLd8Om3TImgM2lv7WyGotVSwLuxVSHP4BP6wOF+Igo6a613EoG8Epv7qtE
v4q/RpnbJ6jiAuSXe0XNwstB+2qWNZFzOqf8XLbRihybMyk25ZPBITGdjL2j9t+p
DyzrjtPSYNzpz7Nsv1uYKpIku6EOek2ckeCegP96eEo=
`protect END_PROTECTED
