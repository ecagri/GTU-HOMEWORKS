`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SR2rCFgOsY98c0Se3nQkxIFEuwCdU5FaTqtbK+DjC/5zSJ+70zeRYwBmff3eX2eV
qrQYfPlH5T6lPS/IdMprpPtgrtoud1IbYkw0gm2LlZEJ/AbH/GhsqJ2Ej7ZdPuEL
SkDkL6BeFBt/huO9A4httveQOVOG6lItLOJVIHdj4/5aCt3tufTlVWj3IDNSqawg
mMUne0kdYlsY5Axt8NktFyWhud9u6TC057XyyrCQjounTJvdVWEG2FJTfHquN2zr
2F0fr1apjDqtSN+nFlQ/trzquN86HgV9UDzKJcBdB6MdqFrPjha3HyS3Q1Mt/WQT
PrLGHuG8/dx4EaUm9Agy9HgLGgJzNbwbWCzq3MGVp8yTZmgRk4yqwzhhY6LKnXNY
4pOv0jmbTLDLMPUPm5Y2vAqdhm/AUfBQFx0rXraBW6uXbKss5nmtuYPVMmzbgVbm
CXNsWIZiZor6gEfzqyNCDUKqkW/kVILCYRNxyj784NUCAmAkrv7tcMaRhSoQG43t
QLkCDJk6QRjWjnJYWzmGHyRdg6Fr6n3xLWjaVWzUI11izFvTq8J75/XbjY2TZ7lW
XFijc765NaWbJWM78Hy/pW/p3fACAuKkTi6yy9HBXTURLUrEYnEFG2Uqj/I1bC1U
rhtdVQfZT9Nqe9EnjemMPFbgBOIqLzG4tvpRfiRcY4GoHxQGipdZwDXObwznbvNJ
RZNOebh91gvl424LtkL7mXy3e6MdRn2Q1aX1OfxNIwu57KttWPcL5OD/Sk58mtAv
5sj0f8d5o5dAqzwb+tCZh+LhlJxy7yYaShGZ7JaChvqiEbvgtDu0sPZlP0XrPE/A
2Y61v5m3b7eHCavF1MNABCHCg9JW1H6CqJRDCjUmnGvT4H/OU2ffXzlqCRCJQ8pn
gLt1zjBMOF9pStfGhSaJi3Cx4CSD91Y2IGvKuQrWHGkxgva7cZg7Dr50SKYGo075
TCPh0RdEyUN5dpUDdV/IsFEAGbKaxop5hNK7JgWKXh9q4uQtdHhOqzX9fxk4VHPE
oBE734PQi4Hl46FMVlnEwOdJ+6nMdhO2M8E1Y4eOlF8h2GhLov6GZmon/dqNNd4t
y7GB6nYstlkqjNZ8goINpeJVAg/j+x48nrQXEe5Uond8kkT8S34NQorc53g/cRWY
VwSPNuGqpCV8HaXu9LicNTcBbDRFXxPfiDPFGAmvAe79PzsYlgExtPhDO0cgimIU
RymHrGfyxNGov58TLS5fIjrAntzs5ITy9PLPJ/EwMQMVV9lX39draXXwqAGPA9mB
xcfMXi4MUHKKAwtzfSqCnLM4FARrzAsbB450AitUTEVqFmz6d7xMZVPRy7UnZpJO
ExnQXb8eZ2wOtGV6kRrVDpaCCAFizubjQgv7WShy+U78JtppQt7MpqHjmQD9UIvr
o7ppccUu1ty/r3JX58BIbGaWR9YK1f2/PPA3T+kiPSI5urvQSHU1W+XEsMe1fT8L
aJWNhJNcyxUx9ch6NAOG4ix1qhCxvIv3ZcjXrVF5V5F4Qg3g00Cxxe4tXG9JMQr3
QyVgmaBHULPckhmVVPWABk97ECbkcA3sNd5F9snxr1JCyQESfsNIzdQRpSvlcQxT
4cTl4339Tc3rysHAL42CIOr/6yxeWftOjta9ItkBW+sIqv4xgtMN1qWwJYOq+qKt
JQ9qoT4PsquoH4cMwv4+yxiD7QD452hvcSjCmBLFQ9f298vTsTuba2vERaifRa2Q
Si/ByoZ8bM8k5CPi375oJ25r5nYFwI+BgYt2clb8oSjcjyv8Bkd6LDL0Is3MkYJy
GBboGT8sUJrlAXN+glrjiA9cUCGaI2sWYRHJqLXaK74HGZoUjkBl/WGymVfYCpNl
bZpCGZXp0CHCBvyYAcFRObvX2CikzqDxCEx4EJegU4ZxKuIf04IsFYku/yqhv7R1
Cs2N9ghv7wv0eoyoacFkeignQfBJx3Flml1ZAMsjGppmtnghmVGYR4BPEK3Rl6Hs
YOGgVtZbkDK4Uqo4Ezt9eXZ5TZPGmMuMgL6gm5Kx+CAL8KPpl5bpJ9Jr68YqLj0b
ZJymAs2kZCe1r+pdRRUuyafjCNhMLolsXgRfhCHO/Fup+3pdIvyafVMwiH7qrFs2
x5BerYnOdSMtVwYgELwNmH4u7WsB4HAyFwWSubmdOXkmqHMK1YUqzSVpOzRd5a7J
rTyuGMxYbUSq1byBJSy5cqVKdHJsPVu7tlbGiqSYOWZ846rx3nD2GRMRUTlcg1Rj
5a2lfRNZ54uR3BhNyizIeHudw5MXA9V7Qrg6+A+8E3Xfi+MjOYzC5U9xnBRs3DUk
xy/VZqQWCObAgI1DsiVSHvhIWec18okQrJAabtkHopD1G/erFCr+itthtfBCe1KG
xpjtXw8w019YGUlMEAizT/U4uE0GfZwakEOi6I3B84IOHRTYovca+rLeJtE7zPYg
Fz7Xz3fpQ2UWNGHNUPgzBw==
`protect END_PROTECTED
