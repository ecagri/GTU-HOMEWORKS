`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p/2SHz0gYaR2/iXyOtjLvR3Jnh2MUtaabzY34vu5FXRHlcONQX4CC6awxRuRA8Xj
tMPvTi34NoCN6AeCxeJb43ooaHWGOSpdTE8LvDObxerogsVpQydgSUpGAeuAW8o2
yPRC8kD1N0sdJxzaEMobwnn9eiDYJlHmFansaRmUz0LGMprMcV92uzshfuczDYa2
zzJWwiRmQIkGmKDigbjtZXRH3o5lcCm4JyWL/tPeyZVIdNyXIke0SkO2M68vneir
Zls0Wj614VzcJJxja1+eOMbB8D4qvT0pWNvCdzLIpu/9kHDCuZf69hxGjwJO6W/h
mEVNGqbzk2xwNIve6oXW1qq+PjJtOQfEpA23fhhInb4++C1YLKScQEypMZKlV2TX
RPa7Hh9X+/kfAh/BQ2b4QCoSC++Qpf4TH3J9Nh9uUji8TgcW8Vfv3aFV6sVvABhh
YOeMEbYJ/rPE+u7Xw3vVIp+ZUFsRgS0s82dkema4S1SRl03mcNgJU4DraBDWdSAv
B+VDZuXOFEfphiwiDRN8myWULXQqf9YWNEPr1JvJRyx7UJR1mpwGYh8vmIrgHZt/
X1YPezl1rKUpRZp5EZhcxeoxO5m50JiMq18/x+VuU9C9SZI3COEhYRVs3ILmpcv6
7PGqXcQotcQE8Nif2Yjr+KFBdX9dQXNHfuNtxhf5fRjIAuv7YsU6x09phtYQ28F0
QcBcfneOTtOCdFu4st3m/pacK+T7kyUAeFuFfso1FhjbMR4kIHXfb5Pggte4RJw8
AlpQ/L/CIRUh239cuHiAZKG1q65HC7VJUskG+LEgbVh3cdtCR+JFXph5kG0zGXRC
CUbxxlithqeiCsS9vMJBIEnHYyt3Edu9EU5ei7qlx1dCNcX7yRKGwzCSSQZsC6Cz
13Aw3DVgrfsddJI58KLksRjmGPR1UoDUlU5tI7HwxpqIt6hAQwdf6DyiUSAhtpRc
BbvJVvrLwz5Wo6nyjQJ3zVisRuHEeJ20DsU8T54HAzD0bRApIOwFBwO+guL7D178
3HR3HVRkOh+ETxcu+siHeza9QJtHt/rFrQK5l5rYAjCkpA4wfX7En1SIynOgmcrg
F+4AkcI2UK11u5g6oAa31WbUOK6wQz+ll/AcsMKxcW+Oya7E0FQyqmGlCUAGbNfx
7PieKR/K4ltR5DNq9teDt3zqLgiQFAwrfrXGyCDb4dYw/rreO4qiVeSmPIwsNvEB
VcclIt9QohMdFgVYSnkwJyptGs61A8hh1Fvkqm+qBvzFryhFYICYCmeymu8cPkpP
3GmNBUlH9CIZS02V/CjFbA==
`protect END_PROTECTED
