`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tOXaYucjoJgRBItKBl2iEEivfbLJwbOIWr9OXwHExp+Kc1HHovAM+e43DXZjbCzW
tUpj83xVJaw2DbzS9MEVFO+v/4V21GA7HhciVEdke5ZkdagWBGj06cUx9z5bRWSa
LoKLj9WzZy9HwjP64/YZ+xkA0QRi+CqXA1UXCgxZgXhdaR9Hz85kFv+ln8IoJYQY
zPfKo+qQNX7fge0tbmwwqK6U4++tuAkSwlHssWzGdsbjwFc7zZEOiq6yxBDiBd4A
4oV4IQ2qSes/GqnSZj16KNc0v6ThngYPPkYUbLn1uLviYiZ0Um/3SkqrhrLLc7G+
GBreszgD/9g6xO3cw9Yr1HTYBQTRmLgjgAWsBqfkvFVgtlm2its5ilxHLsgbDs+m
Cyyk8lepm8DDMhdIxF9xeUKR9w2fRzzoiZ3B8eEzaLz+lyZhbY6LDTlcsgZeU2tS
IBlzqvXplVGxVvnHkgrtYTeSSHg6mkJhg6GdW8vKQ2Z9+hbm+XsIBCuH9lAdjXKW
zIn4L5X4DEepKY5AYMT/1xuKmXFJeFKp3Iq7yrRZ8pndKCCkHhtZen4OnH51zd+J
YHSBTTTUdojMBI0pnkVEPijIXI/CYreNQV66W8iSWI1ttjV/8K7HafBudIxkg/oj
GTq5PJHysY/o6Ar8IqTD6u0tBv3URpkGn0LMIksK0JoW8I3aUPzoclnjc54HWqiC
8KNj2SYaKMaChW40focuKtlL/Vo4Ag6PTlTDUzSwFJ2BfRL7I2UR4ZNaBu4twyEF
t+Ix7iyTWWJlGptApI4XPQXH58EcJZRkrIo7nCuKFgyGCW7R96B0WUQ5pUn+EYbi
jAgqc0/cjDC6XXJPcej0XXPgvmYi4LMh7tWhlSkQxJCuBOqXZsHeCL9xbJrz9YJw
33pNO/qxuOasQmTFMcPwtYSPfrRZRWjtBuUIkYVb/ZqzwBvsEByY40gMFJDO4/b0
bPEfUwXxWUvb22zoUrMNnWU5NuEI5tHLbU4RDvGvaTiUdqC/lNffHzu/gdGEXnB9
NTS1dFI4RKmbAX8DGWRTxZDE2mZxQ+bTMkEhLt2utgvuFGpuDoX57m+Wy1dOj7pj
mGxEV9ijCjAQUudnVftJf2meRFe7RTT7e9JbHBXN9R6Kpg3Kv3bI6hJhKNy8qoTr
ZJVf2NLRZ+KY9wqt9SxJUha7EDAs6mzH57f7dSrUSTgcEkxZv/czR6/talUTYLQ2
fDPiZfuGI080OKc2zMX9y3bBh2bDZ15D1d6Htn7kMZ0BIEmbNswrv44JMY7ickTs
TUmixSvQUuN+ckg5WjmCgx9NWf6nw6Z2sQ3S1cb0fIF8/C9nXEh9XyJvft3gp0L+
reSSLeiWKzeoX+Ailr/0fpgNU7nphGsnQJLVegECsLbobjXTjQUJpxuV+jFo9CU4
PECt5bFjvhiEVnaEOvgn1GYvpqD24aVQAE6ypjAHKMCeOSbefT2StwRzJn9EUkC4
OHgy+sq9jumVjbleQnad0+fRZBBr/hIuzGzoQrsck/Ko+tadZUJSYPjsqXyC+UCg
m6QaxdiniAY/65+EiHj3q0qSAoMqV1J7pkWhLGgA8oQu4pxc2kdV4jPIe+mnDwO2
IQwBzyPdvaG2MctXQ4MeFNftXPsnP7t9l05LX3tIleQIPkTCWlgZI4NAxbYEOLD4
8si5he4OuJlHi+tT22tIEDu+F6DN4OltWUw+PEkjZ+0gANp1hCf2x36d9hbFBQVW
gKQ0xyEPJ7ov9BkZPKKvckJi0npzr1oAtaeaZPA7eAonFnmvYS5KDJ+ie0LkImUB
XTvuB+QjyS1cyZI4B3AuIk6ip50GJied0v6JNCUySo+gXseSwQvEWlyFwDCO+wd7
EvMKPqTYKqPEPxEJL2EzbHBkyUQ1loZ2iA3AuaodqVwabxrMicL6oENJHqOJnWY8
fa9l0dq2hChubapoM6k0WzFVOGHd+VsuzEr981B5Am2fkKtkFBeDHuqVr2+8/ox/
1Mab1BAFbV6XbZTnGWJ4BQqga9Zz/SAv7IiTBUrwuCus/7qTwlO5yX70Pko+rtiH
FYg3KfHlzXEJYKPH+f0Pmn8Hlhm2UB1nH8Z2jwLe7Jamy8m3ZWnf8JthN/84AHM5
ewJsGdOSu229+zkqZC4V4+sUR4Z9j1D8iohSdjCZQxsRE7TrSkiu6GRnPkwBxdc3
m5WC3ad07CXLqcn5HwrmmRMmr9vU73tg9d2MZq7tviSipGLe/DWvkM/7j3aGx/Hh
Ze60DBZRK7RR+klmT4G6VhPqikwcAfKmsYzaLumhSfQNqGfloC6zPbLb0l0/PIhk
iZCOGcKKMr79X+5vSvuBS3F22p7fLNhnrnVuLDarDiNn2jxkCTBHQjL2/8CBMokY
kcwlX7rNiF7IjFsOq8kT/o/eIKh6jojKP3AX9v7AdiaM5HLOvyaHj0OAcylWpcbF
JzfcKTD1IUSjFgojunHw9SuausloFlT/An3t4ipVJnzQnKHRpaG0uVn+mLTWvhSB
FA/FxxIkmNTHKOnxrHXVwThyoUmnsoEwCtl09X0Cade1QbBHV45BAujKx19nBdAZ
I4D7xvxr9TKlgqKGnH7WovTBduyueQDY+jBqxhmuBK5IjQzWYJlDjF/RhLMHiOCH
5RBjKA0qef4ey+dpeK8fZA==
`protect END_PROTECTED
