`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YeCGfA1Zfi5zE03wdR7jJhDglXMhTRh4BXb9pOq5xk8lprxN01g6geIV/vp9Uzeq
Q3iWFRmgN/KOXWtrP3bvmkDuovV+pD3JR6Fz/d5FEKFre7hWqWxu3PWz4T0OZ6FW
xajPpatG0EZt/2lXFRcRPs+zxwGEDAo5Mb1shNdp9IDgNejiDgKpziYoB2PyHMho
P1okjUKlg9u+woRL1jGwL9CotX8CkkDW5+EBOTZh7pmE2dJIVc+5S+tfF0C9iQYs
ow8+XO+EsFbND7JN6ugrRYr35VcvSMAUiOJPpgQASzLzjNqddVtxjwMMncVFGJfs
ou8wVWc6ExyjttDdS8Z4m8WvAjiDsYqKMxmJI7dlggMjSENl5HVroyqO54crvLWv
JTxjZvmiG3pFa4pyIw/Wc41lUeoMo1YAG/l2KKcd1/qn/ruYlOTfaa4HwSkBFs0X
IbGwlOe0ogbdg4jC12ZxZy5rVA8IofNjb0y30fgcrS4b0wHcmj3yMRuzkLsSh8g/
0FNnBrG5+iVtoQuHSoQ7ZWChkawmjkngVzP0QM3ngRWSaLfsGzppwNWrxBVGjbNN
KJ1u28hQG5lZDncIZK8xF2R87kQl1+jhFR3JZguJ4BgRONVI5nriTtJr12Y80IXi
FuXbqRRRnXX3WBTqERW+P+PeX6l1B2MxLScduFQvduX9oB/d3JLKDt5oKWK6+QF3
oQKodUMwA383KM42sS+EGi8vldaByBw1zQVUl1wUz9QrxZd/JCxU6e1Mu+YwxzZY
Tf056Gxnrrm+sHVTdkIGENAj6rtQjlbErztPoL6Wgu9wgQD54S0kzbUSHb5cDr9r
I5qfwugLQsmLdDQxr9mWpjeR9Y2q5a0mVs9La9+QW4bXuZVjQWUX+t2XLn4k2Zx2
5pNg7KhqkD1+szJIJsph2L1NOPPe62miBO7bKBPSrGGMQA/1YFy2waZZ5PzTJBDu
cmNb1B/7OmeHrq32hYJgKVszOccS44anK/ECXPfZgzVOX2Ng5EwqsMn5K4anOpqn
06f5mmQ1iiksfcHiKEkPGpku+egMsNwDXXUfUeLSuO6OsfOMu2DfZpSDEOQJbCXN
Ln8ulnBSS2Fd1NEWTihEPcaV5XGWjjg/dOl4quO7ZAQdpbqawiyWTFmgQgNPWo5i
qaWZy1yTRcOGW49cNj/RA41Qq8yTlkB6o8OxZieHtn9whXQqM88bZ8pamabeC58A
7Ckkr9WtU5cnymxRckFIIzFfPXOImksAEm/7gDyixhtPENmZ+zz17S1d5q29Pcyx
BgwpKOXANAOHghB+VoPNkbntGEiBMBLGi48b//qUPTfpKQJ+WcjfGDiv6U/t/61R
xEg6O8xKb7bNcgSmfDkqwi4ubRyA/WOoAKfknuLxpTd7RSm6wfb5noKZadDmgjXC
rwUvsYcql7qLEEPkLp1vQpzw7jJiOhkeHs8vhUz7MhNnNOouqZ5x/gHAwmImaUAZ
T/4Uesoz934I2Ojs68APkUHl6YZZPjU+KKEeqVMMiNbpoDT3l3HiLUsJrxpCcmo6
zQEqywlcL5hngPTayOEj0S9J9RVKbaMJOosG4Gs6zQ+W5nzGXN85gVyex+gz4PiP
1p4bHRlXlnD/3dWwCce3cpT8gaOjUJlYyPuYd6C30fjWhItEvahrs4CZbWM1E6Sc
9BqHvaAbheTvHlr1yl85/dnFtWpu3XfuEvfUqVJaz4A4Yf7LUA6ii524NaBvysNL
IPbY03FAQyWdEBKtPt301EIFRY0kEpco2VeUNlAXi+dElezavJZ5ZdYmnZKlT8eX
1grKC/MKzMtl8+DPUP1ET0qJnj+fvLXk6rILysjV0UgfTKnCXcnHBLqjAsngX8YO
iEF7NTT+OUWtMUrpcxGqXh7zFf/vQ2s3rRokd+p5VS/IlUavbAsATF23n+M5EFgU
vtaFK39hDx7fLHpFviNinLiaV1Y156KS3ZmuGvo9TrFGxGCYhJlGqC5DPQbnbKrl
SlKQYM8aZ+bA9hbTMt1HBxOJ3ZzMnc4Koqj9BoNr9nGplBjKR3khzZp9yMZ3Ifgm
h9SDRz5hpXGzoB+NB40pgfs4B+ueLfpApx1yaabY+imoQdJmKTX/M4iT5t/VkLv2
CXOaCQw2cY80Yg1TsHI58sPGehpImZDnisZw8ITbbo7He4vkpqGrvMZ2+YU0ifye
N9qM3cJUGp7CU4BhpSklnWwSTmwVqgbvK/GLlvIxelXjSvcmgZodrDQxlGh9xa/T
BdWlvdLWvEQH4BTkdu79RMcjTXRgl9Q8PQ1U2FIdDxitwQaxyiHGvHHmaTsP+Yia
e08I8ltw5wovKlUEmKzFOtpjyAxZsyp4AjBmatlOkEmgxiJRR/CCRxkgJeFCCImd
BP88Do9WV1gtrCDSxpG+W7nIb1QGcEY+DrU7bhKA8IJ16G9lbfKyJlZ+/w346W0k
0JCYQKcLGRPx82Vovd1HZEnWfnkc84qoP7zlprYy+/Kj+oMEtCd3t1M3HGB2RACA
houVxIPAFHFE2cbNPMZqJo2ZtugdWqTBH0S/h/wI9rqy4eVHVQXckZNnWAU4JpKx
0WFZZm/5gLCDDdMtksLJuzHvBGTj0RM3r//c6MOe7/EXhAzIrPiGBABQhZXF2z2L
tIi6OiH1G9OGhsGtv/ZTT+0qfb4jOZV3qucZofDf5rvUuZav0PI6etspA3+6Y436
dbtOFlSl0C+2gepmxwTX8+2pa7ffT+Y0YNSW82ZznBdSbbCEQfZHBxg6PaRaLzNT
aBuOv5PCwpDgySu9soM6+pJBWEyE5wB3lrIKYDkhoc8atkxKxVYOJcuAVcU6MGnx
04PLCGUB951P+8T6+y+xQJUIDvfz7hOR3iV3ZZfzjOdP7h+dacRZvMmi5+k4UmkT
+XqoTQVLyqdLwesM4maxAGv21z4waXAecETrs8+Ah8WBtnVMRlyQP+SDihW9O2l7
Gen77NIycC3OQ0yrk9skCIn43zz2T40aLiKVoQlG0hddJBGBA9bBed9ycTWktYMU
H31jZNzqhTgJcDhs/ksBiWs5x4GsNKO9sNx8hAbEhfw/xakwD+Td9XSfd+TlAeWe
t8OKGOYdr1VjFa1Xo9pzemuHGE8cLu6oSEAVcRaAUDRYE1WT3aBJWMAQs4Xosu0h
Ic+jdql2jnu6KBE8q3ZQVAbS2+U0G++qAHjWewTDKWU4xj0uwaIMhQqwgF/KfHxG
OtTWf4jcduMWIY0cJbMf3O6q6BO1K1nbL48Dd5JTKqx+8TvZCc53+uOnHKi6NQjZ
0EBu96Z++ywYi0MpsuNfYiq2jIcwm38ewi25kF1kFxIDu5a/YZGDa22+hKmfvdLb
P9zIaH/CImgt+xQGE1QKx8HI3CH5wDV0eANy2RNGV5iJ6BsvaqTLP1k4cVdNBzkd
skNbe2s4zTo1w0GmqClguJ6F2/NkXLgV987AoX0SY0RMkBVR2k/pVIpP6Vj+qJMg
Ex1WNEIOQvznzsOH/YxNrw/fmWN4+8N9M/r8x6sDemslVnHq8d2mJTICyPZzwFGT
V2Ey2J2tqNwnqTZyCgIp8LrODvNNgOhU+CtO7gkEzK0knJkk+i6Qau3+l69EI6KZ
JVyyLlOmi4n+b5Gh9lg4NZrG9EHQMVFtQbKr2AgfAHqm+ZSwi0MBUxw/gP271Lrm
m9YnK/Xtxc21XVwXXHccBz7oBXcpX5Cg2KNgzDR2+6oZG5LbbRMGgilrZWrcThlb
cbVG3VG8un9MTkevcBIU04CCfGnoX5/WGrJQYYxgNB0vNJxkYYAZk3RnDO7gx3NL
+Co0hH/bcincLjJ9KVLEbybIkLTkwFxIf+YvtKtMmNQVs9R+/kOf0eNtAg5AfD00
aLt4wnhv8YEI6VOQMK5SV99GLm3McBh0eg9Tyv0XM+Yq+peQ0sgLgkXsjPr/rie9
lfIw30n+QczlP1/tyO8dkz+t+aK8XFxd+nx8I0+8183XWnWOB7BLP4ATvznCHuT8
1N62iKvZ0KSbVpNhfT6xl6OW/QcYpS46XOIdUoL/aKhn5IgY7vCe255dfEO4s7uw
DcVDpxOGWf1mx2LTqo5ZYG2YA/Ka/MjnaLPAV70yc92+SfAXcedAfoHQBnz+Hj3f
wG0/dwYuO9MPdceVjTqLMB6OuTFQ0KFfPugsxnrTohwulIDhj82Pl9UfQ+GiaUht
0E44/5hxp2Ev7z5f6Vc8OlSWD6ClVjzHXYBA2UjkWgKM76NLmfsD3jFa+Sei+djj
v0oOGPG+Kb5vYnc+sCC1p0ri78Mcf5A/UfAamM6+0r/cwhVt5pr0v/1lPjKDsAmQ
MzUdAbOITlNXd6wHwok/+/+CvNuk+uRNhD+WG+ZKSX53j4dr6rBIEtgrbAaQEa5U
o3UBSn49AQ9Gd+CNKQnnYQjVbSMiFMUWbatwrn7xFmf3+y8Sis4405+lA5r6t+Ta
OBibuAdneOstGoBEU4zNdTHGklPo3t8yu1hGmYmXeNQLgILzK1slx2o2AhmCs6Ua
F2DXbSB+RK1HuvPVgg1bBqMb4Ul6SU547qU4gf1bjc3stJa77M0B+Ul+8NYaBRPd
Inu/9xQmC/7PSTAg6ldmuBfbegimQ7vkGy4QykdVrr3qsxhvYqfMe+G9UCETmqzn
e1mHwPqCSrM0DOvXKjYfhEWWlEQ56a81Gs95kVtUpt6CxCMLhsp7vLyNIpXpTFIA
pdu8OZBXl3qgFbWcn6NEe5dvqgu1LbsKX2TSx1ya3TV6O94qrLPbf6q+nHejSY7b
l2Qg/3fK9jRFiwsI+6Nmhi+AfD7IpA7QuClQiEuhHPUD21vsJm5k9+7QHHrYAH2l
zTM6NSL0VOk1G2roKm7FS4CDD0XN2dk+ttNS2VdF9xIhjGq8pDvQckl0xOOyYaRS
7hk+YFp7sDIOFSbLEzKYMk6NdtCO1nId605JdL9vxKz+Q68i9PAziIxYTIudSfRw
QGBdDioKv4OxTUN+zZ2/8EGaXQ8Q8Gw6XJeTSKDZRBLNWWlLa2jWmPwwW0jBRE73
FZS8FA4zxdQI6QtnlsAPIWlBpvn4u05ogk8rdy7rI5shqy/Cqr2U3Wliz2bvyLqZ
IRzEX6ffEHHnx0cuw4+E7+lUwevyabhuq1wsp9Q6rYEC/tFrd2Scg1r/JOFDIyAx
MQ84ghkBtby8g5xA4/UcfV5IBSl9YiOcNLRbaU+venkG9168Su+yn8qTb3ejCclg
Cr8qkeDUCiOSxXVeXVAlgt92oAKhy/jTpueUH23qiZU/75XbClmaFvRP/n/lIoXp
PmWtzQrLjsWcwx5HlQqV006E3l33kYxqYIVXX2FXERJtaWzpZ7zyQogQV9qsC9si
Bm7yvNTpP7TY0mitEJqU9fkzV6qlcXUvhZSmusYmB6Yhe2whZPRN/9XN1ceWWTG+
L4b7Qt8oiCnX68c63JIHRR56acymBw1b5xGxXYugrPcghS8DZNneM1+ybqRALAOA
6kdjiL8Et+jdJqVMS5hiBtHl8toBK8niL/Zlj+rCNfPjGqQ2JKcOeSvEcPY23ApG
EOeg2j8ekO5tcSTiX+omego3gYa+b5SGJxoiSdkkAxfvXQDOb1qhoQFClF2IKJOt
tbj8xtfZwQmxrwHulgIz2821tdEBS01haSyZtbdCrW6i/novK0WljyaC5HG27yK9
cTDY3N/Qy1JPcnGAenDKN4GlOr2FehSIAqcZkD0bJsqhlphur0cajwIZ9swgBBf0
WNarOKxP+2LBOSXPIBnJgxVlMihWlKaEEF5EgXg/CcveGWHxGfFiVmSKu8D9TdvP
K8paUbu00H3zdoOAjRyapZq0ClSwo1T8QPfKXhh/3zKkREnXFFzTT4yZSmRHY2c8
ed3ZGkHNUmET2vhFi4ObQ4Ldptno4hDOIcHhYaaivDMPEwsaQyh2LUiFpyUhVUTL
9xvpbLhpqgMfG6skCQQm8KIrduDGgp12oY4sfp5CDHdepyDjZhdjoi89ZdvUuUIa
W+RzdkklreO4sxixgOLfqFhsV1ENSbAiuBJg7dnMh+t1T9NuoVKAMjDYTIY8BACb
qWui3xaa8rALise9TM/0gMm7Ra6b9+IiXE2aa2TveqshdttKqXJluDzlXyr/7a++
WqCNxfNuxtgVu1KpwDmIeXxRyLh6i9sMZp3a+stSu0lCKkOVZVkk4g7DCpfGkXyT
rhmS/ZLm66uPEHLi/Dz4IdMxoNm7ARkukMQVACE7I1FYRvFW2keRgf2HxnjGGPGl
jnt5Ig2XvPy1SaImuZPixM8Yjq5dZbcLoojE9PpvqgC5EBonz2/RAfAyE63sh1N/
ZYwzMko4e8yoMNNO09C/kAjxrqmzxVxvVf3fl5eXlF3Hc8evSi5ZStux7Vl/11ba
OVyUABQnL1d/yssP/MEsdcExDbjkxugaWzi7fI06RDjvYo1d7ROvW7V/OJBbVxfC
t5SquzceKii5Vk04q9aW2NucCT1MrLvAZ6QNtnKEQpi/BkwDAfZdUl5nHFjlrJWg
hh44s1hD84TjYVRaXFYbuaKd/4LbsMycb2FHxwO+YPl5f0Woevc30CsBoQtUSzxY
8k9TcmrlEEJQ5qquz9lP7HhPIewQTb+mT+nItgXjpBQbT3dxQhg66vXi7sl1285c
OWX1ONvxFIEj/b6PgXruwjMU5p78EoORvnmhWKkRAtnCieRxBRV9ZS+s6Gm27qa+
+a5I00G90kUq/+H31cPtoqFzlIWxRXe6bBz7japJyrV1AlbtL/1L3iqu7c0IR5Yt
ADoKJtzC7oRMeaW3PW3n+hzx0dVMKLIxPImxim44EmI5bPPMsLxV+d8JgXIebro/
iYDz7pBCTSo6v8BHo/yepE+1MmMNRg4LdIv2Fr4Pm0MzIMVL9Cg9ft2YHtzA7T1c
TvxzSCuqaFFAs5p2Du5tDnk/m+AWAp4FU4gliJqOE3TY4HKCtSluoSxdhrbOpcR/
hxrLQR5nmk/H8p8rLwN4g115GpMqfob/zkj3Ha2p30/vJp5t9vZTjcXbSuVfDjV1
5HORUWOGSuYVxswxP6SEPEWN+W1GTNGRrLG7MdqGkFjyj1RwKU8NPI+p2gNeyJhm
JioZ7LBYPXZpo/n3P1NVBt6etu3co0hsndzpdfP3QRxvHktM4EQaSu5SWwf+vGzS
CmnVM5F8unNm8AR5r6LmLrcRiNPF0gl6l6l73wUp2f03RL1Q6Y5DcEuvZsEfFvNG
NBSae8ObFPqhSvJ8SisqoU3NZVNuVP9CYnhTqsAPhxxRPVPTs3HUgvovikoWaVNo
JMUHFQt6o0pZKwyJ0JcmrF4mysGLlmDBDys8d754a3q6uQwlNLyDMUUa0dOWt09C
SNFd6dArPsLOaixQc2GtMlNcxpYVxRNRugyTFtBN1y83wV4XI+upUdI0Nkp9bMKY
V9th0NOSSG0BWJ9jjZFYNmVQGkWQxqG2Ddsdf7mZ1k0oOgb8cp27vLUBHK8Tyszk
5k78baM4RGruzmHs9iEBAFzZBjFkxuXDBzzitCU+T0/gtuLU7KcFn7UXsaSsBLvY
Qnd+V57m+DitRaLLqwI2R5ItO3TJgw18d5Rk01HeDJJIH7AC4tM88wPmj3fiTIXZ
WrdUIw4kWlnVnAMXp5Bw7fITumgjZIdisXfYOFA8CtmJOF3920bTX8jUNCdaajMg
xTe5nBjj88z+A6/uy7bNcwY4dwFLUbxDxWMCNsyZmiugcT5c/KAkwqbuNKYXTUiN
0QyF8J0vv8Cggp0R+qh92k5p/YNh+aYwOiuaAmp4ePCParXm/6Op3sy3MtmlP1pT
a5BzL7QjbQGE6mWyBnwR1puzBKW9EGfW82Rv+ZfhiZP1XaJtnrCihdQB2BO6T0P3
dR+PKyzpWZKAlhKdacnq0OofZ7JVbQxAHnNvW0B49vjWuFsaVc0beeV3BaC9kiEe
paEb51pEYWT29GNAHU266YJGGnm7WoGT6G2uBhmu0VfZFzNvFP2/0QJF2lV6L0Ly
v1MPEmpZlAe6x79LGV9FXaorA9zDNpY0TUwNs1TjBUZTBHj2jb1SQkDuKuuBFKRD
Q8Wcu1DLRILjsCWlaHBgAd3SqbZSYNQnfD5Azb3TMmm8ZrDWaPKm0FTMObdVMbpe
C38ltANlM2+3TLUJjREKxUkMWx/S0+y6ycw/kEBuulf1J5Si+AFW/q/1neLepmce
awHwjli5oFt2s7J9yH6fAwtDcfLm4F17AkBIMlxVsmWTmUs7wlXNMTSbGPbzE9ac
e9yKsGRpeVQxw77vhJKjwyrGiD4uamSz+J1wY9ACdIPYAxF1Ber3Ge/M3H3u+87z
pFUDdPnOzCfGHJPmLp3zt9WBq1I8y32BQRx1VaN0jjHCAtkECkK6xoJl7ChWhRdA
YJGizHcBsw0IGvGBkIT6ur+rFUTblyDvM/ElXvq4rsV8hqDwhjzdIYvGcILAfWIt
1meW61G3cmo2DapDbUqX4fYHZuGr/APg4SJmbsnDeHM8QkyWS67MC/mEa2URau7T
LHbOU+TySrwpsJYPK9dBWS2XiKnnLDO7af/eZ7ogAkgLvk1eLBfuB/1nHaGMrsvn
hfqrOa4Fr30wlyf41LKS5F+y0ML6Dm3G/HyOLFXX/I7UHiiRazzKCKAA5ukFpO/q
2P6o8YG92lal7xCPujO1eEIP2wQugNmTajpir5ldlJvQBoCngUF3Kdd0cgazkzsT
a6S7ZmcS4BK/+SvKaKUtgKTamR9ClebACgnoW/g2XNyy+EwYU9+Nuu9TVGNrEGFL
s7k2fiUicHQqG2SP/rvtnTwiPmbmO/Tz25EkQPj5m8n3dlY4LbJubxtrW+72szWv
FUFG3ldW2jFP4xz8TzoBudx9FbMDdYLCJ0ZKwBZ4QWFXhJzFwXX1onAKddDmf9+0
mdJakaeMvfxjDuPPT/5DPXx1BQv+k/dVMI6eVyqVrtIhvUR68ToDhjwzlcM+i91B
2pXn4oitN26i23wYD7bcRyvahTkHxhfJMKBMBq6DdRZiUDnU4hHEM06H9yPYAdQz
lMJe6+lt3yJazYvROxAL3+xMDkGZehBCH4VTsbG2VbTJZWY0HWNB5t24J0tJIKi7
za2IJr1v3GqEifetANC752EGKBvppIUEYFS3de8Kt8YTZWmn54Tkl5J9frIyC8ZF
bW0Zl5/kc6W1S2DvWPegF6WlZvbDASpYulIKsG9NLpoU3qBqCxD1DguLDTqzp6wR
8x+k174j+N+aIYhjifyzxTlpipmfcEp/7tZ4kZG5iNTgLP1Qoiz+sH34v3FG1EqZ
aGMvoMI9ikKBYFqbrYKkYTG+peaGjCe4BaXe51jUjRIsIXtGMUtqWrD6AaOvMakH
4TXh5TuUDUbfjvlfzOafS/DTUxfsdpJz4+b1YKQRVucCQTxKhU7FdZHDjowRTe9y
swg2bj2o/2OaD2Xpo1vDObXNQacJVOtaztHdaTZbj7yOL9zFt2gOJ1G8p7AnN5Or
5eyJ4OW9t1h11YGpN5qjx4SfoI46R5xVO+6vp/CyC2lIHYLvxXdh24xv5LoyrhLh
/HYPitZptBB5lTOVX68Mnqs7iLzjdtkrCsNttNL1YLG3MIjJSPf078Fkmfh0w2pe
iaih/J5lmxpI5ENT8Ab54/z2DSSPdWJaFnFsft6PiO6/zmxMMv1/+UUeMDiYLzYu
kFRHZhIZlMraFb+z1Zi88KInNlzRbFZsUwSOAmBX2Wf9TBI/rsMuCvLXTkxa7iu4
9kgUDplqX2spxquxzjAIesoX8bA6v7cvcxyqAacq/6jcG47FXmpoedOauvMgxONH
zI5pZFfdV2hmO/JDuwnYtkn5EClTNqzQeW/Y9vjfOHa6RitTm16RjWbNR03gf/6Q
K267mRrS3ob4BAK+ZUjxZIF3x0A/Ec57E0/McHJt/6QPfWedjUAGipTYP5ZgZD6f
SxdzTT/ZO0ylHqBIybsLCVmmF1znkZcZA4zNZ6meuYLeXMmrRT1TuZBt8rdGlEpp
KEGBKY+ePagMrt7xua+933ZaxZyLsDaSfMsLNSMJRensqJcee8Bt9RKwUTZ38a1E
lL1DPWAU/LAHiD8OvmdeosO4BV6wIG9HbcS8L9xL+AqRbOu1v9HgQVOc+jx307xP
1eLxr36FcuHL7uYKlEE1tg3bZEq21kfKP+uZXH8Te6FngrN9IZ9BjnptJ4aDO8xE
kMsOC8FlEliaGleTJZWZeLL1CzHl7y2ZmCT+mTsA++fyZVW6otpL0I2lL2QdQMCV
2Sp8KRx1eO1xXXmQOhzWNxfinkJJrbelJyz4yLJUuvFtNhDrUOYhu6C7gYSzIc5A
E29yzbTMt0b+Hn6w+Id6q8UReJZNupHB0b3/7nY5ysUeXuvRYrONsxg5hSJIZ9sp
1+PqJgy2UQilrdjUxOw0DI7M6ZbfW8Rxa44oU9l0mFML5x/sZQmngjAC/rBrieD6
1VaoPVcPu6JlaLj9v6AQbsOVLG5WJAr41GLqQHxHR8XTeoM1G/sEjFW+E0u9UKvM
12Nx/AJdgyGH8pCn52Zc1W78tUUx6Rcqzdz2OZTOqNtJ+tMCUCg0Pxw4Kqz3Y1Th
HSEW7GC31szWf2V0WDcCn7iWxLvoo2tq59UK86NUQjngsl4Lb8oPIa4iBnwY1qwH
bnwrLkimYwCKD9ipmJfCDVhvGelr6iy+QYWzIPU1wL5ZFf/mNyOi8i89hdfMmlp8
6U/xlzje7U21wPmfW+WM7FiaUBThN3/dQo7MsllggR0ufh6S++h76YPJu6IDe33K
7MqEBjiphQlkfa20Lb/8Vmuob52i+stxcPaeqopXoyroY8e/y0hqzBuJuxayn391
djiOp9zuEmEei0HMfDWx6wfjq4GJjXJpBCRSNaxhKo5JemQH8pqaV/BHhplqBqUl
pIajCYDrbg/74YPdKtiNjn16wV6qUXoCBqFRlIyaFVi7cLEOXOT4d5+KgRqIuJ3E
DYd9/y86kyma6aJX71WJB4pX6tSK9uGMV4DEJ4Ycf+jrpJdmfepn99706Ecyncvl
17wlfIye+NCp3SLSHuSYIIk+GtAnpc5sbYnHV3cPNxEcTaPtTH0NODzfkaCVHnk2
EsWqeYKLHIBS6V2ZQqoqMkY2dpLCxQxCerWURWS0EIJMVQ1wKakCn9pAnV9rn8Df
VXp1NhW+0VFGNd1eWF+nMt2R0Kofpb+a50s3qhR9wfasiPnDsAXllIAznLYJAAfc
1wOvwe/GOh+MgNEEDSCIIO46zsblUfbGyfn7e68053RJP/48dmiWQYHmPu6qvtlE
LHYGF7GYYpkZvt1oxd7sFSc1BZtoZSLlCAALDQ4AnxuXXA0CdxV+5HA/LlOpLnvb
9GWFWQy6aK7zF2b2wgSSofSaN1COukvtIBYWTcvEH0SSTb4Nbd7HzLMsRVjr9LT/
CG79A2HoXxHdkd7JWPgw7N9QwmqvfrS9t7u0MYDByS6wexeZHktPFtfCZRaelBSn
Lu30QHRlBr4PWMa0d86BAT/ppDLWfKRAEwgdcZsEnJ+ZVz5/wzR8LfWnw/L/FRHf
uHR20ks/cpJioDejdzde2HelLLhEGWAEmlcoDKRqnYB1rgItH0/ulOC1BO3ElPhZ
R2G07IQFbM92cx8QvILBj5BmcsREWSrYHbpse33ssrKjIgEYEXJ1fek0wdW7E0+b
99qSct4L2f+PGUrnTs+M2AcZUERwdrAvlCwGK4T5aUVZCyWN8olr6HKjfAqiIdjB
Zp4sAjlj3Bf97YqlsIQI3kGl7sFCCsBZWPm6UyUs4TEK1nVzvDvBLd+ObeXjKzcB
rGhaAh0GpOfYelNHNsKSk6r/RbrXVeyVnypzyDxAyuukYPy0mUqeP2hPfdKf4piJ
w755qdE++rt1U342ENLT+Hsu8+D+ysMslFaSFFdYt4Tv7SkBXO5IojWihFq9GAxy
jYGyb65TWZ5Jjsio87cpaAYN8wjjOFnmB6cbYKErNPB27T1rz12+lExJJrG8x2VB
nB+sBZ41jnbtI4tONp6TdNwBkjCbIHd2ruBtvj1HwGB5FSUCeq1mabM7ABwxp0Sg
QMX+0LxarSUh8HVeTDo0A25tL55wR0cW8+DgHoDvM12DgLiaZMw/UA2PR0DVCBuZ
vstKwip5wNv4t5ximBEDn//1H5DnuOP7tXmkFnI0+e5wH81noeehcl6wxv0DNZJr
5sL6HRxE0lp9apxc69XOmWN038/G/kDfWQB538ky+PgS28N/gqndFilbz72w+BFr
lsWvF8uZn7ff7QmsTtNF1HqG0+pexJoIDpoFZgjFci9gi+zTAHJiuja608fRxWJL
43uoy19i1ZX13FP3zab5dQKdK6ZmYP58vVNn8ezcXkA9PAjdcegn1KRFnFyYPORA
L/ijpRo1vQeVeiqYMjfYVtKqAzsTu6ovziPWGWRCWwlkJoMv6EAH/06ebPTupcRH
zKskxLO1R4ljJrojMT/qGoTB8Ni/Edd5uUuAGvT2JwimJBnDy/n3MEuEew1WdHNm
PryOtD7a9eQJORwU0wCEy429nnQzOwtAuaU4tkoJPZVzoivwVBLqbfwfFBkBGBbg
pTFfV0UoAPHSoMSuMcnvYLYsl4aoiau2o3T2y6vWUJQKqUzrcctaO0/PXnStlVKh
td+xxykGE5QjXZceLAt/MPO5jQPC2ncW7hI+MWpyKWImuMkt9xPqr3SwHdnsOJzx
Wy/I/tHZRWM8aOfM6nd6pIj4gp7rRWYrGzQua/mjqkirNT4SgW/zbRb/yrMlaKB3
NFlrj8V09UnEr+y1XL8+hDEvxVnqlT+4ajPtKTgNHiihFJW8qCKfgk4FRGYz3H/H
9vqjte9WI9iEZzd298joWN5SHRK8VyZkD/Hm9QHq0DOF0/oiAIChQ2H2mu5LQSHE
4mbot/26fJQW79a+p4nuIQUKgBpzBNL1fQ0ZSE/3muutJPahjKGUyaojKOQ/HuMv
s0jYhD1Bo6brb8wxxPHiKFgfSA3dea6wImWn4KOkbRgEKYGqSUjil/L4HKNouJdz
jgQac7+Mj3BN8JGYZFLjsmUSGP1ZxW4Lds7h45faNlQDJrLNbEdE6L026O7qvs4Z
7s0nhzQXLy0VoBQexKjvxjk2zBPmPeR5pwp0+7/ipT3WTc7nUYLgqre6ryOVyXc5
yHDamZXcNW3bOrBkUxYxk5/S+P5Wmpja7meVvOeyod5Dub7GSEzkm43fCYp96/Zr
3d1YCAWEz+Ox5jyRcy+gL9LSjDd5k4g9DYjq3AUl3C1JRhy6rQvsSymqc8wik8F9
uQAh4ET7yYKFNznafXvvzZmcF90EbVUuQWom3NNh/ysbqBLCaXuIem74uktlbiiZ
1j8jYuM1tdvD787Lp1XyQb2Orb7ah6OJrpqIX3qE6+fIckHFvq7KbL/shlqNTgN2
WabX98vGdPu2iUuFwO3y4ECRVTrhe+g/5lw3JdhfQyi4Zh/vtWtg0NQjABwJvZLA
tFFQmAfYTZCV7kreJU5fbMefea7L4i+dB5RkL4Ts6dafqVUy3fVYajdNPtYvoad+
YzAzNbh4kzbeMVqmsduBZdcxzj95dNPzdxN2d/5Me7DnOmKfYFFqVNCIL+ioGfWG
r10GTyuozkGShGgALjXa3XZLk4oANv1RbwjSqunuJSPh0nJBqVfYtSoAt7p8st9V
fFkkuestENIwmFnndvY3WCW/Ed2drW+PAQj9cYLGLw5URBP6sBa50nTVAqpMfO8P
i7+bCmiH6OSWOqvQ95jP4zGtZDxm2RH/hV9J+abr8gnbZ5KYKe4MfYCknEu86cgV
C12RW3wZsOqlwyDXseFM8rd4cHXryk6/yEv2nTHAA76CvRDdXs49Yp/R98y0CguT
5gbGQ7eYOjcOzYpkQUFK2ucq05JAEIdV4F9DD/y5nq2Hu1jSi96PwChybqLusWph
gDm4CguGf72hhymsbt75pD2RzkPzZiFaM2M8cubSAQ/znEC5048W3Sg54P32opzB
u8r+wL+g7D127dxcK6GNJXEYUai0zL2SzPOXRD48YmZV7IbNQ6t6iFBfylABYQof
Mrjm3pVkwWdQaBjf8k6uq8Bird686pUxtTvaFaoC82mnij95zn9X6ugInTHvpTy+
qBfLRzYOIyb4xprY/t7fiJgnD16C/tiHP7Pzc4AH7UeVB4BIvA/P3vRu9EhwNYEw
Vz1psAg98+DWjE+Pdy0nrlMnrDrnVfG2efXKlF845P6oc44I94p93hg3x8Tp/EJV
3PdHNPA8+xkZnuvVoaKxZQmI7Lqydy2YefF6HeWN5I9SH2CBC95yoIzJsFua73RX
mvzBwbIgBxwtypUMmoaJxoE7iDutX8QtE8hbf/G/Vtmj6/xgEk8wOcSERd7uwFq5
5Xm7RKVtRjlCxxGNHYgSdeJdip+s+Q5TaWeSM5dj0t/6uLDvfZFdIAkQ+s5vOG+S
9Jin5bH9cbt+Ef+MG5hdWK4ezQzmPdy76UHjyuNTaypSp+OTB1phJvNu+YokR5v6
YTVw2yS54sPE+RD1Q0lUIEyvAL+3KWLL95JxJPAGEaB4j75n+mPe3BazD+Fml8Z0
08gqHGFMn94FwCCkq70ehplZzQdOzNI2VP+b7N3xol6FLgBRBDAhgQsZlUbQR+bD
H0ImIoUbkfcKu1udH67yUKDLcCxULqY4J5X4nLPyGfMgyPbi1A6xZLaE5gPkgCOU
5YR0Veh6ieisyivxHrM/QOzmNqMGdZmwc5k9+G7lUYwdIcPEiuUvvUnjyws/Lkmz
cT87aXSbvOVCOK9IIhrCsE3EsytFoW9zGIsQqSqj4Jm8hKcx+uCZc420iuwL7EIo
pEJnJpekxz45+VAF5b0TzUe/wTu0x+Da5oi2YUKLEw50NLDT19uTHPZuMgXF1R8Y
yfGMXi5X9xJThM/S5dWADlsLmL6ECsMqlflIkEuvRin5wq1Hmj2kjOMYgeDv63l4
vl9AwuQ4m1zKz+zFtPIvNocp3NaN5HjqMRuyRxAln86UTC/wwRs9SCgZwy23ioOL
3Ebc/A+LZNFocfcjmwiqiqeAQkZxZuOIKfJyGVn2j21pdC4YAmp4yKnCodcJtJdK
GDomI2WKhaWcGNYkBes23o3MtJpbWI6AJx+VGWQJay8YbihsejgCEHjzWtOKqJAa
0h7Cb+MKHVzNSRLmO3kW5l+cK2cnfUjiolAxWunsfW6Cje/6o0tIwOC4XLm0r/9B
ZzTaDNSol/90FaFqU68e3WAs8Dj7SsUMNk38EX2FtDVkFTyXN4sm4PsYQOGKLr2u
Q5cUDrB8HByNW4IQSfq4iGYtgqHxKuMvyv2KBdFwIBXtVu8zqwQZAbuJfJ22TYHJ
FxLFnCrvTt5Do2l32J5HMVC113uZxKWyhL49WLI+bTx50KMq4MbX+MSrZWeiKAA1
5jLGC/By/TEaKWFBhUu96olHlRqLrJIyw61tBis8T6xhDNbJvQEB6kXjtOBTCG2b
IPW6VCBX4xOiO5KlXrzvWu9SBPTJivIUX00pRaqx/yxWTFOtGzhzymjZQwpQlEeT
1DGFIxYn8xE363uzowDC2aj4EIS80FWog1fI3dzZpVPtfyeZOcSkrVuIMuVkRqb0
wlMQ9Z2TYgZO30Q3fYV2IrK/n2GC7O148N0clK2DWffWXrGVpJtxWNSVu0QapPY+
vFMh9/E6HScWrdNJj1vIN84ZjsGGe2z2APnvW2zNQs65o1q/OJso7w3QFbddaWg5
+YABRpJwq9g9gU35sBKXpkj2cYkvlj4U27durITJrp7XIFCO9dIvHvbPB/o+62dk
qNpm+EtfMl6FHCcbrRtYvZS56ThNWiU3+A3peLHbomqSVScvL2IV3nqk97zSNWNB
/R88k9fML8rbBEMoiNLSbokKl2yQXAUfmRcJA3GRO4otmjBBKVXPelyQXv+EGKUM
cSY5+P8RK0BMcCEUAoSbekuMlu4aayumkfTm3Qeip+6T6NoCw6PW4eEEBoPQqmwX
x7XLMSBBEcgCQqIPzNcDEsE3uLcSs/mr4iluEjdCgof5FyLCGYj7UgN4SDOEtcb/
TSUlVpI+Zavmp3niQ8/kw0j4wySg+UzTCfdKfO8oar2/QVSGHj83N0HcSsb37eEK
ZfTHdfSYS/pB4zWKmM7VDj1z6NxzFPPFRlZkSTmb/5SB+2/6xVpoYnxzq1Ju0jj/
yfdaA3+SO+zJgsE1zmDQbVTcID3CWV/VY7h4zqzP1APj/puPz27Xw82rIF9kcwJg
Vh1vc1xi5DnI8qxkFiPz9aoFO8JjwVAGAxdjGX/ogBtfn2QpVqQSsADc0nruR+Wu
4ZqHPg+ThsZ2O4viL8Lms9HY1PX0dwORwlNFzHTacD9GDfK5avBA4R2DDoTFidQg
YUafbuVZ1WmfV2CZn3wofdXQOcdWedkh1YF9nY4/3CPZ4CCharqSktRMBBCqQwUN
wxL2m+KbOhrhgkXsfWNUU9qHpfuUx8zZyovgbD3Lw2DNNLwkVn6O0e6BMG1rNuCo
1hLfeooT4btzh1WDiC8rroa96E4jAUjQ6Or6/Rcs9WHxZPMK+6qu7l+asksamTjO
kOhmf/Obwih24LjYnNRsXkRTNZ9i1pfV9lz8JPwDtseSSYCqzU/JM3XH7a4nlY9Z
zVwYY/X6JxeX6uLGpuze1irp9CgHhDELhAayGpxvRym1hNjLo+zccDO19ECSgVfS
mWTveixbwPIjtzhDKp/cYPTEjRJDRxN4QuDS7gA09n10Nah0IMObpeR8Shs4Kx+b
y5VAVGNbGmZgtcwy9jTJWfmFKisG/ehKvEoQc1mImGk=
`protect END_PROTECTED
