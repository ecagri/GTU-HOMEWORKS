`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k9WaceM5LCtlD+I1MQNVIVnJdqCgX8FJGw7tiDG54l66C3ju7HiEQBlxC7l7JkRh
ugM9CFfaUh3ZBpl+72UCiwrUmpz1uRoDtAtn3GU7vmXCmIDaLXixZx6zxEUbMaBt
723Pfit9S8uChJWMln1Lf9kRGKaHg6dx8+OSAdHtX8B/bHieW2wX4f9+olYhkCFB
/7LyPkHR6HMewY8B7SklufuWvrHr8lyr0LPAgQGj03aUw/k3+RR3wNI+So6Sozlj
/mu/RIcMxk89ajE/FmqWa2Zi6W54N77cqVZupK3xplpWCio+foH6puMiJeekh2AB
0Q7WAw5n69LcU32e3jvvkswApUXlEjcioklMrkRn/efDKhIOKBYGQ8wh9vymNjhv
8mcew9RhF8wKCMKDCHYXC61U2E1CchlZuertg6MH3AJP6tBz+Sb6YNLZ3dIsmDMK
lVUPE6RdnJCyUwJrtuKPXQhKbkfsmimpPQvWVmLnOYogHzwEIFu2XGaTf28uTvUV
oFYaKclMISLueYn9c6VmsRMSX1pdvMAWgTAwO4qm9xtCMg6Wi5yw5saEyM0bW7Iz
/v+6CG0EZnim3ODrmX4Nhaa5Re4/dqYgODfs9FmXLCxYdmBP1fXYgIl4JAsHcXzZ
jdspUydxZQvQjPALFSva9LxapOgY1uZ1RUkRMWEMegAfpXrxGpT2DIG5hOKcLs/G
CdrOTI7E1y4l/r1Zwd7/mna/urKmLgqB0F7xr1XC1C828U9eQ50X9Sz1VOPAe+s9
RJSrV4NqgAVfUmf6G65Mj0PZP727wZA4BpFly/z6PB7fS3CCl9PRQzn84L/G61v9
VXYKuvblAVkZYekMRCMYNj+RyyguKOG97rAhyzaiJAKuzZ4FP0wmm0NnlEjhZqBK
BOSRGQr+jjMpDxakmkyEyqhxHuRiei/KI7KH6Nz2v+fw1L29v1J++yYSy7h5iWeC
Ky7F8p3CBK0C1Y8xBIpvhQZL7pk9m7puA/CaZAtdvg7CGp73d6y6Pb/5MVzOnQCa
/ZFxKuW5xrxOcsRN41BKzdbor7PPBJjk48GVUaqhI/gpNxxCNNy9bftVe4KJG5A6
/YDT2GESJJcfBwY34iV1c3cz8/9ikFD/i7AmoNE9ER1MgjdsJeLCXQXAb4cYh9VV
/bUlmJ4Sl7SI71HMQPnentdm3A6YNs/Hg47qgrmKpMnNX7YP6koCCvvos+P7S8zi
SgQX/U4hYdfntXsK9EhgUkt3hQkUpDj16xZA0iKGQECGc4LNDlXXYWITfL4uG2VY
KNWYHZDxtwINRTCfBaIc+yBXeJKYdqSCSKYtnUx9MIZBTB9ER76xyqIckobjJd0o
j4exhZ6qdIuYASxZkLYKlh0xpUjaa8UKyo5IayLBUjvPXpSW81HDwOfjGIgIYpkA
BzJPojR2tP3k9d7v9vv1lIFFw2MswZKwDTqLzAXTEfXnBNKowuszZsTceFwCQ95j
z2lDg7DBYrQWxiK4tRo1TL5RurtFyUcY9m7XZBeNLm1puuIqQX4UF3wMzEK5Pkom
pl5DPK8vFJa8LrQVrETCxF5n6sCtP/RgLiSNPsftNNjbB9U+Jmkva8FcrVUXjQ33
eUBJXinM0/YAtJjit15Mz2ClTPWogC+qsTIRl7gIGt/MSK5LWQw2r1mIBM8CroB1
xo6Rip+JHQkXnmJqPdtztRYf6xI3+t3RWS115wI9ofo0ZTgDEXVpAK2M1uxYj5TF
czMYmGDU032uWvz+srHxujJpj3FGJx4SQcjcqIZzVbR0wSeSGgU2LfGoGpC270R2
+4A1XNPJYzXfRI2YNYEjIoCdHzvXM+HZgf1+pd9sGLDPjdAoeB8I8O1UXUNvnwyX
I3OWC8rAe86RAIglbPtLAJevAZIscFDivNGP2mJkE8qCrHcETfGV6U4F7r3160Wp
jviDSJJzi/nf1vqqi/Evis+XiiIvF4B/o/RgalVCvTVw9SJs5rWCY+4s5GdGgiwV
AkIvZo4NmeoyFDfznaXnrXNWMJUFy4XGf0wdF7RBT1AhnJAs6W6K0asQAvDRgkt7
T7AqvO9KFV5NXnzPAawT9On9z69Ajrmc1gVUxkISu6kA4kbJIS8qOYgWdgFQuomu
+dvrMbpPUcWUvez+R3WKU0a3dNeeDhhMwPV4KnDP14pldZCC2Y2Iuk6nvMAlgg//
KeZwGKiuZzkaLvdd6NoTOu5ojVJ+hKzIeoMLwczKAbZ8P5uhWbyt88eKBVNj+icC
Y5vjwOppiZfsciS2YhOR6ZaDqI1pKENGTu7/DezMkUciRtT5j8Ry30wfdwP36/T7
OPnJxVJ0coPhmtW7gMqy3OUhLsdFuAGQTYhnBdENvQuf/6PUKJfBryLMyz+55kyZ
HUaNWJY1jhPoYSJYTOo9H2f2YBrSjobQkIcIl53XQxljqf+lPu1wmydrkvgMClkU
xPjbG2W5mlDq1VbQS+qLMPqGCPrcukUGm1HhaWMM6P9WRJ6Lu83CxH6SQSFriW/L
rPGZgbg6JsOQ7YraM1QH+oWvxmWsnBUZr4DKzFaDBVDbXnEgRawNbi6owJ4IhaIm
2IUh+SzM7GXmb1m6qp5vK9Y+9Q/VzlfyWIvosLGOHwHxG0oz/3SeoDlRdlEXAbWc
/aBjPhV6MEh8YMeCy09hocwTpsCUohNFAdvpHXuIkBCi70fGOSgH69FTua5s6V9K
WTvmpc9q+ADD9sKMNKZ7MfXFDeIHS4jPzvMzHsh0eF6LfZ2B4Ojd+8K0quWVwDnX
3lL4l95LCLQpueoCWTLvwpoipwtjhEbO2OWxkffSyko4H89V5aigWADNpbJ9Ih8e
E3gfSmdS5a4ZN6QJ0oAljHaCm8tqdOomnbpkEg+KPOCteoIVF+V1dQa1HR1CMOHz
+IIVNQbRmJ8gN76K3Jgiomb5kyb/m3dcI3J9E9pfdeV70iN+Y+DM6dotOZpSBmQJ
e8CNUMv/7wVzOvEpkaq4IvtfKrWTFjXuVqDKmT/0bASEj39p4XedggT5Z0xnJgf7
f4fHMAR7Oo+taARGTtRpU+jqUhFh3wGJ1mexJFvOF5Ive+I5ax/Czpq2x9Gmo0w5
AYAMd76ANCHWfO8n7YKQlK+/oLxZp5Ci04C7BU5RycDfToOX4ogyFov8Hz5uio2G
cdc63FQlgjqvzr7AmOuK4OcSmvvsPkxODKmKtZSq4maJfnUC+9nZX7EuMZY2ywMY
aCBVxLNUSUIeJoRVx82prKeIQafy/UwGbuRqVG3FemYKA5JuvfOf28EsQj430Xqm
TDfoRMcI9tDdEGNM/BeGqzPAXgtFJnv1ip3XOPqfY0Rucpbs1GTHFlE4pzuF+Wmk
cbSJzit5u+KSlt34uQOaMdGvFNggWB6aU3E+J4usJL2IgeC7MK+3pzL4Q093x+54
FYZUrTowyv8HbJOt3yVaQubIXN/n/mz3s1JNz/DoFUIC8bTsqKKrSXhQH09JsNLk
uCQrgPGFI1oBBthXzjF+rwyjCPsxOjVfNJwo/++1mQpCQn02lj5FyYIu/SyIj3u7
8AgkzT2jh4VK0mKLUBAEazCXVJgj9Py3+0geIeaInrEpHm8ZBuEBPqGYiUQrPPJ5
N40I6is0m6G/sqWrAnKtSHQwayUFZUYl3nrpwZmKZ6OY8viWaa3Y+2j/QqUOf/5R
FH0xIGv1vKwIPAlY23gG0MqimuJ835B1ZKWt+UQdWlYZIkQPhn9dlkAnEPAS3gtD
YNreMdRjKUWojYly8tYVdSP7r4nTotY6gnH73T4lwSsjmgK76fyeC7E/DgC+HFAk
beEa3AzSSmvv0kUKpjY4n5iWPGVE9ODbpm236sJn6HamcJ7uiMnVDVpo1d2NFIRj
ylz6Fz7oc01l4tanjuKe5+HamcN6yTAG7Ta314OOLmnPg0gxumpbvUC3FjniUA/t
sIDWwClHY68c7S4+1uU25kpa5XLsW2j4SJ2N94o9dV9iGFUUQv1wMLUN62zYJm0f
Rr0zTbX7RTj4NjIUb0hkRSsi9ja2AlsP47JauovamutWUWC4EV7nQPt9UGWBXTPu
LGsCpq/65LyFaPWcUggNddDTOI9Ufin1i8voDaeAasYJw6HW9utsjrA1WBi5m75g
PO8N4IN13nRtIBVxA3esS9rqV1YdQcUj1jtBfJDrFPfJqW+krUh/fbDF3/nf77SW
p6UUMGErndLXd2R+xP0NxRIAfr9WDGcEeXIQ6PIHfYEXQHn30UttmOmXDx9bsC81
/6S0ASBbFV7CWObkhs0vD6T83RN1tHOYqyvBCfDN+hm41OzffxOejq1TGSP1gdpH
DbcC364ZcXu89e0ZZT+ZIfVtOgqLdoomfg2wio2sZohUjHvZpVhDq/bXhx+ViDf5
MO0rwqKVBo5p9VTYmK7f8W587WruI5FXqIl08XKRq4+mY3My3sZ3i7WnrP8SjVWj
M3wHdpqwbj8y0UslXWqbfBLTpBIss1yvwJdz8QV9YybZq2YqfeOqagWcqYvqO31n
AgW02L+GxPeJLoDGsTRP/u+SkoKGaxGHbJWZYovy8Jxlh9KmPpvsnETsnhbbxs5E
L043unlaixxJmpe7niKO6lTGlrNWJdjVG4m9oKEMg8htDc3h8RhDkqCWxYyJjvf+
PR5EzZSF8Q2Vfx+Izdx9aSIWrwPVnAMyiU5yL84ZEUjo+s7tJPqW5cTg+6dSEIFT
LfEDLXAhTO0TzUjuNYZkjx5IiiCcbl9F0CKtq/L+ucAamKYKhAMBYx9r6QZYYqkP
H8cI7aNGGDh860mDjmECc1PsKUCrxkUilX1XOypWRCQ0opFUSoZnpRSVSYB8Tgmd
cU1nwxQTdQMJPtKkkLRw0G1H1rJSw/1U0esueWSXbjWFeF2+EM2ITnyJicGaB05k
+LgP/JFsjw9b+H6vyWHl+RHU7PKzAG1wUlkYEdjkLddbwZieLA1KQlr0+cj6xG6z
4991G85C4ouEOO7wNYucMnZsl8hGmF8wtLWIQIrp/Ala889KJS+GBmI4nrfwgtqh
0sFXxWZLmaiLluQmOz7TiDMyLs1GakyEAE0XSxqFASPAzAIbL0+/lhD8KPub4dhc
qC3Q5gBUhvpptKK5YoA0QR/wmcjZarxLnJm9wqdck0g5ybIM3ThbiJ9uJeVVCTMu
kB2Q2lA9ip2WK9iE4iCaBcJYsQFNIXvPwQFKnN7j6c+pHHY/5RchfA+y7RG6NjHO
BH+LoKLjFIbDHssn1OdEoRS+3t1RkI11xlwj6x8KA2IhAPoVy06OqG9kl6HB40eN
0p7V9uM3bjcVp3/aO/ch3FF2Kt8v2iF0yQVR7ndEqlUErkcnrkQgQ5c4Kcfe5ub/
tTA+JPu5jNPv8BTo4BPXwNv7/leJpjKZ/2u92nhcppVY2aLG1ZKJ2UVwVv2AzDuO
GvCSllNFm7aYkyr9MaYSEySUn2B30RJkBSEyuO+4CRaB3kAw2m5e/k7dYd4kPC8F
U5b+xesvPVnkhEkYZaMlwPXx94rUDdo1xcw+fD5+L9VgrlOtoeRacNtHC+Y3HQHd
al1qOuQ3bLzHNxuFWOzbUrpu4RymBsMnSH/VGoc80cdYtSGOc2lAVbJrym8t4uY1
WxSh3C0bCWo3Gegz5gx5GuhIdrm1eOvuviyH1hbwpVJf4piJq4pBwwfMb2X/k/cL
fWVcaXeW+vZ/G1Rj+lxPV3RPUaeI6XNLtMXjQF9N+lRld5UBCqz/6XpWxUEd8Aw/
Xw/nifopKRQaV+ZFpCAAiIoq8tZIHSJQEpsjfOT4UB0aPLJEw/XsnexibVty4Dqu
KcfHIfZ471h3pEnTmeTAVR9acFuTOug3EZ8Xm3sUEKCkQGjmAyzWUWPs4efzo6wB
Di2R0R3DPRLoML1FJHoeLwmwsaq4YRuLJI8IbW/HXaxoKHb4RSimKzYiO5UqoCAk
Tx/ryzBc6d/EQ379YQR9fSOb6CZBrkuPucDs8/iLEZhTWt/0t/g5ifBqSycQaqXD
yVveYRBE4AezNwjtUHPiJVh+ZLb7ytxDkdUBVGTcEyM9EDkqvXALNnvO5eWXlg4r
FFsCvNsrYUcZFmnlBIk18UxQI4UFXnSUGZFLjgEVposHytvB34iwxZEtCwenXxeP
FM4vhFKB0uCzcV/XrlhY/7ulhwuPVfXRdn+pzLN2i5RZJa83MPZ/KLKadAozr60y
o9HU/2yTPTrSAu7nhjPATExVSsv9cPL3OXLIRqsvNWY1rvxGlbEqwFw5wmSTPH2d
jOY5caTW7XCojBIY8B434MC1VoQkAp0Q5Dhy3n+oPRqBNvlOY4U/Faq3TuPD15L8
3Ai5JHv55SJFheAttAa6OOFhA7AMzcqYPVD9KibJpUGG61liBHCZyOg+dinbMrMM
4ijijlzeqHehivSIS9cBo4vciwgrHdBrwhu92GmeEoywWnfxbPwsUG5AjMSG5w5S
eqdEskiUk5DOxCgqsW4PPHLUcDOdIEKGUniYWyJkuLQkss8p6gETwDhUKxU9dTwm
nqEsrpRN9jjHE6uph9cYnRR6prtKxQn7BfX/1WBEMqqrLj3gXh4gJidsHwwWronQ
bpFusrmjh58Am0qCkwsPmbcy3IZGWAdoJx9NA3lOkkv3khUyxNIpLoX7lv/VCn2X
TO9fdx5oOzO2gghixwPxSKGgp/XE9E71Feof8NiaFbfytlwzZwCx94yTLklNT3LY
GTSHQuKIRkDvUcysMuP4aM30eW4UPJsNmFDhovdOtvZktiH3hekHwMWSVMXWSyo+
YoxLp9kPgp9Yq4FGR/vJSzUIzQnX5dzdVEW6duPUX20=
`protect END_PROTECTED
