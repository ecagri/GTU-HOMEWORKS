`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yUjQuaN2wqVJdJl5/l9CJ26xrHoPn5bUZO8kKmwY4euFI9iZF/Oun1M3KhHXuJ22
cFSRH/Rt9b95yJBdx9BdzQLjfA09VOM90jF9e9OMaJUiZXu5VkddPMhIL/iB+VWr
tXCJswLCQL9EnkgzdypyXWsEaQIGbaPqa5tmNVQNbRtHKzvvdg3pQCIylzpcGHKn
ftUMega8uqoam6FAiMpLEZGEEUQKDRTNjFVzUz6/VeT8tshhdxBgcsYTUE/apUj0
sDPpgPWzgCRbCL7vaoIIWNireOWT2vF9eEvB7W/uqYtDBaJnVgJRgo+kKXIoWJpG
rvc8vhYPPLapl3N5M7Ozm1WvOakaT4+7vkxI9NtE8O2P834RDb8Xwl2VyQOUOjcW
TDZfnQQr+zBYjhnXtU4r5HI0WE8eBqoHr9vjA8J42fK5x/I/v9pJaLPWQcxxkpda
3fvWTcMHE5R7UuSH1w0vjbtyDcYtF9aPREItdqymgqfKzwbRoMXEC8BZLbimHmYr
VAEyXHsCRpDTcipNq10phqWptkDJEEFOuQxSDDY0LlnPJPQ8pNrnspex8Vci1FPn
eEdT7GiFM56gywHCcg6U3B9s8knTZwkV+8LTGVks3c60M5T4LCypGJyyBhTpoo/M
V9kOgBlD5rbaOdrHMwgOhlcDSIVVq6T/RUA0FoELkVo+ifD2Gdy1FP8o2kFoHSEq
sXQd+NcefvoVqopc7RHFyc0KpKINeuHUZmgyrvMgX+CYhCueLjWjSrK4YdTw02Jy
UU8iZeE/Ifz4imshOp/pn2vb+70qQUrLAeMcPuE64R9FgMp8vfd1OkGMJ/e5/w8/
g7X781AWf+wgy9C8w4Xx+BMMGgUR7PWJPYNCW1k1tIGCFXyrM5oFxeWtGwroLvo1
qe+6/m1l7O7PelW6DfCEtxuxgib0LVfVm1SnttwdkkZLJYBD03utdsQUmifegb6h
WrMSVvUh5E4L5ONUhUd1gBkj7wJt5DZT+gdqcCa8XW2Ux566E0BS8rCX9xJeAoAs
jRcLZXjR5eh5DWs75arDPw2olX7Wj1wR5B9cmKrPWqe33MdgbjTf42yHbLg1ryi2
`protect END_PROTECTED
