`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XEaAjv7Eq7hAzyHhCapav4ydCn/G0gdxx8T+m2Hnhl/TwWZfLwub/CJI06HdjfUT
u7M93xDxzrTyPgHaPYjWfnGYRqEvAbmGyeHalPoJlyODJcCF5tYWSk3K+ts2peK2
iD6Up2NrjhtaSGk/nDxHo2CxC+SsY8/XUKiZyWp6B33dDhYRjxEhotb7VmJ92t8o
PCAY5DwMRuPuFGDuQdukADcI5Q1TsI8X8YBuiG9HB0yL+qf+2442qpIp8Fq0q0Pz
AEJXb0xrQotcOERPh0LBLez54a/7tBy0uRfq2h+GLxBaE9vFP+B/gvi9QLM4n93O
3wFxLwh5iQYipm5hWT0c/8vCC3yOtcIOuXRBse4wTSm1kKIj8DD1ghUx139YuIUF
s6rg2iB5rysMGdTLHGNewGblLB8tRwBTbQxVxfSRuYxf2zvnpeod5vR89vSnhsYG
/7bzO3zpnDCrDQA9/icbGC70ZfDAIwOHNH9DR58HzCLmwPZOjC9CJBeNNJgJnIq2
2pwn0w2kgF8k/z4Og6EwZ1LPvfYBF70aRI1iO79eSdN4ielSODeoii+zNqpOSOP/
MBwcm4rndQ+y5N/W6mdBg2zHdQXNL7pzRinkZk7T1tlAHk6sLMr9ekXufTfUfHiv
xQ0BD2TQByvlFKuTVKD3Ntk9uHXSgtTWIOP/7pu67NuBkx9xBOYF92y+WXxkgCZI
83YSyTd5njy3ArEiXRWhlSO9kbMQjOWiyFSWYcw8iTU=
`protect END_PROTECTED
