`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cGob6aAMaTSbPfrfvddfHFpIagwwxNbfMKjNBSdvvUmjIP+fhQAfPS3MNk3ix5LZ
zZuvFXbK0X7XqlV0hWtAa/4e1S+E2hkxDTz/SDDp2WZdoqV1FLhN6nLo3SHU0vEI
sOltIAZdPMVHpmquDsxy2qsWCFTy6iJme+SKjM0TQhhA9ws7DI+FxlPnJITLdV0X
ujzkUILBEF6doCSn09grIQvDN3OXm6K5o72bs1Izm3G/ZZeFiJBi4b/b0qmu91vp
lSbUst4Z2/q1Aze3wXTnnOjnEgXU2nZRQbWaBF9inQJ7gJu/MU3+qpGtV5qZBZHE
Mw2E8ekJzUbxhg31y+UlDbDuoTOmINOe3Isk8cK6+kvzaUp/c091WkmivY5oBjms
ZEB752f+APPy+MS1bgcAGn0fEZEbTYKnUQent8JmOngO9yDor01CfTvaFhrVAOo+
uASMUZsMSenzEGcU391fzIPO8fJ0xNyBCeexBWpCudHLGKr73INOMtVTYOhsIA5x
jukKR/X4gDnxN7kpx41ALCTgSzHkLFpgIq3OyAi0Dk2p6hVoXfzhdtumEAXhoWMj
d/J+gwdv55RiYeXZ4+lDsq4a2TYYdesNzY4C0JrN7iJkEhZwkV2hxLBRylq+d6DK
BvwgU/eG973+aqXYjScQKqqOiXBacfvQkXm4zI7lG2HoYCtMkRd6n8yyIVF0xqJ+
tOUPox78p/opK2DQeDU6qyiSovpOWQ9evERRvTM/O9KobtjGugR59jNUEGv+zonI
wznsIkPRyON98aGR7+9UvgnBB61QDM3A/5ANDZCJcJ/l6K2bn0XJFQAzFKr9d+J9
xvo5391w+eZ0TGDZCWOgw1KH0mULmNr/YgEOwkRcJMIjdzNPacgWgHtkRewmILnC
DvlGvu0kJOrhwaBbeR0k90chaDuZsEKhGTpGoVoayeWyr6To2RwVlaMyiMBaNg+p
6B729frMakKTXnYs5eLpvUC39KBP3ybWbfaeBJLtQDkI/sWhqO3XOag5nBDCOMep
bzMJiz7Ft4afQKlbYhL3GENCRfGSntJdt7fddd0IyZETZuvb6yLboIV3xCuOvy2Q
0yKojJHujnI6tMvXRk1/aa5I6zhMkYPnpvRmVOE1xRpWgq1ks3UqnAg+ZF6yDELa
Oq8zoeqYNcwpn6pL0jHALEyyhev2Xze10bM/MNlHPqfhVXG1ra3K+BDMbC494+cW
JsXBAeArwUOVzwJRKP6gyWIvdqmYmzoBJRRQGVVV8tMu38FPEYvAXpGxzlB3hI9h
y4TNZTol0SYl6UL5qJsuzGDlKvtvGJ0Wz9KpGjyPvJZpLOkfghrxpE7aE58HwfgW
T70fNwSqaKv1I5uIaCnE9LzLA5BfDyk9GGG3ZhaGx6vc9WQ2cblZgCl517I6nPU8
O1H+nXClmI61a5W9dFIlkeB+Uu0zR0+nqPtC7NbJfP2g9ksY90A4+xgrJIWPs0rs
k0f2N/WFWwWDgPobpUjJeDcFp/1NeevrnbsVr1VyYfctNr8EvfLAeILOmTwwBZdv
lzBhadB88oQ4zTs3fDlQR0hYSQPGWeWljC1oKyUZk1p2UTtvID+QOotXna499m63
+d7W/D7yjKCLEI9JYSoNSTRYOndbceUKE5NAYhK8lCFZFyVMIPutT4d2s5Tno62g
GFBFyh44VGKLKICKaWg5aWXb861p3Zc+DW/0IKihT4ZELXH1R9QgbiG2JP0raq8Y
YifmXzwl6UAoLFPKrGdcT/epZwg7TKnKqNmomMmsmQ00EpIzkAw0mweKC4EChmRE
hIguXo4smKYTRspNSqdZndAoLLvz0KkLuwavEy3+ksmZpDdJ7HaBqPvg85+xoO8y
h+2h6HHEKQtbD2AivZDlUKy3kGQDNYPtMzk1PxGCFTH7KqimhGANfskKZtPLH7fv
7OVri7sjyEWIU3lblnYNWD9B4hNcWjHkJHVLHnvkdChu6KL/IkJ+chjTZIEV1otQ
GMtAZeYuRf5iRjQGifKJ34z1rNzN+pi7SlD7tnvroOmjPjGkb0uzLjbWLP1uQZre
hLFCFaTqBRYS/fBWu5ydb9DCfJPPKIAJs5Ftj3ALD82kSKCh4R5Uz23QJamJcBt7
3B32bqyr20P7ias+kl8+/guPgIVZL4Xl2enDqxbw0sG3BfY+AHOvX3bmUTkkt1r6
tq4e/DyvJLnkVhBDH2KbTWu2bSqhYUDwBT74yQxxybkFfhIfu0rChROTAS5+5G3E
L8PXc3PiX2xlYOmE/foukg==
`protect END_PROTECTED
