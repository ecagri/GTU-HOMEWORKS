`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zGvya9hmCELNo/8cgi4BnWXsSIsz2h0CHuQ6QjfdpoWIyuxRUHD/50fgZTuLqOVd
x2aeckCe/ChBJjk+lVChsRRHcEFzKDEcjchZG9HhhE5crbUyzZVoXFquYj2DFXb8
5cPs7Ixw7n6Rq9MrZ5UquKNKfjBsanhCKtm/kzn0oKa7dPhTBn0RSplSuVs2o73r
gY4MSgcNm+dEHsWIO8XJxLgi/axw39Srw7PjuioxsmBWY5jFQGSIGIFzlnuy/Z4z
P37Pux9sS91cgAmuyWA4MiPEqg4l/mxXm/MACcchPgoKKngRDEk2+v1xRZ3+RFL8
qiAgk8GlClaXDkT2txVZfuuDHbn+wYG1yJXX3Qz5s0fhOa2p9/dg3sB/ZFgIx1Rx
hDYBmN6qVyuRg7dxhi3mtFbEWSdmg9BEW9Eqz6Qp4xHo41QDTvj0x0dXBmyHJ+LU
JGzOTF6apxSTyFLeQd7MExbEzrzFjFEqMahflqpGgNQG3xLVuZjZS9ReCkPeOMgT
kvdEIyC8qyHj8e/zbQAqkQedskcIVQozjZ31aS6RhA6J/ujk5PuMeeyZRSRqmfJY
YlyfP8ZcNw6vx4C2VhezTGrS2qq3AiSiBcaICmpv2GVL8CpTQ/cYoASrgcC4kAu8
yclYFwOEkvVMBW1ZFBSfH45vk2UYKwgd/80nP5VmQHPwWJNF0fPCcJwfFS1k9wl5
SKjaEO0+39cLRZXi6xTMf8jdf3xzuTygyicnJxXLAUfiLnHK+E8QE+tQR0+UTK9O
19Vz7IuflelBHGZ18Hwz/JSmbCTDssFnkzSA2cdrfGw3CG8U+1PzLQVxfVvART3U
8defgeySFz6c9AU3akK8osfvto97NUx6rjEDD9eS9PG0hZLG8S3EGdB+evfv/COc
MHLpMZ2EA0QPC8uQiKdnFRr0ITapRZmlYHTy5sYuB//r1MjvdtDcA77dlmLF43Ri
GSE6omgx58ZK6AP4fr5WEbi4CsAyHMZGzhIrH66JKPaNc+QjZoMgDMQGJk+GLcn3
Ur8whTFGYQN/YYed+pGLypO76bMZn2JntiUax56B/pK0wRlzFF0C4DbdF6LvHXku
9KPs6IEWF3cfl6Me8TG1r+X39YQ1qzpxpJffGD4lsvpPyYoH+5h+D6AgnjgwtsEt
RJ08bzVjN1thxSW4zKEyosfkXUA/Lgt8hxrRxlymkDdhVcezT0iHQPbNp0bw0nKA
/oP4ZMCuCSanPx3bV+VkzQQ8OpXY2rXvSeIOW1AaCW72PRtlfqyIeidoWv2gpsJK
ZTzQAwYlGLVL1C1BO+VQwPZuCoW/OTPB7iewlRlzZiDUoixyxzR0R2ShnN6CpdTO
uWUjLKS6HFXYLL4O0aS9yET5bzUHPmU4/Lv1mvAFnr+8ns18GIdoZBWtf3VyEtM5
EVqydL598f+mSDfxfVA1Ig2JZqzaVC0AmGDpu5KCFHmGmXgd630aewZenUbeQbb2
iWAMYf0tWYa5iVNIZ0biChyk8IGkckRiIqzBbhtO+bcMQ99begmhisIzSBkj1beL
vvLc5O0ihshPnHwWfPpjFrVVNRLE3Ku0W2/9aTcbZt2qyCph9CbrZXM2A/K29ufc
JqSfkefzpPFGC2Kh+teYFz3fo9ZFtpno1UWUwnKdUqJ13S5Wc380ZuLP/vSl9K0m
vZhAnap/LHRN+gLOlZ9dhfbhWe1ou7orMnZhZv6SXLLetE5lEP+ALE0duWoiORoO
nZbVi6xAR1x4spZGFFK4VLQm6QZggKT3L7macrBXQce8GLBidRBu3vz0ERnQ1g9K
bjrov8wHGiyFnqUB70ZIwyuvHzrv161Ou2SbzHwuWRHHoQocvtsBQ40ubfHpj8JW
aKgeM3UANGjbRy69uI2d1qtdx/PPrOQbTIMxhlcZu33S4XMcElTC0SeV58ZxmRcD
`protect END_PROTECTED
