`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P7Un25DpMWGwW2nvljxh4IUZ9vVH+EQFZAZrvzpZ1IzbZyzL6+mvl5oytDNi4W04
hcCtlBvfqbZsazEZX6kYrqYxBzNpJHT8mgHj0snw9ULFwX4yEZ2Dq1UwsfWGocy4
lafDTDtRis3gYKwsxFtCKoss+S1A9m7gKQNYyg6eOK09CQso2zRnCWxJiNDitg97
w5Wd64THntZWCTGP8hiC9g+jaNrbTgBZl6Qca/ZXNSI7/ycezVMv61FFecun4Maj
mEjBPAxHf0Aa/Qp4Xldmqx6Z9hmf3T1Pcz1BKujHmy0JQWeLYhq3vYuvMnF5NPnP
gCOzaRk6VCs2uaYv3oEzOf21MP8Za4Dqe4izqtykUHkyqp+1AKJt+Eq+zC9v9oua
I//EMDd4vDBYiPezIi7b2plz4CW+8+YzZ946mKEFYYdrfxoovmSEa2+8eKj36CSI
XugAMyh9IrnVy4wMrW7OA2s7zff9geQi4p29x7k/yGFqG4Z5rUv/b13ofLQR7hcs
qxWLBIlmAthm4NJx9CnnGc5IXLQAGQN5xF0looV/JriaE9ayX3FJeSUsNcZOJunE
VrhUZotllKo3hAnjznptaO3Jvj/whL8a4ZdtcAXW2n+Sqgv+LBlK3dKcCfOAP1SF
dPH7Mz6pDbmscY282dBpjccMPDTbSDBRh5l9RDeNcJrEeAujrfKl2UpnwGSnsto5
IA36laKkidHGawVCepjNja0wylhE1seZqKgU+LJUBFR1D9XJ6+ipyYJ8hvCZDL2z
pp7pC5wtlaW51dBeEoS9+CHwQ7cVV3D7QKCkxfVWJXauHZfVygvCo6MuxDB31Ss4
ikuHZAaC69zHnaCI0Lhy8ep00ceI4bvwsExLS7MjitDEMqud9k8hlupBUzxDb9Ue
uUtFup18u3/sgcJdgMmqDsVkI2+UvfXZ7eVqY+Ilr6W4ey1ELQ2QRjCohzBNrkR3
purVJji043p5Juu9pNpDU+ZpT4Q5z7HlpIsJVfDOvcaO8ZjvW8b1iWkt8x1PjvUs
YC9RudxKxDNLGig0iYbq4UATrCtMZIHx/Hzn0aZRC+FEXkRuS3JsfedxZAQiQ4z4
SBCGPe0E0CBSK1c27YM76SIGbBZWnn5+VoP0bgLSpp3ysBDkyBao3p51+c+UPJzC
L1flcyC/zro12sIXlnrF6A==
`protect END_PROTECTED
