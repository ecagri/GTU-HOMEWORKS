`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uW0gCOJKYTe+1Rx1o7lPIsz8KRoBBmqnZteAnvY7OOesY2HR8at1XHGo1BVW5obS
O/iU73b0Y483ESqcc/0aR9dK/E65VnbN1L9UVINt2d/vcw12iEyI/v8SzwZgFAqs
gD5nuihK/TcVhvbR4R/ZmNyY9iQ3FIeEi7kzv9a6OgowMSuWi4bzeH281ghua6Vc
VdnyYCbvIsHd38d+QIsnhvmvWc251N+KAnGUMmWLeRg3BS43TTsHAabzrHRMHbQ9
s8f8DNfMioFSA8oAkzIclzV2CBwUKFHmmdjJoFqRM67iR12A8zCZ42N0kY1hQMmb
sGiQa2MykZfccqiLZbih7RiFJYxwecds03FXlPZLmk5STe+nfMBotor1br998F5T
`protect END_PROTECTED
