`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hrUv+NTPPPIHJKcXRmvkzMQw4BdypBQ9ZaK+gY3RSTfQn3WOpLekHXzlA2j5kz7t
c8xkbLWhYg7vZnsI3Ro3zPuU1M5zRsreY2gai7RDY+mYVBn2feJ3iKAZBcnKwGXq
snFnIVdxyKHLwuxIIoUWv2kbGjSaKiFOMNLMHoctz9IQ9kGThOaC2zx0YLADyGLR
`protect END_PROTECTED
