`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kXfZ9bJ5PhTm0tKIE2NW7JRpxMj52OQZMMOfw95becgWQuPrvOtcf03qep0XcJN6
ax8kQVvPzsYMoFehFeWkpLBrSM7KC0faHjdBpWn7G2mdHPzFgWhw8vLX5xRrOghT
k4P4GQVYnBS99u5dO5pap5IDcXOEXGvBOOUD3/ArgnX2pv3nww+Aa2GvdV1scaKM
Hrvqq0rsbzT83ldqCvdyCIAKldlICbNqv4ra6LTB9Nl8QfrdHSdxRFOjVKsdh+sD
zpolMZ2PQMBbSl86wWFJPZ1XPzUGEIDgG1NIu8q4EaxFDijdtkoMMGb+fSzmcNuB
jEIL9PTVNP1wtqgaDoWlOtB3oLdiXdTTOQKcWFI/Yvxi/rfZCjfMqNlu1xSqSuBf
ZeJzzQuvMz6JB9q2F6zvlXfGhClVtB6SrMDRjpRiyUNFMm/Ga11dfUrSDoFQKe5G
C5mplwhIVGvEhnAnRHqKgKgkOAgR9Dsgq51FZSeJ0B6c2b5En7sS9/cjYKS2X5fC
DsKqU9zJKKnTmMOrkCUxHPkw5URfHPM3GphIGOgHn9pJG4kPemT4C7WEWSFm+/+T
VQl1KCSDanmiys0VdV5YrC2s18zm1yMiOSEeiRsZ9Kboq5tclz34HBXUacdXRvj/
FSW9Xu9Zr6RMy9i4R6ju359Bp20t2lUH+gA4jQQCqByyG0+br56iOqJdQlGKAp58
WLYc+1zZnLxahhMfjbgbJ9mMEcBCfq3Kdv65yGHGB71lwAmRpdfFNRxapOKFDOKV
gvJWiLX76xNSf5rhC5/GMOnp9bd+25PVcr92wo3+Lg77wgprXKRxMVu/Fx8y9Xvl
T3pXmejkx1mWNBJPhOenO8jkuZRSRac1Vu3ChD1RSPoLtfHznp/buTHxmlgKVwbn
E5Jsy2yvcEYkeGGLo9Ak0xvFtZPu165+0OD/IJb2SNMa3hkzY+Cqsq/5DUQ7C9va
dANXV305SMkyldOi+kcYw7nze1pMQiTPyNR9ZrWU+2JWRywNJcPeKWWxR1F1yfSz
7pYpTnDNf2OLNEFLQr2cc9G+eNWT3HDNzB5uOQsPJ7OUI6YQUprQOg8w3jZwEdmN
AVgb7BPjqDDOFDcuWdjwJx1gaTQOifr0DCc7jDs6abVpbyjXGkfYKlR0qORbvv78
TGTcncrMfKKD53gylPx94B1QZrxBCQ6xVDi5Wh/j/OPV3vGL7OwTUxAF66gFa2hO
TMbN1+IXjiEMmDljXsIQwayc3LBCzQPzZngBtMyHtyQpzQtJlYkIQE88tfSEDePH
EomAjrzHVnSaWyTsZEkn+OetXPhu+eMCVIRHm1ngmKgfwCsCAehwuz/yk8FTxZuw
iE1LOCs9FfoUU0DAK84k2n6CfzUuYxSX0FSALvZ+pvwwOj/OPrcftOhl7YLFRsFe
pjvuZh9p3x7kcszzP/WifKE55IFeDiPBGJ0+0XALsWLHAbJhLcOqqAPUodjQdIXa
4CWQwBXIPk4rwjYoXOSsD/HYda+mJW+bAYffhXk/+3Xi8Jp7mUBdlU3Cs27Zbjys
9QWY1vNo8peky47l9Ifp2Q0KhJqybmuTikxuZH2zUL2gXhQXOvSci2CVEsxYxSPd
wS6ppfhJn8/EevJqQ9+G/Vd5AOEgnPcSmcsSBa4m5Xd3fWFwjml48Ns2RpDzCH/m
OCu7zhvznHxV4OrFITxU4qjQ18r5zkhECtpuLtuI2u9p6SgePC+G0pFv0dtd37Bb
x9PGb699F8lI0U4T3mSWPMWhGwt33yTuJRDrmSqoa+J01FxYobBLGlyhWSTmCQ/N
Tt88mJjF2Tjr7GS+v4+pKFxc3yYtxmMMsivNMrR2Bke4HxPNgtNlz5JF3Y10y192
piW0Wd17aMRSGSX7q8AMZeHvW7WnyTiS+wGkKFD0TpcAFi40jzqtQGoeFXhU972N
wczdPqK2ZnkOsFHGYIWDkEYgwkGih980l2c6ne3oyyhtdb9s0NFGsZJdfEdD9Nyo
gl0UxLdgE5OIXWcyfonjDoGMb8f+60XWw5ERJ/hgc/72lFS5cYnUsTo+Xo2FKWai
bKF63smGL58zQOe5aMISFGjRw26ShejM874t00YSpveYNF+EjHR9oM0ikvzBsQdp
IIaIxlQgwUrqo5omrQtI4JD8vfj/uZ97y82pxbbRAt35jZsIqALc0m0iy65L5GnH
/APQ/xu3nOzxLfUB6r2OKZ2yiENKlI+R5V5RY2190Bym221iIe/7fuELZH2UQ9pg
q4CAvn9RQoQDOhFPm3PwsVTOLuY4XKLYju3TrkW6vBU57TAfe1vKDrnBzQZUvJO7
b+2dxDqK3MQQ+bus0hWn//pzVdJEkF2lWtrwyjaS0lpjcBfxQp2hquFh0fF9opzT
pIWZCVCkpC5OQB21SKbj69DsHB6SxDgcOyG/3XS0l9xB+ieHab8YgQdwvIL03ZC5
xNXUbFbNYAGuRgQPWdYYHDAbzertel8Xf4RxgybJ3PnKHzzb8264QxzuhwAzr5OZ
yVDeFEIQlcUNMVlD+0zgZMaoaxL2p/8qGZVV8LT1rRrSuaj7uqKeqA6BKI9qqAXo
mHXV1Ragd7GvXK8G1qqnsS+ES5bsfxjlhVITv60TN2R/FG2CeaZIKV712zqQJPfM
GSku4qh1eZzZbau7S7g7MysanNw816kzwEa4+T3eTTT2fwm/pRbRrosuaWlAn24p
4jdxMM3fG4yt6ytZtvX0htLISnxHPntSfzyW7LqeR6R4BXApPnMJLKLd4wYYpmJH
Ey64nj9rhhJ/+NdjkjiBOpMfMN+W/Pv7X+pxDdM0ZXevadNdSOW0xuDTUkQt1LnJ
XBxpY3zqqlQ0/7DLalhiG2KWcxztqyE30t+GPmFQ7v7eSIuO+vJYDGcaFIztpl+h
LGutl1/ynJenmEurBl5NyHoiCCbCYyFbKGigzuI/S5xmZrUf8dr83ZTOkAiIPgyl
cWKGIsrKwCSEBxXoCq9Vl08xrgT55g4bUS6ee7lKShJ66od7xbYTigCgpm3NwEME
aMOZCDJEuBAIVA4S+o7uG4z5I8Z2bNqpTZo1vq37fyIguGBjMG+34DboH7ZtkI8E
wm2wItjcJIVkOjAK4uXU3xIzE2LbZRAFlzxVUHS3dlh1BAZpaio1L1MpGDLB339r
WXkL3vtBJEzQidbdwvscB6EGyPBUP9PgXaKoojsdCQIDHSV3yH2v0kutAyycRw2g
N/hNZzfGRxdFUcrLcIgeGkL9iJE5msU5psutGl+h1cBlNM8hvIQT00EVDKM7C04U
+kUmtW7q7tn3E/mJ9yChqMAEOdWMaHDvI9JR9Fq9i5g94BHNUXEOX90ziaygP8zw
YluBgRh8SQjTxej4qIiX3BF98ql+8kdnTLAoS5dSGvTqBvmlAalctqaDAFWNhDAa
0Kxfa1G2XJQ7e3/jkAQvqoWWuLsUFsFRdRa96TXRNttORgaSLtpT4KN8k3M5dJfu
lRjmPZ56s9n3tblt7SAQSdA+J2HhrezAL+Gb+5ikKO7w3fKsuiWwpywTDSUuEMx1
IcIO0jTBhhc34OwWKPukBzLt39gXo8NOI4gna/HaPosOsF8+SJBGezSu5q/gIopH
KGQ7DDHJcC2Y/C+WyKyXOk/PhnIFaWE1rTAomkCdx211eOuAWdqCqHrEtEvhoA6X
wTCymj1DJh4Z+ht+Yz/WdHww5Lg6UcnuN1W42UJ+yeG6OUrxa5a7/ug5OOBKqYw/
7qqX+rr5hCIVwQLRkpruvCLCbyAa8Evw64oSm6ywS2NNkqUPYm8J6oKMsRaGI+rA
heAjlXrmSbr3+F84bO81YjXGbr1t4yblyPV23xy2Jy95DANuDPKtxldTa8XSo4r7
M6zLiBsfbw+uxTsJ6AQ5PHpcDE5WQ2XlfC6OMfzoty67tiOG0ID0ZkH7k0QHSPpr
EQeAGsTmgYvvV7DuarO2yguX7jKct5Zs4BbJQ2koVG9G6R8LZijzGvLse5elMwMY
xx/aSLmfKjOdkx9J5Lfi8wK7VTQ9IaoQDYSNdA0S7oKR+A6RoWGu2pJDKSNs5L9o
BPsmNHcQy6i9k6z5VW/7KmyigRuHoeuaGB4mWUz8YA4+fYOUxigDEC0ZgflEI1PC
FjyUjPkisKG+oqlcf1JCeQTwvf1ivINEoNGO9VNUHVOCOxvMKJkf6c3JxLKd6VFw
vDd0Yp1NHGrNnm8NquAUo4tHpRHJI1ZgFO/Duq/8mFvJYj6Ocz/bTUJCnTMOyuvt
K7B/Xt+tF9I9OaolSlkjCjxzdLp9hMe7BQhtXGShTbS7yLLUJXfJdZNT7Uu5Nw/S
Kz/Mg/lRQTiC0GnYHrp5hRDinRQHy7qfhKQdfY6vwWL/qJ95K2QO6wKra42pHUMb
0BdHCJyCBa016GtQ00QmqQ2lijFdxKyjdDa1nZFR7cp1VwB53hz5x85oj6f1eH8M
MAG/OsX5xjyIYyC24cYc4slmz2hljo8BRzatq6a3ZEmdClZiF+k+6T+EpaW+MSBy
e5A8O6OzJfFsDYr6AMGMW2lzqKt2KOWKbKb/fPvwG2gMvWfWLCc9yVKMdpQB4ydW
nl4gsOwIVxFFOh+0y/tTTdqs1F/ElTTy+1Evq9verLn5eD6fq5fX/QCPQzHgdX54
Jr7MpgPgjz1lzIW2hQJOgVDULUb9wMbz9cb8o+PyfV33t44w4t8OMRDWdD70z9Qm
kwojSgc3LU6xbCPUa3N6KNi1TZQDlSNyJJteKaYSsI9Z4WDVUydsw8gvC/DaNTVi
ytGqgV2dw4CqKRUHEb3FxAGCTsy9rbEGVTx9UIEpa7KYfiY4iuNVA81Ml5Tnn3bB
YguUm3QzlWNTXZEAdBwKn8wfv8vjb/l95GA3vhrkvqOkZDDAaE2nktGfxyeiqG1a
CGEda50m5AIJZbQS0nWO0HUNKWG5NxrE7riox5jtr68v20teqT9ya0s9JrOzDJYr
QgaPjYHzU+k/qG4x1rNF6y2L8zOCeJSAdvhY6EtxY/xFxIOHnAiN7Xy0Tu/tVVQr
x+b7STeimRhHU/e+Zl/XLHZbngIVOw1L87XwQvkQe+rtgZK8Imp6Mk+IgY7ZL4UT
r8KduzsQdLFsZpEvD8Qa8mZ4PZ81/Jqjet9t8oNpSqDC9dXsL//9yDJApQ3TS4/2
0U0W5pfhXnj5RrFY0gkE6aFdGTdosa5VarHZ671+MXmXPuU+Zz6gKAoT6irJY2HS
DqJM8MqVBI0OJkPOXbm0EpcN+6RpenbtC0KZ7kmn2lV5rxU6fL/l85dH/cDVeSCs
fz3lJWkZrNXD0oIhbkryh4KugEZDZR2WrtrvMqBCvCKt2KZHKh6r9gxqZkXUaHER
LTSm4jwbLnX3wNyRVXO2Efjy6m7xq3Xlux4dNeB8ExhcRz695DOmTeYjZxwcjP1x
AAPb9n3y9RyuhThjYQ/463UsVsg1KuhZVMpom+US7WD8rU3Booj5Zoa49/vEue5m
JwwVVRTi/+MLhthc9efz9LkUjlR9pCEgz5oeliWkhLnl/p5ZkcyCFfo0jSGQ7rPP
Udc0aZl4NF61axe+x1L/VR+2vo5uM+VBNfPdGC6CbetlAjF/uQwS5MIRFw2+H9i0
ezbPLVYCRO0uK76OUHQgqjaBnsarzz+qBkOfoYNf/nv/tKct0/ThO0Nls064MZG5
Y43hgXRr/olVQ6T4iLd/CvqDOtGUz3GOF8OiX6PYBmKaYntMEAs3jzJrV45vcUxb
FxOrRg1Uo6LQaAyO5mm1cyUc77/eU7Sd2Zaf2AHrgj5wEeL9nwwhQZ/129KYG4xa
9TcDoG9CJStCf03c7mhd+8UHgkip+tFV3n1hiBaj+XbEZ58Jbd6Hi8XKDIsGK/9u
g9sBqH0DcQ7+JVRPgJJg9B/7wkQ7i1OsQFkNjgJl0KnD3I74wZK7zca1evra9lyU
4LmW6xfsTc4mmqprvlDa8y0MFDxy/+awTwPoQnwgFyQ2Zui5FbKdLMQ94g7eNkKq
SGVyZVUAVyUeetTIO99bvT7JnO61X5479eIq77zNs+djvsxhK4L8Odobd8nPltYH
D5z7vNUVQ+SgSoOZfn6nMbbxSYrMgpdIcFy2/dMu75Y2+rpd3uY7JALl0otmL9iI
Mc1CUQPgfmRi8UaqPVogiABWAd3SP6WnMtsxxE3+J9F3883uexrY8cK/aVFD009O
wyaFiw+m735I/KoH/kipCnC6OQ0mSkEfgUb2Rl6Nw2YyfyfZECORblKrbY2XrLOT
37l5ZrE22YsN5kGXRxzit0G49IVXV77Yk9H1VM/mhA7aa3R554OTAnbshKsfIKe/
Zz/fy2mm+iBB91sSIk+LjDmISnnPjnzhI7G1E8T2DY+wfUgG3DyZg4t04htCAuNT
K9YVoU3pMUG1UiqKXYDig9rY+hiIVTZnLJRitesbOWWVm3faHZu+JkP+xHs6QFsd
5A9LUK3nXwgubddGTnthgTNyf9O6cweyQkm1ZNKkBhVq5mOnpiZu7ajMgz0vjRPF
mmJVztLWUA4uZW5k6sv2HhSkGnEhpXKc8m7zTnH/MUT4jNXRGOzPrlcUqPU1nujA
Jr/VtBvflhI/8vJSRw+ZI0NRw4sB65/CtdczKoNfjqSW8pHPIlDyv9qckX88uZws
Vv1kYimXlhlzwuipoUyvSdWe0xIbKbg8jk/NNyybWDx1iPZh4ppV5/PXDU2QU0lL
bKW/Vz7NQLN1q0mqIfuwQQkA3Gc9P9+6XJTJGz9q6//lidNlVzlAQWHd5GIdpQpJ
GxdumOxOE+HusD7P0SxI3cmHsDPThmIYrKmViSBQnRNk5Gdc994vojmkYpC3Jv4y
DBTwYwpIDosMOKujFQk1Y0l8TRJfLouDi4NKjr0IrrfxZEjJT5svdw5+SQ+QGxeD
E9T7E7/kGpu7UArxuwtkH2ULZZIRpBODlUPC0QFfWq5hDVGXI4ZPySLKlfL5JFY8
RF6myO+PcjoutaUZO0Kptl8YkWwiYgVojZvytm48zeVypHgkcQq4UKjy/vNkgp37
XDNVprGhrzh34BtUevjywsNJx5/0RQEC35M01rhoy0Bfo6c3fQd2p7qaD5V5TgNu
VtD57IPaeVt4ZNoHNf7jfu11jVDrsRypLUwWvQeAu1aq0urd45I4PamWgGsQRh6h
Ys3pPHXTCeqd0cC8uecWiPms5dZ01fwAe+1jkh8AUY+9znXk10e05m1TX+VR1clb
DSXroDIEyktrD7mmoWTOiigdB5f1SXoxQl7t1BwO1VnNxjDwk4Svfmi9icGHgSuq
a9JOhkm4IdoBrlFWtaMM0KEeWHvdbAuXhEfC6cFNdGZ1YPdGYGRpINyqZLHUFmX1
w+pw384ozVEhZB2rkCs7Bhel5U2dj2CydfhzhtpuC2vzuGYJWYO8/CmcxefpBQFy
txay3WgLXwnksNKqUcp3NnTz+ogpGxy092m0PJ/w1N/2qfaXBCVIHlO+Re+iFg1X
M7p3bzvfWbrHxAhGYJLHqZ7sk8F4pt1NiLq/4JmTbgeCF0l7P4CWGhkmW4KyYhj7
3TapjWI6SU/KmaBjMIQbo1OZhfTHu0eEf1lNAkBA1clOTablTq4uH8zfmgxIY1XH
AdmFHVhbBgFxe0SaOi71UQrmLmC0fTlnV/usFueZijruSTCWu4hI/8y4c1bx7pGF
tM22X7VjZuSAecEk+IcTds9tp/809zjIflPVJDuCC0Z5qLczwqPN/SUl6DZh1hoe
X7dYbpNnFw4/rxCpUoUY75M7xBM7ZAmiLFZjrqeKigaLlwDuxJi8lPE8TpuIGwk3
jnUYk281RL35BlD7lqBTF9eB42ZCu6SLPcZnnATL6ZzTnajtumG28/poFwnoYFK6
ALXoB9R/8AasMiTv33asYT64qfaTyTuP9SpxYZsaisZ3EajxrBmu+0k8MpDSyQCF
uuepz4VihqtyhslD3SH9SKWG6apToHIUyLFAs+AkLN0koJtExBqP0I/jTeEnkj1p
2pHSTRQbDlsPMhNCQBXBFiRr5s8skyNnvBXlicnr0rA7/uCtHaCizN3c50SdLte6
ELCWq6W1V0R7zEKwrwsHJhl5LG64g8UN72dhNGTlb/hjDXtwHrCu/567f3aLjf/H
UgYOV2UbKSx4ZPiEOcJ0uqzXIoFDPpYJ/OdIZkFesSwlFxc+/ILTYE8f18e+cH9o
0+h3JaPVpmdmVTVPRoaTuLVZ2sq2U0c8l/L9cNU6j6qZASr7XN2wtTt5xlpwZ/jb
1Bu9np3uWfsCi3B9M+pt2+0zwrxzakl8rZM8+ZS97awhqnNoU72ZokAVU4PYGv2l
sgFMIk9SHxGZLpKwBeRbcrMvNjM9BtC01vR+OTTK5Gw630nwC++N37uV3nALlg70
6RkdQ7qQen+/Jo2zzReDw2QgoJ43fufIQR9UCR72/r6yhEzkJlJSGsSHZxrUs9Vj
8XC1rJwVYhzQSQhuURRxssJG445Kgz52l6b+y9c9pyBm7Ot1okXw/+iRgORZ/bnT
zP6wAK9mGa5MJuSnFW8DOlI5Kr+FMZtq10gGr5wA86CoNL3dGygxI5dkXNNQ2tUr
S2befoBQUDqvl2VNICIy0NZPWtrsDpw71LHpZxMHJYG/Q2xfB4KchYHQFaPRgkxD
N4nRKR1oWF74X5C+QoZD1LTE2l1/OhIZOVwpxGBeJ1bssdrOHFb63YhxS7p4mNbs
9ouAzHe0h3kBoVs2z2PAKUT/ySdgcmNUTNnlqOwAouO+rAX3J4LKVj9EsLfBZ9EJ
uz53qfIOJqp7G7r+mBvhwmC5dBdQe3h0Kq7j5avrvFfL3HMDOvAedX3yLSN+y8c+
ej56WzyX1dK0MtuvYaH2fEpGYzcJrf/Mid5xcPzrqUpsHvZkEZORlX/Cduk71RUD
19j0KfrbGLTOeIAWgHkEE1PdznWZdAsKH+h3FjTk+VwYYh0VH1lvB/MhjHyydT9S
S8Kj0NENDKeT6L/fLYCK98d8AaKZhernmXwbpo4G+FsxO62Vtr12l/+xXl0vTPDo
QqjtZ9r5QUjF798wt/ZO7Gaa0T1CGQq2dPruddoqp5ipEW4KqNMio+ABhNqW/A7s
Sl99wOUTr899E29qThytPA0s3x3K4b4aSDO+Kbi/6FRdcqLNLjCnj97yMhAN18av
nRADpvnyHqSAJ3BwO0mdXoxX1lKAQin26+uX6ThEa95mwLQhKnE0yISC3jKKUaCL
MVPb6YszmKlfgco7LO7MwJtg97uvKPMqcRzFiiV/qfmQlcrQqG3mwvTnQtpxouDU
XzEpBWjyPT16YOvLqfm40kEV64SsmYh2epvfmYcwcXDBt7JYGJ0zgxiqScZq4KH2
0kdRg0fPfHdh4MZDSdw6Ij9PSQ7h0cZABGdXyGR8q4AnPeLrafaWAkOrg3kCASyF
Vg2OkWOnzygr6s0dBOpTorNYUA8klHf0fcI3P+v15U1xNG1gM60wQ/TU9y/I7i+/
EakbYpRzSQ5oA3xMsYoXjeuBhNhbMWox9yqUFvpPs3RD190TZJPgT1EPb4TOKvLe
mRhWfiemO4sws3dK+IGzJjurOVe8RPLq6BDIutOODO29FklLRkNR14E7tGjkTRVa
f/H+pVbAo/azAa10RUB8QFXbJkBbNWER5y/RVYOyLlZJUTqwkPetV5FFtVMwo95s
pibVGVWLYE6ys/BFtyTOUCfV6+L3Q+mYiUAal7nOp+8NZUjC67fwMnwpK2pJiQFh
eV691C7Ml5zguuwr42mpFh2t3c3sUzeKi62nGr5y5jk9BrC0sSKw8ZROKTuTk8AK
usb6pZIoMbKeuRePfpb+bFJZ54toyVGrGwdp8aWfGAtxG5w6lOXQFivb+lyBDcGC
NmAMjsFqn6LYVDSzev4RA/3AeeB5q2rs3iDmOxW3kVmgxmA0N9awxR0yW+WMSxBP
W2fJC4k3VCDO44behfQJaqZPuR2QPe5JlekCSWkteJZef9iJhd4I2ENO8X7gh5NV
kMBRYzqDsVAdMMxXm97pwTub+yOSK4mkZNWw41qAWA21HGpQSd2defd2kNwhNKqB
wJTupi2KI7pKwyLkbTf5gS7MkAwv8rGzXBaIJk9w5S+bh5BdPgUMkzXLqLL0DoYV
btIPKqQZwhZ31oN41OvmqD838a2rPF4IejvrSGsyU9CQLIfsaPBAB6/CWTTzY+6L
FZR72vMz/7Ow99a58mZe+AlZITcBjHzFGQg5KiU7VB2b5nfJybiXa7ORRCleqVUO
Pj+FjdLEXO9LHq49phA4GtWUoIei8rGdxNlL63/rypzSi+LA8ivQW6/fkGUEuzLR
sLdK8IXWh1eKy5RWQMdJm4LEdUstZrDjlBVWYkNfu5lt8kodnedeia0zWZdhRqnR
Cp97tMJbcFuOkUeeft5YyKR7ODovxr4tHwW8yGu0lUTH8s8ZJ1+WdL+UJBISfbDu
LkZSVaDJoPYFi6cAwito36kjrSa1R7uPpqa+PFAWOBUVJ+lw32REqJr8n9WAyg7R
vmnxNmeJUwCmQMQGVUZPzas2wSgSdZCrtz7+t4S/bVPJ9k4Viu4A43moQqM2YC2t
wPwfIZB3cVEl2tQyVkCBfzbq1K/XSSoI3RcMuXSNhlD/UciSDumz7K7rJISJH8X5
lykikRRGjAOF4glxBxGX4lZaOUCA2T4CHy/T5IBMUMXKGF4Shd4OWbqkChb8L4+8
7jIbldX6AVwZ/+Uu9bifHEKwB+aecrAPMTQKqC5c2Of8XzVitn2r7zP3qSuccvhN
ZedhWWP+q0cp1oZY6lZdXz4ICvJgcRT/SP/Dy9a11jj1IFrcmfEbBG+reBP1/NUM
77QS+vg1PMcTTov8o7EOze8kzkIDTAiZ41AW8/PDRcsGyDHxh1lsAbu3IESBD6xp
yJyJlcqqB3TmbbxpMdFcuNoDL7/6uwnUd/T63dr1XvMx5zrogRmA7nrWU2GbeaCw
0jYOEa3DCTlnyuqtk1RPskXHbBzZDM61hsZY2l7K8YNJb1MCniQ+zomQDdsFuSOd
8yYCblSKAwBbmiYm6bE48Z4T0xMW5OSlqQVpdCOvsuHkrM3TgUlw/L1PPEZb4wRU
7ByBdyYoMxR5z+lXU3df3fInzrepuKt5DjR3i3WlKgNsa6BR94jCBfzo8k//5MkI
dAUbBUUmzfOAEsGNYjbaNaNJmuqR4unq9YrBwmfCNn1rJ8nxhurtG2iCdoR5LsTg
bIh7aShmAFTCDKWESo3GIiMEefWs5bbTGE69wW3ZPdm6+aFN/f934A1wiBocrAiE
poMLnLfRQ2OFe8YI6rrB3CFXOxcIrIWK7efoK0yPEMBJoJs1IMCaejO29IAZqSNz
MVIyUt94UNeQ0ui1BayMpGsVVWIhVPd/k+vS5FcbA0IStjSxzuT+OOsSHmCowp6r
JlytluT+EBBqFhDXwkI9dstY8ldn30D2L0NXQzMUpUx5aw/eHXMxZNWJdpUmhzFW
NxC0ZXaFlrfLFnElU1eNgGs842+C/qKzv14gPdhGLTPqTHs9hLBhdu1WMxmEBv0Y
V5LFIPasytlBJKI0DL34u17x6QXE4l3tBOyhgp2tm6NL6BH8auLUHhxptupvB7mH
fE3OzPyH6w/9SnkaPojYoX+0ooheB+iqrJy+JFksEpfQE7rdRY1TGNUw0ajC+i7n
lFPt5qEzDY9bu0OLndQ5VwRdR3UjinwP7T6b6PsLpRrXxKvcm8HS9kIsxVdtzap4
N+6m5+CNtFdad2nW0VJpGcgp4sDrI/4zC3lZsVsu4kAnl1ilXcPdT3ZDOA/8Ul+u
GWE6iIz/IfFNv3Jrj84XVe270AjSuGyXYAS1seF/gvvBsDA2096oPdXl7uxmmZvc
VBgTUVjzEXY4NTM93aI1RRDoWoq2Bfvy8j/WkY2SsB+ztmS3WdnVFD5e3H7rqehi
4EH5A68Ch+ZlwevE9mI1VCJSgyzqV4YvKmcwd1rOMm0QFqSEhCHhXjshJVhJXK3i
BjEo9VgjpsWclLxsKHrEW3SIeH8uQRnMEyy0uILkc8UWpaa1+zYp07ZH2ykCEelO
3wdoJejo8EncLGZEXo+JfSG5bMAlLwCNy+HdNohx7anNgL3ESUol6ndbzXteKpd/
oarK4BqiIHoCGAesQyQlghV3MNP++R26ftWGyASmtJ/yWLVep4vm49/I6Cdz+DSu
GI+O6ur7SJU/MzS9pB8XuHHNrVByuekNgaNXnljeIkE7xsfZaeFyRaqWgi6NoHKn
jiLYTQELwhXa8foulZisD5o0EAzHO+QSSuSEAeEEmJ6490hPHSSHqaeS7onJ5o15
+d5cwf2zYSukXhiX27k0VBxZzNeI1o9OmEj5UozdM+0VEK1S6zNKMrJdn4X2S5PC
62zMuDhTHq/cF/aixfvXCiU5KvaLn2G/3wDskjZqZ97aXhun6eMxl6Et+03ZbU4R
0AbeibKAACufIbQbU4RQn5UtE67LZTcsqi4KGbiGKwTZ0VHOCF/m0eeiTb9nHB9v
2Z6x6tbAxUtedGx2vjcCNlQKN8YjsRqRWKcRoHUOKUZ9yd8DF5NcEkkgmyJ4KfI9
S98HtxzheqXuh6EQ7G02PInRu0VIGOgSqtz+9Yb5vLrP3E90l8PWGNMC3ryfUk7w
77DIdiTaWV+8UYXJgP3Ul1pfOp5nzE5m4Oub8A98aPvXufwy+afD2NhXRhbRQGH/
jWaDW0X/ABOgZmJniS2fM7GJ3xWTp7c9qR0m8CGbeLelgaHtoRP54vCinKtWh/ML
1BtKxBuaTuSwIdFVGY5GO7ap6vfzu6Lgmbz5YX7C5+lkV+6AN0lITlEMlpkg3HdK
Wig6lPTE01uJ/ApbBRJbi1Xl2F0aFsffQxzF8yWxZXXvPonjpZuR2wTbo4GLNp8T
sxCEXDn8Lu6gRwigWhtwjd5LHXRhqSAUhNzE8QhqWPy4zDWQK2eDVnvlv2045jMH
jslOS3XWqBIZQFUTjLFe664AxokdLqau5vOwYPKg8h0uht6DHfpOszVU1voQKkTl
SVli44YJSOqvyPXT0CzcQUWJCRqKF2UXKL3uYGxYMrFnmIuEs9WjQ4XHyBC+iX1g
bi3QKBturQEoSQhQKoXzKuKo76E4PXhQrg2lSpu1kHNieTFF5VlU2LDd7/+O3AuO
hLhsc384czLKFWB09sL9/6bUDv6C47noALrkxqJ6LSQYIDAyW7gL+rGIopZbuUQo
1ZcKJKHcDf9s73hF4zph84ep1juGwPss4Hs6FNrCd1ZgqJYx4cGoB0PmbHteN6D4
zCdhh129BtEgZcTlyLEHGMRFWCTVNFKSfCSkRBEIXfHlzz5I68wDuhbDZ8uWQQOr
xqu/PUgOOkwyi0tu7ZcpKAPSm764famN/KUZnlNkviZ5fpCtzzIkD2+O9d22r8ey
hWXEnSMNW+KT5SHeHOa1hgQq+Up+PnfRdysTEtOTr3N/rvSZvLPxqBLWuRvBQQRx
CXOap/vY9Dmoduh/ZWUKn1dq4uo3bERUQe/DQzRSkX/xDaZgAd4UF9SDszo/p0ci
2JZCYae5H3t1rtM5zbdHXrcvUWNdGK2drC5nH0YGQ7+m23nqbLOarVaYWWYrhYGG
A5kA88lZCdxpFfOGYLU11Thu8BNDzJwXzRuCvEStXpCTlHdXEEYHCXPbuiCo/+Lu
C2WShlMB2IZXgEWUkhjOtchDty1I1tAry8eCoNxIIqIyEkPnTBXXN5sjWoksiBQh
MJLFDarQrtWz/co5CCjuu8Gf1I8uW21/mb5SZ/u0oyaqVy5Tb/WWxqs0hhGzlZiR
vRZP8dwm9z0PkXidJJ+L0hHRMNYvdVQSzDLFUPX60egu2ZT6+V3E1aXXmTBwuqIG
okVjYzQxgbINi/e5KBl89tPpvUCrXFnwZonEGwnd+j+MIN09wps1xMMttvM34JxZ
stUmkaLKZB7zhv6444Iv+pfLYI/gfor/121VoFAU3GOPsU4VmivRbhvMu6vo+I04
7KN08V0vM+CPppyrZ5LWHcbzDr4xJsCC43XaksejEPRv+iliv0b8J4Q/LuZ1Gu5v
pgJUaIPJQbkBjDHMLCAFXOa6efTM2xp+b5VbLIJ999V9iiaXMz7DwldD7U4Da8p5
45fx5bVVDIlkQ+pDw2djfTucJpj6EMZGNmZUUuDbBe4eFwAAUhDn/3iFAQC63dp/
biWrMGj2xSdbitptpeJ6x4CjjhT1CmpK05SibrxY3yHEOLsfF9+sPDlQhHT2jzxk
ZWvUh3SjE04nUwch/XLFc2EBjsoGfgGQj/oGCLIc/pdWGNdWU+AbK9Ae2rWDpaa2
W9jj2aWRSIQuUg11n7NPfPOiLBuZjueNRtJV5OtqEBOE7KtCubSpVUXzU10fFaU0
5zNQA1njk7PErk4sz4YTggmRWjumwYtvS4+O4dpaiAFaij1eH5uJztxQ+4mANvKG
qF2zf37uHIDcwlzWZ5/v1yfpLSUucZTNdTV9fgsRMSP4/jhIt3n7vxy8vHWFQli9
r2fDTtwLIu0cE+1AauHbNhkg1N8Vfx3lRsBZAFkN84x8eO3MYR2kp6y+7/h48hNR
Dbw+TQ6fniUXmHkWBnmSjzK2ReH46QJfMwUcvfV70boHVdB2DIIL6Wqc0A/s7h66
CJxXkWmf62SlekSq34xP0vbf/5ROJzuEBu42UEUAhFfUsDXJaeyDuCpd9pAdutnk
5MHZCSfTNY/XCkx8kpVLUQwkijHjTGmOt2KisXT3dWPMhLwwy2wtDt4+gLIsilTU
QGemMBHLe0ujo8EBwhhhNliw39NtlS5kEGp++7gqriDAhkeLmpoOoRakfry/p3N8
ratxeZjwhMBuPmrgvS11nq6mALUVyPlNcCqeSwDHhT2K1VVZjKxALdaCigAcJSwo
BkT4jjpenYtlYpt+ZkaeszMXe9eQOGLjspFSSu51Dn4ekURVmdrskEjao679CRMP
on9EegD9nGMu7QPhnKpFZjbm2V2gzB2qTktmx1PjeckHh2LORkMUrqzrhOQmChf8
G5f86SGRtGSrvsyZMakCiJqvMvlf9EvLVFe5TykvWg96AIZIAEr9Sx5UQRL1jIHw
9PbQZ5G30PNvaZ9nl/Hhz8ZrM2Q6gtjpcSCWml5xZFONJ2+Y3HbOCKhUBu69LgHo
XesAmVp0kv2z7Kl2P2qXbuTAZnxFUvYRNzDTOCe1LHuF+bRIc3xqfyirOQEi2VqZ
Eje87bXakTROa1kvJikDp/MkczZSDiG03dOzT61Fl5GXeEDQIKX72j/MwDST7zgF
EtZ77Mh3/RPOEKBtiklyTz5Rw3/ZhmHviQ5gV53U/QE1ohay6+I3KKnwn1pSGFFN
pxEXvKpoD6YQVZMWxF83Ytq41CEtQQXt7GdTEACu77QLi80kNwOZXQ1sdOO0T2Zt
8HzV/NAeGNhUFnyAFOmPpfIMbc56yBt0YHuwKetOWWUy/4rZwfsFH/sTyc2XjWix
Fv1+LSLzNZq0ZFSVIi/1fHpPade1eGdPenKbyuYkVOCDk3mvM9ZUBrftrRc6YHd5
tPUEh9MOLdrD9QRdeDTIDZIBXPfXPg3LqCUXMzEHYuY=
`protect END_PROTECTED
