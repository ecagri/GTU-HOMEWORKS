`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jGCuFMfWPBsgPQ0iXwvjzjxze1UqQDL8lNUlq3i9XG4/FBPll4JwtiTZ0XcoAR6y
8rCbPS/545uAYSSInZKHSi6AFBUPE56ahy4CgHiuhZJSTJy5tLwZn3qETChkTmOt
GEkXeNEaBNNiNBLyGx6TEVw5ii4lsE+Y+wYapMoqCbVzo7X38ll1aU/vrgs7JE4t
BC/eXGSp0O6hCYFMeB+CpG8DI+HwnOH3mR477S1MHNR2uE8Sod01Mhp0t3zrHxvX
VsukrTagCKXzx2i4LdglfV3RjYgOm8K/PLnn4CKzXyqheMMWNck2guaFQwqFz585
Osrfq6csZsKgn6B4NLBS24Irs9Xt3fsVUc8CfZQYzTUb/Por5HrNFEzyG7Yv7O8w
1sORyswG03TAurFCZZRIYQRKY6fuZxXD094lKPRS96KwNff3+lCt6v2+24idgGrR
Wn1lhYC2bnEv2PiWcEhn3+d8WyrduPbS1Rv5H4p9ZVc=
`protect END_PROTECTED
