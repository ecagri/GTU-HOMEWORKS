`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0bN7+LB086ouNl9Eyp9anC7D0D+RWRSHzqGPC2Qo4nB5ryyqVmDcKH5yzOcFYfb6
VPNu1xWklJfS1ThqqhLlTfpDsQO/CuWCEKQOuIOlpvm0PG+JYUVAOaTf5SuHzdrg
C7tbmhi7c+B+IdQf4ZCA/vvBxHItZix6fJdbY6kId5hHb3rZqZl0jf4IJRCbaoI6
PbcLjU4GAhXZvdDbXAXGTthM4Ku4oksl/lKM/To9NfTfdPMYEM+JJCTwlRilKBsg
1AGQNzESZDPKcYNKXBpyc+ANgHKAT1+qO7nOsYLvi3X6N+8pm+Vm7rCvJNfDZivA
rauEI5UwvNk7lckgtK9DIPdxLtcFMyCTrvurk1qNnM5tHXl8vU3BfR3UjVP2yyOO
1Q/8EG785aEoz7Uh368WZ/hOxKtPxu7O5ufdeJADubZo5BDCTXE1DQLeSyTYF0D9
1QokZz7Sl8aM64BmVzufr4o27uRFzasax/LI3z8Ng8fDHXM2cnf0JqSMhbVAksoq
63Q6pZBugh8l0G5VXtBweyVAmAdIEOZxu/nhK9acKwk67puaYgsyeLDinF9DQcZR
DPqFb6/LT/2A8wRYU3aaPpuzgX0ADfgOhUBEjPbjw2KnA48rKYNk1R21yoXIkWXK
08BLLB4zMmKgOI2lBMMkGyQBadntLVQ4uZ3y+a5xcmmN4dH6s7SD5evgV0gXZ8DE
dncMqJTzzcZx1q8LJl8RJFMJjswY2eJdL3/y92ZiQkz09Zmxg6xlBx7m4q0JciTA
m2TUHEfv21MMtJlKr7iD6tHc2IPMIBPmFcf9HWAcu6VGTLCQDz+yOGu9J8Tdo+a2
0fO1BDvJuMuoiZZB0Fl98bcUF2iRDEoYGsbvzjCDX3+fww2sq6bGDVeFVl2DTHdJ
cZhuNpF9vclSYthMDSBZbm0t7qqA6Hluc+TMBIMXVPsY4970s4SSc7ywqx9RIScm
Gp6aJ0KZHX789x3Su0zPjlDFdsJjqZsnwJHaYhDTQRXCOmPXSKoPmiTPQEqL3T1Y
hsuuJa2rIc/IlarQOqzH8cpuGBVdsbrSHlc6pJnxCxSpxnWnurdim+j/LDuvlr7K
VconzpsiJnPzOjqX6lkTWcUYluji7qSKrjsD0+WICufWTfepaZca7w6dfT1iFiXO
td7U1Y6XUj02yuZZo8tKu8mI8L/bpCYuuoT45kJKNDb1q216DjTsMLFinDdFh8i7
QjDnid6j+QEg5T4Vs/2mMd7dmvXmoZ4PTpmKqXEcmX8OlspGipNWdt4S4Et0xDjc
PR1YnPagqZWZtZx5RJSATglIQqHo+1/E1XdE7T/RF728IGolcM64OlwlDbM+4lN2
UCIqVtU9SxtSm+idTyungJKSv+AyBRu3vw8VhZ6wJBytV/F/9bNBS4FqGlLxdoMU
8jNMbTrT2JkvGfb6L++jIxnz9aV6fFVUpR1IMCmKem4RWIdlds1AERj6r7tqaehK
2HNPWhqpPWS1cUTZxmnav1AUF8KBoCk27eX9tx/WV0tVCFp3+b0rAdDk3Z3JWYEw
uCzZNxdK3Pzv1bDDi9IqsWo6c7REgnXPmx33RuILwMWO21sOmcyx7zUDHA+JL8UD
G48Hz3aUDT5TjmFiBgeT8px8hAqI4y1SxieikCpH9xnv4bMF8x8RZsiXM2ZbWU/v
TXBSFS2xPfMmNMneChokbK5p7F55Mbf98I9eEhr4BGLAljUhPQBNTMwRGT3VT9Wm
KkcVoJPuR3pfBkaOIY2gf1fJuCPA6Wydv/nyqVbG9wGk0CyTYeUuSc+sN8+Iv9uN
XxT6DTRUSHldxQRvcwIYuIY4iGAMRUettCjiUk6aZBvfJtO2mJIaXe+HXMt3acr8
s7eiAeerBAXSg1ruLx8zUoxD0Rbx94M4ODfvMc441nzGml+4Yi5RIQoeDbY7CoX7
6QCsJZbMyD+OwWnQ7LQCHZW00mX6yAgTe4ORR+xFH678xOX40ArGg8DmOxw+TiDL
70/Ndj+qt5ywH65rDBSzxTQXjDx1iJic724hpo07ThDrvU7t4RO8qkwHBmwtyVlG
MfhYX31RtLpQGpsCIKIdoOP5djGKHV1Ru3WG1QWfNnxMrTRnDBCo6EtNyi1ZQ70j
s+jHdWp93dYZNIiblQ6qkWcdcmzs1Zf4StJYHNm+7do9dE3B3uusxFJ1s19gNISi
tW/ggzaWweXWh/eAMp09oCeNNzu9owRhx7xcQhCNbz04+SUd/bvbPk+cYhbqvLt3
NPTeKrjDRZ77/5nxY6cbSzRfMqvb/vkph7vdRQ/gi81hRo3ACn6QoNtWit2H1Yy+
YJydeqXPJDJg39QelYAKoC8UR8mgcReIb7k7YodWTDX5nYWGHipi8BTukiqSnMAm
378/KEY2mvvHA4W4ucylWjVbRKYzgCpQrEwEGgwhc5sg82YeAeVgMpxd53Up0NJD
C0TYnysgoiRvYMR+7KQtL0zBVCcJ7Y89qFEXWnkdPMVvcy5sUAWrwNZFqp1d7Ze6
f4gsqsb62Bi37eiK7MpaVOaEk41bLouNlkgA6yVUy2PqCA80evTBNziWPStFr0dn
M54RlyKC5BPqEAM06TeD3gmPoIXG2W9aYK9Hb6X1pMqV0jlSc16vzLXkKaLKnQn4
CtUn+7fb3fy61RzBQytu/R/we9NMcUvx0jo6XSIRxGfr+ET2RiuG0Mnt0DWbPgzO
7vXJACmd9xEE6ALWZLMmC/7E43dZUDzCLj9OJV1xJhS0+DQFjj7BK/PZ+gGN9Tpy
SXS4ISS0KUhru0J4DCybRTfp18xKeUpaEfjqKHRg04vyV0zms7sGVZYwb3E8C66z
W/hBclyitb4LwWLEu9hJv6J5PCVlVzBkqOD7oT4Xp/Xo3rLB1PkZ6EuuHbmRceZD
fTmLmZyjKm0OsDF6sEb6sB17driA5rUS6j7LMQntI45DTMjcjMFTwfa2kG9+n5I+
4snVO0KVLC9Ck2CusnzLiXgxLwXYnYDsbJN37Z9YJHmP1LP27wDZGwSCeWIwPCLS
xzUiQf9NECRDSYttzVCO0JmDL31vXy+bfo4gUC4zSQJw+4MMygaTP3RdN4ziPOPP
N15nQX1O9ExyO7Yqdf+UOILd25A7ajC+aWacPAlOSPH0bDW+M1o/NTVeWi8O2Z0c
eMaj4G461AhlD/NC8F2ol6EKfkAjwwomxq7NHqG0Tf2UoAj+Mt5/ilNqfYKShPL/
9WArm8q7r/c7ecBIFQcCdpz29UkglD6kg6pezl+AurcnD63Hjv4o1B+98C6EAkL6
Cjy93JNSJIAy2wtYky7T8Q==
`protect END_PROTECTED
