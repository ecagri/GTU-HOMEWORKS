`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ydx1CwtSu1fiVi5doROtthg6c120xxMJ8snn6BKCqMhnZfIGTsRZ5/grmbYEnb69
I+bMYREXsFftXejCRV+e8MsxC5xGFSqb42U0U+ycoVTO6DU5a/VE58wn1SN8V/EU
nDS5j01ue3a5QWvdkDLSX5GwpYRGGuGDAyRbesx5tjuYxN/A57yn+Qztl2WNZkaj
6uRhgsphs9ZkHvtRgzJBjoT94l2voF/qrd3wZ3IIQVAwSgMgeOBvWC4hOoAEqsQ6
KGaJcIXlWx3Cg8uMnuPN2Z4RL8GpsrX7+3o+MUHYR5EOskVC7aNTOtXtH2bOESfT
y8vh8TCnPF4UAoYiBOaZGXANMQR6KsPVzEaW8S0U3gsIC4smS9aND+0JrD1s7r2i
RtzE2RV3pgCbT06Rf1Xj0U2uOeZLVfCBDO1AoRm2GQ7cE/PNXQW2702jLY1fONqP
p5SQUT3BCvXDeCAYQJX00Lu5MlJ6/TgglJGGZ6zwH9ze3HMYZOlBRSkHdn8SwdGd
b4zMBmaI0y88ygtPULmqtB7TQp1gY0rEhukuEYz1PE9gYl6fHgJ/ER6bNBEjqV06
ffjNnTOZtd96x3jt0uI1Ltb86bC4QQ4htEozW7CISPrgBTJGSYd/bvGwxoGXVtn9
MFKUELrKflzDGHFwEX7yFdFTsbXnlbQ5rE7WSAxOgywdL9k9m8LzNwvuF8ejRy9t
EqF+hHKWkVKE7U8VJ3YtRZ8+5pyr1KYoMfMLr9bXiPjaB3xlsOJrkna7AiD9e+3s
CmNVK7bvwoM3//yiUyb/xBfjiqgvDooIhZDAN3FT9bnxaKWP9VyDTTZnS4ZVo938
+UKeMGeeIwSnbGaro6zbZ5uGx0RAb2h0C+Vk7Nob24w/xfrLEhnsakiFjg8PxnUv
OCrNs/a8hE1Q5poiXzOVzuSZgZ5OGro6v+80E+AFjQTgNaXSirvza7F+E4iD16Uc
8VjQ9Ry2kUv5ZgSW9GagCTDQ4iNr8VsbMTyAGReRKv/yJDFPHbHi3NpBwOjvRlKj
2uORsXwGy1whqBL39M4BGAk52pgbmCBWprqQjMaTLKngUQTAGG/eZyvOqFEd+0tx
FbmA1w5MI4cbqFew3pgTa24CkvcvaAXlzfIxIj4Wpc2Rz38o+7+75Lsp/tg8RzxC
Zyvb3bdgzav94PXsqu9Zd+0h4FNI6C45aKDEBBfi/bgRN/Gtqo9bgPIRh5Nb8lnQ
nyQslyT6Nlpgwiveaxx8SrVPu81UxDN5wElpzskU7dwjocgpK2BvDMbcsEB83Oyq
yG0/TIF+5TDymZJaBh+55gCVHDEA5lSqsNxd6b/SQl2LWO2h57lYK1NoMxneAtYe
3gkz56rx7W14Be8raCv0dXLrKLojcQoaXM3nbUwpqfpoH/6MpRfeOJoSTX2jedW6
7+18dMPVN0DtC14jSEctOj5sM8qUcuDa6enosbh64iPW7lkIghrSbPathTo25SJh
N15wg+8NaIV3K1KXtGSwOIiIlk7Shu4a7SQ8GbeuykicVXdQ7RZzhagCBtfokC3X
A9KMbYHMytcBSkPUPv33xIKl29JZScTeRH21+LS6VBilbasng89O3Ym2E4wJJqVB
S1jQZfKvi4ZPm3LjShmIGifVOVDQvqbH0sVzVcD3287gvgnzcTzfVI8G1HoLvafv
4/lfjzSkWhhyHAYv1r9ttmhYJsmVW1fkwiP/Tg3tzeFfzTk/nhHpPJNGKKcps4br
I4STtFQlworfLMWPh3luLThFFkNLtYlSb3gAMyplzi535BZ5/eYCWEvxo02xDQHC
`protect END_PROTECTED
