`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vKIW43P9KLOqIFItUaqoFRfUkxCYV3jbn51xfhVmGPBA1oYW0ZoG6JKuR8gmlN8w
LLXOmE6Du4mBlgAQpOFtKQRKvsfi1At0aHRGq4BHfitLWq7gDNd0SrN31z1HDnqv
iNuSWUFZFoHkroCvTa+AuySB5H+EbEKw3rqBpNCSKcGvj+lahRUTcYEE3PsVvmft
Yal9GVJ5OV+ZycOXFbGw6d6lg39++HabQtA78EVDzIi5n7A+aaJuXGdk3ADGW+Db
QtBtQXnXFYeoOyA/ji9LcXR4FEjagtAYnWzA5byq1j7A8VDElx7vvnGgVYXbjKwG
guTEysiUYyYGdI2PDVs5bCNPoTijyij6x9flLASFfc+9mCtJCTqkSONoF6WQs9kf
L0Y1Kg5Vd8yPx7pQTnwnnmSGxgCqgegDjD87qj6q9mqPRIDCluGxOA5cJK/uUXh+
OB2FX8/WH8AI76Gftip8g2UeJY8eQrL2zOJzFBTmA5QHZDkRup9L+NYMRdyqKFb+
LdexAxqkyadiV9WmDOemcvBQNt1U68GsEr3RXHIFiJAWyU7ILzdsLmZn1o37GB4p
pSBRc90Rp56Wb3tVp/aivdEvmiufwQqUnYkIFjX2DDtkOy+1m18PlZnAPVPj0E11
AMWuKDR2SDqyVfWaCLWK0YqaPUdkEPzM6W85mdW12geHJYecET1J3dDPis51hd4S
TWeT17EBl4Bpcsa39g5Hj7IsSFfaAIlfD44aPJeo4BJh7yTEDt+nnor98UbvK6Ks
VBTdwx40uuRBF6gj67RFEmOaA7ItoT/T1qlbLpzXyC5Hcxh3VM/fugnX0EudzkKf
pAuPj+wWwEAxmrRoncZHSg==
`protect END_PROTECTED
