`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0HRXwDddnVk/iG5GixtamPhwz2hKXwVWf4DRwzOajI0h0EJWwUxShTPQ8JA3WrGz
5cHTaPZOPYSkECZRtKWQa3geUpjSQprCZYXKoIh9fThvFBCEALnbgv2qdtJGEW6u
fH7fbBKKKWx+qAf1HyX/gNgfSucfoBH0ftFalqgfkHn7rdYKvEEyDbNRHDfmgpDD
OkTCll+NXbMQADEO+Xn5uVn+xJaz37fJ2lFGrqDheBzKfNHeajWSgGOvg94GgPrO
59SqyG2oQgy29kE8SPWErAiEJ/hbRxgsbM+A/DKwovh1NVyZiwMcMqj0Knw4SQS4
89fe+NbTDg/qVRj3m+iJyqxvUy9u/eGOzQhb9xyFX5h2NF0MKluVtbf+Q6Gvfbm6
`protect END_PROTECTED
