`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z4UjOR8DBTIaZMDu04GqTVgDNnc2UFwy48e9VCIEfkXj35yvxyA0C3bt0omnCoNY
NG+O1AwNfz3ezNbrzitFjwa5WRZKvXMDSqhFcWmqwv71ICDNjbTkaOpR6utw1Z5F
uyjfOXGim9Y1gvuuceAaK4p2dKOefhx3yvMffJaMQXdfVhXI8V0vaveBibP7u4mw
x02gqT15on1EQef9XOetoHeWWvbyXiu/u2cD/DomkyqZ0D1MssZUr1c7R0LgLj3p
MuBAjGZ1P0JdgaKEMHzIBquH8sV3BU0UVTYKXEObC+r0vc1rjm/JigDdSvkbPvpK
xekD4YnrmmWbHOcwnPW05f1qBu9fM06O6/AGGbtfEoTfHYRD0V9RkSLHux40lFaM
XF5SbY6VADQLOwosoepGcyOdxR66cUXUwpa4rmdnApl8QEpKjqcz/W73sVQLufSf
uVGiA+bHg1w6M0uI72bTkJzk2q974Vpv0wGbMnwrPTTzSVPkRonf0ivtyoLlOrRK
VfBVXT81YW8GQug89Ek1o2v85XEpW8dF7zj1qtpLliQ3tYWQKFftKcQ+Stc0n4KS
gKQclFwHzY1CTTR30YRct/IdQI2WyYoOqfM/DrJyiZSn9U3aGsbaq/m4quUY6Pb+
AArl6wz8fDFmCmi7Sxj7JkH2LjlTalo0OwAs58KkRvppL8Ad4k4atoishwKDsDzW
SyLjUfQCoGYuCyEuqc1wPAcr3gyvSU8cQgtw4C4kbtdW+JLOOAOKn4cScVug4tpN
K1o/AN1MrLvTdzhuy3o1kDmp3QU/K0kEVCN89jrJf85Zf+xOeiwcK7csQJaFcgV2
fV2edEc6IA/aMB9UX+z/McXzZi7Sut9UoECe8RTcJIm7JURzw35XhU4nzW/KXapu
g0hHMe6ImcH5Ni9VHpsTYk88wGUVwxnkLq/dIbbMWakYwNeW//R19G+ZvevohdsI
zYyXvRA/OtkOTywywrzwlIeU4Q8ukpdg8Gz1r8Jsq4A=
`protect END_PROTECTED
