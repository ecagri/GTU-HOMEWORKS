`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/LUtAZfANOn4Fqo/KUmX7ELcLnNvZx8NboiXvrfKViMVZcTPDhYrCJdxRhQfNe13
PV4fg/oczSN/fJZW0XF3twhRCMc8+vca1KXjH+guSyzU50vn5/WcqPjBRqsJM3Id
0x4H7m6EpOs1ScvRk5WO7CvzUvzE7ZSLQe09AZhkpDXkVHuIuY40juA/kxSRGS7v
udTcsUhFs9Y6sEhHsOGRCCG/Dq7HNr3pZuWb1R1ydMoGAq9ECfneEoQoabSX2jGv
nA6BNBiMxC2TcgCFBmYFv6wvTWxzSx4QFYX8b0iKQyCiBH9gWttmm8qN+nc1OPc2
E+8gJqR7lhIQu7qCi4ZmP/mehgYvGqgLYwkJ7zMszA6uW7OJTLHLtllVZsmjsOPq
Hzwyi1M5rKcPhlxzTw+gJf3i3Nf+rcZMeVK9BAq+nXOKGhm16B/aBAEBaTmzr6Ui
VwDjRkgb8CKaZVjsOoxDa/aOb+O+c1T3SDsIPGjsK8+LOHqtZFb1wUi7puVYskbk
2YGOzvqk+qXET31PRRrski9RQj3/NYowCbbnOWdCCwIzEMSRcCZSx7UkwhR/SbRv
aZnJhfs8V5onHXdP6053ly9t+KA2qSFWvCAg+S2JkU5h1cyLLSlzrXLLAg6Oo9G8
yNAGFcc72VYEv7vVCgh33vsvUCLSDqax5+Luz+uY9WtXiXFrEPES8lNdH44WVsC5
WDJx38EMwDKZE8Eboi3y/WxLlR9Qd1D6dnfcjyYvlb/mkRzaQR4Q0tu1FayokyvI
MbvLfiprwsvkpWkbuV6+TppHDoNvoSQ4ay1rhHtDXpxdOjbZgj584TnsrAQDjWbH
xQn32KmqTbQRZkvj+cPpuEtqCIwHQWg6U/MPBYUY6Xs3TyG6TGf2Yp0NlCTiYgC0
CqzcuPJof00dgbNqCZwmDdGRiTGAAvTUlsw3o/9Z/N8zInUnTQIMS5saU8hNrAzE
7YC99MeiTXJ2zQ5zetpw1HAJgjIPVJa/qFPJrBcmumaqcuUlYa4bddzE+O5f+01f
YTF9SJot+GMcl9fkXdS+AIqOnbUA4r+E273lkPvuqs5dXzHDk/xsJ/KaC+2p27nG
XziTSYSEfN2gzj1Wd+xiJ8ckO+EOwxzL5YADVAi/ZsTUecbMzI1TSL2/ZvLWn9Ox
SazXCc4Xc29ojBZobKiBMEPPS574p+/9+nKLWYCcicJPz7HrCMrq/y3Y3wEbekC5
cTz+Tu/M5ITOial6rAj6KHKoYu8sG8zlBOZe6oGSGOMEIu4KYWkqRNTUeGhQfIzG
oRl+r+P5Z124Nl/UptJNpmY9nH7sYPykbbRcHI6ZMWLE+u58jxsU3V8rMAMXgMqR
HGqqqLWgvURuFp6d/3iSbBuaBOWh8q6sbYdS7hUQ8J/szlpq+TlI6d+kKzvdImZT
eBMQ3pmsvBD9RRryPrt/6FsN7LhB0JBKFCYZT/MRh0hUqx0SUytwixrzwUo0LSy1
KVsL2ZTTdnqJI++7hd4WFZpzE3Q4u7rlU7KiY/mBgWPVSFoV4vJ39uC4bnbY5uJ9
OLzVj0crse7QV0VnNDw80Kw5z2fZ/UZ2wWTZ+k31jlkJGUHQnoqFJh1A0pKmC206
UiX+0t4NK1lCuen/01zfC4Egx92MdM35VxTYj1WbiTbc2dhCDmA0nh5bO6nWdTT1
yY9bGWg8yvUKBJKw0D2OePtpuWTvVQuIsvpR44cXvh2/Qtmna1py84ozvAI/7T8S
zFlxyNG06CKAgpAYufB9/Wc2XKQ0wtxjZPtbIj7w9s1L1o9a6wOJ/rveId9Tk1d6
1a033xE8Ez7/DFM1sHxSDGOBj15LO8cGf7vdWDg4KAYqnrM3HJinGJkALOl+xqLS
2zDNL5r4eFbFaiUouktFv5UVoQ66e3/ALhOc0UaUyBv8Ug92Rwp9Ts8WAGas/Ao6
ne+GmF6jjni1GyR5EWCfsxL1z3eiF3cf2D7wyLG53wKtlNs2nclfkxJ0JzB/Itkc
QvddlPWx5TT9p8ih5UMAcQR+B9gOUAGuG3Y5yM9XWnJvwaUrT+P0vqw8wCCjol1Z
cDdRmrmZn7Xv8V0svSAzPHrKnuIvw1ry+WGTynlAcRaSQgjGOKTARH5dlX1lAnyN
DezNPmsRblkpP9EDShf9S1AAS4Yg+JqBSTuXLQYMNDoH6jS2rv3sEQVlPQaLHi5P
tfvuSOA7ZCl+ve+6iNyt/iVCJRQEdeU7WZP0D+mfrJBj6QOFLlGFMj4kGGbaXkrh
wEze39rOjNa4ZKys0aL2aIkBSpnCHuG5i2UxWvKiqi4jufsXhJsYc1lswGK1xp6y
s2B3EG6/q5axJ7crwUcL7+MjtzIb9Xl38u28jQThJcUjvnu1YYHP75eTgcwqN6aZ
p6+vc5tb1cnWIYz6pr3O7D4tFZE18uijNWARINF2bwFTLrM2VrCoMBx8LIRPU8pq
NWUGnE6Z+y4WtB1kJIImGnPyWU2YpqNozYKLgSX35+gCXMMojsiY50kFZSioZpnL
I8Gwpt5aByePo3AXsXNwrNTEiFWox9K3axPYe8vaK49I9DB43zO+jACoe6WlHYNb
k74iQ3vnDB5lDkAd2F3YKf8eXzrqaQw/+cZQHthedSaK8HaaLLsN+4/fqP4mBSkj
RZGR9D9oemmdBnE9UG4QwRuEFNRxpz7sscVLyRjQKYzOPLHFPvi+ajvkatGbH405
YIvJFPS92W4Kv9iPnCVbgzOXQAfy4hXXvvtQyrYFuXIPAhbnVYBXfrrOegveENqL
iBIRQNR0+bOKZdUrtYI8be8sIerH5c6uEcvQDPrCWjxzp9P/kOiL8u/vdk/Gu0K1
6jWWdl5bjSFN/U4hrxHBYQevj7nrfYKHuYsZRd3iMQ68Ot5IHgFTHLFNlyGrgVI1
2BOYiTjgx7wz+PGLcHY0IxuLROM7ZzVfKMe3+LDNj1qHEl5uGWorALl1+AkGz1SL
6fUj1zT3YU2RMcxiXaQK82/6EkmViyW5Rh2ITgCGkmbVIC1kNkGYQj5+GsItkQ9K
mc7yfSPQwhat+pc5+tNmIPTiGR1RDckYAyUoY4hg4LZTJ1DefTXPeTIx3B90hzlt
XERv0lpE//usZolQHRl005jX/9B3XQep0b7rhZen2OQQwqCS7sW3PSBWnV92jBB4
vI41THeksExj8SjAbZblgbVvxW4Jy8RKE4qIXJyzjTXEZP56DFuXPSUwR1IVVaaE
pvJiB6pwEDy/ywS+O4NWMm3SQJpBSWxdPRBevvvwVKPlXZr7uAYfCH9eVncYPKEv
wULX02P+CcXJUS3qr25gGMHSd+GUNCwsHxbxttT1a5Hc4hqwIorf6z1xZ9ZqgpW2
AI6AoTpOkwAneGI6pjpI/9kzvSS7wNRHz1p/CHf+W+hp5PIuic2GxFORfV2PzxNa
PkCVpengWFQZyAyh7D+Ho2rcBFYA5v1CEemMO/tgO/VFVlOONjtEtEkrO3QmlQwX
1DayN8UGxyEjIw0uK/tDhv7xWrEsmMbD3O2lEZZvbFGoLDqCJxeVXUB900tsAysq
gPJ+/CGjGu4K2LlLyPUW99j6u/ZSVXA6/HLn1QXDNT2PbiUJCV6K0yMWBPZDAnXv
cS5pPgIBg0DcIwZrMwA0mKwmgMG1IlX4T454mDw6eJmFl+Ka+yB573TNqJ2DaiBR
154H1Ca+eXjDiKAVnLR8CRN/gq/M1PljQ0y8RwJTOULgc38+4ebqsYCUYKmqR9LF
Aee9ANgS7Rc8DlmMIw4xfLrlMUq0lvkfdz4g5n+UfER+VmKI+OVokjFzIyOCeMF5
VUtwW5Lwv52Fn8Rc68p8Jnj4dosNOKmLAFD35pMYmdEuM5DwGFh48/ajp0RxKaUB
G/hR7WbAZaE/uUXwGXF8m+7lenBiwjOy/psE1yKmU6qmpu3vu1xhl/pVustHPsd3
liBI4qV3jAdvayAVaf0ISBpIvA3vzwxepbHPCqc4QOKX/5i03Yq8TiuquGLisO5q
hIJ9jWzftJSBYZY5nHGy86zSkgbusY8mggVVbE5JHHl7Nz4l5lolHWXVUjQzE3nZ
VoV3zyXlAMKlI05Hl6JUXiuPKOBGrM9W/Uq48fH0p+FfiubEVlOKmjguBaXULMLF
MHa/q9uZ9OYdW7VsUW+q261NkREUfrVsBTkgQzuC9yZ6TsgxXUeG7Gf+ZyZAeXP4
iL46IYY+RsgUL3H9umxYngln8YPYpPAQe3Zm5LlkSVbAgvVj9ck2sEvlOJGqkrlf
NPAzBfFae7phnm3SDT5SUQBfqCtuOXph17vSaqNB1yE0O2IMYFt2Yun+ndxu9Biv
zg5JcCMZyCJYo2VsS6TRjebIlJrrKPyBQxvi6UWe2YpcyfDJwpfzONanib2F7+D9
9M82KuTbP5CuEGO3grx4osgYw1wIE9fAjZJu99eYJJXtajg1qe+RgQ35F30BzXyR
yKvtPbdi9xZ/51KvGEgGR2NlHbsvr7C9UtJT8AnCXTs7Nqb27AhaOCeCyDD6+pDT
e9JDssYsXHraWLK6SSbK5cS2LSxNTOn1qBPM5gLE3e43JB+qPsUgCjCumZBILwUy
l80rC7Ua8TSHMOjZ4BS3aonVP7d1L/EfzrSweSov7ULGRDsXhrR92G3a13Ix/EhY
EH2TEIMOIfzSa/SUFiL6lknMxy1vfoE9FGuMc9QN3vWLAjjaVMjRErw6UEZYYcF2
L2Zaz2pKTsfbCE6j1jaFBtYwndVixLecUoXpA6yU6c8wPwOx9cXyo5+uyFBS55aS
CarvkKWGNI8ZIo9HTNGrEGyViVn4NcYUZlC3yJ98WzCfp9eEukwd2O/Bx/yyANVH
`protect END_PROTECTED
