`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uL41bXh9VhsSirDbq/1Vn02F92xLffAr4nlN/SSJ34GzGPX/ebbGm5A/QBWtJkQp
roobL3c62E1Jv4G7+P/zkT52kyj84CqD2SYOL4bJMyXk7coA4YrUGpro7o0Dzkmo
IvY1fSDkxrEiNe/fs4slaO/rYvsRWO/scrVlzGqHqYaUaV3ENziFPObBQQiiShh5
eKnO165U3y1OUuIEcf29FXBZTDVY7ron1ZvTk5c5kcKDNBEsLgjQihyCdGacd8Te
S0sJrg24+3ozUByKEVKc7gpGA8XIkC78SfZSlOa5iupYxd8nLkDcqEGZvEIvvcth
4Js9DwpDGt4UmeeZQWn7z4Qs8WPnIVyUrisJBt96zKD7T1YpEWZJJEk1/V46Hk20
SaGg6fRop854rsrP87rXKz7c07/cGElsRguWhNE96uPABBCXHhgcYJ5NgOyDW7tM
Sk1jgTBju9NRJd1SYs5P9N3vExz7GvHHFWmw78DOr2r0cNwf7VaRQ47U8fZ0AnfY
CgGKvx8lifWtJhJ6iPf/sSHBhkTfKCajkSGObIyPsHhEHWBEL+Kz7Q1Yt9eMUm5w
EfdXvZoz/XQvxK/Yof4fphvdRwH+BQewWUpEtgtgAqwDLpdFBYBi5fSEunQJD1vE
xCip+a8df51/enbFelU8RZOzgPzPx7HF5DLH2xnExfW/wfnVxrONySPngRsaOpiH
dMF55YkqZoxysCt49xe7EyWfHTOV9ohyfFu6rx+HagM15+5XoyEj4P7mU9/QJce5
GCYkgX9D+DmBsc6Qi4oDNWdZ+97ijP+zDN2p1MWnjGzmXtRcBSo+LTMxVPOQhK+C
tpRPnkgpoUlTV5ep/4eOmgxYdISIAOEW/lp3aHHp9+Fn6ireNsTk1LqfiAgAxJRB
ZaXEYrtkSFIho0gH/PwNH2g4aJStV891SXszIQFLowCkhFz3u2wrzt5zqwEsWQFT
NQMGo3Eidyn/yNO0+OwvD+yAKzAMY5KXa5TrFArwFJQ5s6CdvZRvBWDc5R1DzWn8
Gayrvc+cwCuIlsDve8fg7UfaGfv8mnbsuD0iljvc0YdY3Yd2OUSK+cPxQleONl0i
MaLbP4+mnchHzYkQrqmGniej4rFCd5rqFnmQyrlFVBGUQYHXE6EWp16B929ZMCZS
+txPGC9RotiiLzPiVVzohXVn12PHNPggXgPS0+6qsu8wjvdRPVrEKZoTeBTE2cvO
Dw356cZSL+lAzezD5pLS5zo7XaZo1Pa14IvCh+YpPGTYyCrzPZ6sZ4hO26PSot8O
gKnKI0N65ZcilbRiEFLYyjkyYfIvp1mP6EFj5v/RMhA4RimWXimgiILHMJNBgcHc
FwzQG+gC9LKLrWV3aIwx36NzdAv67pmPikUWh+43ju+v8ksyI+5jWCIb7NKN53zL
0IaZtsUrboK7xctTyYAarFajgXe5SUJFRMyUHuDI4yhsKSSCG3JPHQExRDpVRIIU
ELi+nh0/no412zLjcJm/0uc6Fj8dX6otGsjw/DhY6UNiAcPjWDPzOCRku/HypJt4
zMP0QEHKUPXO4+Csluq8/R15ZGrn1YBu0djWCKpjjbUHzK7bQy+5XmYpkWVDAoFC
75vz99rdH8O0L4rYHT5wnIXPVUBS5Ua1wdaIhK2fQ13o0DOMCnqBMAu1WhjSuCVJ
ddBjVzv8X3Mm/BpVHuBsnH65QnZkQMGN4NPFEdSl1EwNhXMgp6vVXOHTiOEmZ5GZ
brP7G7ztAeBFP2+gvQ0NTFqDkaHMfB1DQKSuEw03EbWbwkapvk/6uOf8R1Mk/qWZ
lese51XQj+FXc9ZRx83/XmyV+6ONDP2IBiPmPw/T5cxFBw7iy7vKJsPCUXGWGVkC
Jq4kyp9yBWEdPAnm8769P8/QMRCJHGUJADCkj0ImyPXTQ8QDE+vWv/Q+zsL8OMal
qkXEpdmgyq1Ug7ydIjI2uc50BySbsmjJPbTQzlfAemCOJbO8GM8EgiB31/Er7+l6
3S6/5rJL7pP/Nzl2SzLp4taqifdtdTu+XEXTmJ0ZafEucPblz+c3oRVJkrdXDSyH
jYOFt7qRkJMLg9KZXytT+ND/81I9jaOBHP8cFta9nYs9+9R8lv1zEzhqUeVvuYcG
yR8ZX2wFT0/UFpEcmlkZgQoDzbqQSyO+bCs6vnu8lSu6dsxENgzc40tKXzhdbiau
L894crd6nUfHZ1bN657MPgw6Gogu9RmcqiLDADqtF+psRZ1/q0BKC2WkkMscsryX
+VYxdFCsVPQHv452Qik0Sg8CvGY7392Rw5kSsKE6cB6TDB+OT0a0lQeQpJycB0jF
X7jSgId1yN3AqPr4EMfAh02RoZTwvtpEDSIuj2T0cvKsS4ONaywRQ5YhVnL8IGN5
CV/IEjdWYcWvNXcnrWKnSKRRLRUqBWm5VhI23XLOu+VW3BHuXoqrDlbjS4zhxZKr
PYFJvpOajqAGs/4mfvBKX63G0MgkFOEOl0uZw1FQjcupELWIgjJXFqRgyOWknX7W
waGuOkrhN6jGIJ2FtmCyL2eRf05jTWQkYmtadZi/jhSHFQ5EoWMMWu6VgVmYtrbd
EOJ7ApAfNbFRgbwFWjJhN9gmtB/qiKBo0vJWbRZmqhfiKrk3nZgGwuCJCbmo8/zK
Tdkp/Xp4O4REKExAv4EMYC6DlyrVDBVlkJNrMy16nHhTHxzRM/ylCjQoIIj2ce6G
67dRWcMjwZEaF69tc5bg2iSZ4/0u6zHd7SMbvCQKhe7cPE4cJzGV8YB+subehZU6
9ml/ZkcWaoKYKrPzGXo9VEhxAxUMVj1ml1+aG/Clt4rZhYS46G3gsPInp3O8Lq+I
WQt+9FJV7Okg5+Trk6PtwGARFI8tj8BOQ4U1mN1fuKKPlYlGSdgEPX6YKszDC8Pc
YA4fIquOZZi43ZkG/81Kjxn0a9vUrtMavtAApLJaLKJjN0g5IQlVYZsECee+uI7c
YDhobCCAyslVP2kQnLxul7qyAfH/85EqkQS29MdKaEFqO2zdv0TDx/HsVcuIE49K
HDGhmUTCiYLVIziZfQbK5Ac7qkXgsJhAZOZ5ZmofgOEQz7CQSIbfMOnVmbWKdY2W
KO62skP8aJ8Sir8EYSIZA7Vw+apmvodloDGZkw7zU/U4gN3wHpqwWyV/C8TdpAWv
crOJ4Oylu+wnTXsCozYCX8rcFI7WD/Grsu9P210jSSMrFVGBAr2chkPpXUMZd/a5
5wZCFDr25F3To7UkK9MlbpaNvOnD75t8Y+59/zBmzNIkmbwzauOWTzbS0DePu+/8
BmGvSV+K4t6afF1Xon6cCddgdud1xSEKhzHVq92yls9EHn7rztpnLDiIN6zk5A3F
GwHeCkFYQPAreU/llpge3AsCnO++VHPK/rUDCfajm6M/kdBxaWfiX3kObPgRZKdC
nVomc9xJefLaZL1HyS+C9v+ZDcOnAzLvBz5LP9HgW+6+SV+qftFUaNgJjML26PtL
t5gnZZiHZi56VDDafP0dpcUNuBpd7DphVkrzVhTgLBA9jLiLuosTBmqUhcUr0iF2
BJn2ZA+gR+4S8jmLIYqensGyCv+QrOwfamu8h5nhoggSv2IVBDTNFCS6vu111j1G
fs1t9fxS2MvYlflR7oBjtR4CA8HE1FJAMH+AJP8mb+wGCysyNP9QmYMNxF+nfiVY
tg+WPaAV2ozu5B4lEyGbNxW0dBZ8lQ5QSjltc5H/kR4iJynsG+eqxpwuHmivbwN8
2zG6nu+6eBBwYmpX+k6srY/avClJtQZpRk5AIcuV6Uo+EwSKZnzQvcMv5/bW1VcU
pahuKH3HRhTTRlhoGyH734ZKZ6fFAq/P2Pg9cXAPvMA/5PXmf1g4HidL2DulxA+F
q4Jw0T9DD8LCVfysMDRj6C1pUGa8azSIf4dUGxRY1Q7eG+uAe3IpRhM4RCFBBjbE
qdtwu08m+AjHZRRYMmm66L9z9YDOPXikMTPLvk4Sth9lumP1hC/XXkSnTuD1RgZx
umu9iPO8DvN4gXZ55ljdvgaaUQPc/oGKd9w2HNigOIUd8Lay4ZhNZMxMi/NAwhQD
dRwD5QzfrPgPHIfKRStTo0X8aSLT9ZH8EHNWhaa1l5LTsT+YXXDVw6Al0p5uJdDN
NN4LeBVI1rf5ron0C7ufkRyy7KkEzh9rRyzRKoOlJlHJGY7BEqxRm3xuxof3HChZ
Fwc5YCGaivvw0LImRKFSt7pfN85M8r/m5bFo9WkSmge/UULuuJeHKOITccbRzweS
X4G+Q7CuX5AMimJmO0+k9g==
`protect END_PROTECTED
