`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EERVGW7R6z9f9nqyGhpdRatfeTJqFn8QXnQN8KY2iRC32eY68ds3N9dNnjbvJPEV
Yghe1Er33XWBkap16OunKyJoLkJmHduGDyPK/T4t4/gkPuZkc28i2IHJ6IoEr0xN
bVwp9yQHGxuBwGnxLJp4wEbarx9NVqdji/3Q1RbcaBcyTNbzxyawWnjyeJ/UdeLN
bt8jlYs00ViKQNmyNSJbs5n0vvqythjjjAJgAQGGQbewcJyHMRnFsEi7dTjHM9fh
BWSeZ1pjcvc/NDM7QYGfEzK3YjWnxvgDoYvJnBwstkCkBp9cyc5t87tgRWmsn//Y
DzVAN4fN1pBFZ1p9V8PwoZdjX5qibsPcWkr8IhZ8EzsWfAf9vdXlpkTP/wnI9XuY
0CAqHZqrpX3Fx9z2o5NHvrJS1tvXi8I8qUwKdTT1H5Pb2kIyJQmCYtHYVIpY53OQ
wuPXuar8Q6GfyhXpgrzgnt3GwX9DuwjV5I2W5wUtOjVVE08RfKgDm2FrwvG4pbR5
L4ReZUNn+jkH6VJmLjpNmXnxHCo0mdsVaWuBk+4uk4eICAcT+AlqJANSwqCdngsL
kxfWppcjWad9lqvLTIySi0yD6a3IiWYWN6Neg+s/NEMj0nsB+ijl52eM3uvv1Sgm
JbmWGmxaZ8yc2evEYmdjkFMx+Tah3E8yVGvSjVXmpSglkDEA5dknJwzAHgZq3qmy
WEWjgqVLwPHnO8A8sVC2aNIceHoJHa3kknFaeULonmdUP+8yUvM7uLCYTpGRS7kN
F0+g8BJErGxa0ZRsnVaO97RM5krr/sM35GxVjgPCdYwuuKJyUnZeTmckw2aDWEZk
NoA+GFlxIg25ylepljK1y04aZj+XTXwAL6D80lnaS0Ao97c/rs9gUdUtOSedSEpK
x48vAUsmxrLcdjXiuzpgTCAsL/S224na3OprQ10/xF5ba8puP3FCSY7K7/76cFIu
n+toyvrl3iSa/wnS8fUxiLe1Gem5bikdTZGXUCn2vVhjU5GaZKIpp5WUAX7Wm3zG
GFy6iQWVzxgqtg+n3Zu1JK2Gy+cLDuGlPYwfRpDCTSTfhV+z12Oc1n/NAx7NwZjP
lk3BQ0tSmHvHBVWtrwslX3kUZchid5ZQj6Hk5uusE2GoshnzjOTcKaDUcvo93RLJ
BMH+LF95+YZ1mHaZwq2zXA==
`protect END_PROTECTED
