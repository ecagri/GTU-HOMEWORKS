`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zmLCwqypM4Vb4GatQDeeHmLcMwm2ywBoTuFoz93PCPJQsltatuIhIt9RHD+s/tPS
79/xwJD3nvhin9sQk+DKdek9W80f3qJaw/xAVfimMYPWEzQ5eUnLpekKDxTGtUbp
Xl8bSlRcJ/gCYvuXWTm/2mfMflJ27Vp+9w55dhLSfyJHXCuPZ0c0F42jZ8QAe40K
LECB6FD5zkegDIGCvUG0A2g8tDvSQf5nqvc/aWicaEmKiCU5I+m9DgrgeKJcGsZ3
c0ImYknBwC68HmQOT3uNvqitS2cpP4eKve9RC119R68Ibd1BlzRUTX42g896hpgD
4Llo6g7HYkeQOCWTYbTR2JJW4SALUk2WMOMtEqEEHZ+OXIk1BzU+YO6EaeTorIQ7
rnX9QtpZL0SWNAK/v9F/rdK8299mCvDgOU5O7t4EdFv5m6KpbD1s8qZ/OAVRoKd/
nXFBbMofaAUJwg7OVxG6dzwbnh7+0L1ob6qhPkA+jQaDFM1W+A4YfTNOtSMBh3bx
JQHfjMk3B/J/JNH8Bs7JO7oL7nulrfK0OYqLdA2yD1Kx3LHRddbRwuVcey5lblSe
RNX7jaYyasZThrSGur3ILkhFhUmHp7hhrP1Uz/YacLWq1X5gHBm+B9jlQuxTUue9
UUH0Vrl8hr0omvjLVCJf9h3EWc5F6W/qu+pqMWjdc5JEsoXDCq1//kQBEQv8Ygs+
v1zc9KVgZZhtqogywBXnaJpq+hqIusZ+aAyHryspUnEAtWaHIHVCKdDhjx4fpSc2
DfrA6mrYdI7j6W01B2SWMFaVPklIzvY17MszfnspfdTFoQJeVFXVMrm2Ue+zttCH
gWumzbddHTJ+5XXSWfvTUV1fJDcwuiVrxLMWJtxsE3mLHzy2JBVOCtqe7B/wPguH
SOWL97yvOFKIVLM/YqeltL5g9MgTYB1jERQ8I9xEXAqUaJLh8ah9m5aZwf1ztMGN
1qxpiODIr7DMOUWIb7e+enCdl6EAqwOEmWSISP4R39aFCAhAv0sfs4ts53sDjQzw
gIHzOdhG5WSJUsLIIXNwBpouOVKKiCeLwodAorvvfOdf4w0cxP7BqvKm0VN3wgma
kaaVcDiP3zV92nIoKdC+Jg4tt7QctrZ9Fp+oRn9/wdR9Szaf59NnZ94/kK/VqHGr
sWfP2YSuLSHlWYx9rFQeuWJPsv35Wmbv22asV14tY970qY3Ps4hMmTjgcdvbc6Wv
UKAurfOGXQJN2pSe26lau0mb8/+vGhRfdMeXIzFKDdM=
`protect END_PROTECTED
