`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h+B7FsgnRY6e4cs5iOifpIz2gcsnCjz+FiU6qyngRmck1jkud3q0dEC3YmCZNSLd
dsOfc3zLFg9oFVmyqLb+gskFxZiDEgco49xaKT0I1s54YtHGeLLyjNnHUhb/xsYJ
xacqCg2e8PMIyKc4kmOQ3kPCaGkOVQPEM4856f3IWCwJgDg1DiaNV72bKlX1kjRx
1saurQ4n1PaH6ouOhuGK0aH3ay9pI10uCirRFKGcZ2PfK+ftopkSnikpWzCbUJJn
OxzJOtBrS1FeYpS6+fr8YVN22VFuFT/jiw2VBTG8oRWVlH5NRbw9r4aUSfuMJoib
VciqgtBzQzC2ki76Ji3wgyNKJ7CiuT2pBqgsn5GsbbJT4MV6CM83MSp1kMu9fFBa
o5V4v0cQYqsMEA5q+ioDA/Qg88KC7LOg1kkCq5ZTIYUWBD3vYgic7gizFvkoQZoi
biZb67iHtnPJEWoZzHSfyEnbiiKa56RhJJ8oNrdrzrnLAEvufueGGmPJugjuzGRN
YE1gV5VjAp6LgIWKNmmU1AFMO5TDN8Uizq/8gdKLE/5nyB9CeXX5ZpfjI2Ux0VWX
OZZ4OuTZiGuIwxQWD9hLE+q/h0yRGFsy9XSWFwIFAw3lKiQ35dmhBzZF+cglVgL6
KJyGkOQgppeZdLGuYXsGf38U0oPgvD/G0w0/HLMmWKonw1CQPYCdAdGdM2PrWprp
ptfxZF26oQIjwUpOc7otbJ6oAsK+W+ePrFPo9YOOxMoZaGENNgKS3v4tpMf55RPh
XulW7FePuoQFv/0RQG7L+jTU5AnKETkHZp/ofT70R4KVmTfAiwe7bsNV6UtomizY
PpiUEhBBS/EknLNQrtEFFItwU8dbDSIvzjhEGNSTkDNIOdaLDWmpCmL5GrnXLtxU
rULquPJ54JXNVBQ283M7Ml1U+ZwZjAjpbt2EhWBEUoRW7/SWaiEkEg8MWeNPeQdU
NSwJe+QCJ0tKd3chV3OZQWbVilHPd1xxM2paLcP/H2Q0nIyfw6r58SqEAQN17zKr
NdlTbFKHF6OFY9leF+/m9yUAk1Dnw/7CEeBjIwM6W/b0XW1kv/o0j9o7LucR5APH
zXtdK7EKi/BIcPLBJhw3MFGS1WWXC+dlUwj7y1QcqtHJQx4L6vaHy973edFewJ35
Fy5fJGSD+dA+Xod498qNA2C9POvGHguIuSDae4on9M1yJlyvLPDfISIPoQHpaAuf
1yHBKSFNoEKcH4JUtshpEm6FG+6liFxa//HwAWzMPTWki8K9NrwdcOeBAp3oI2iW
3L5vJ+x9KPGFEyjRVY7jw8nYuvACx8VtJaWZZmzUUokipBBHDqvMmNwi+D9dEWAr
4diPWXzQFJLQVvkeHFulD02Dl0BSfqc4B9/KOjr1BgoDsdAnge/AgGQvPmhEwcPq
yp+2YFiKbgVWQQI+a80bxCXT/YKDp0jGTSRbDyqNybfId8exzae4T3S2j3UFv1pW
ZrEzfI1ySL/8S7RllCDPZYZFiF3cmS+6f0B2gAWQkjGl19ZaAY0xVDNdqvpGve2+
Ixh6l1IeM1gUAu7XE6Ng7sDVE73jft0lu1sT4NcPwQ8CB7MpFhHSkfR2awVw2yS7
hnFqiEHB7e9z+mQ24h1aXuy8Li8VYL3Z/Zs/hD3dptI=
`protect END_PROTECTED
