`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JewpLXtfY5OdOjxn3/UsCvOgKc9s2X0pRcaooMinmGVHPzHsIm/tJgzov3bVYy6l
PK29wVB86T82QLyve6oBIKB5kFGmH+pp8b23KSvKwgdhJ61oka8hTV3RhHSXpZcc
5WGnZO8iv8gsqP+5x8yS3ZvKhW/X5vBSDPpMhuRzZOvMwa2Kne6DjWJyFnyptrtT
OGF+F/AXistl1s3It5tJ777ol/Q9s4UuLIBo0U3ETUxl1vZqcZzuxI5UvjKMSjjG
YNUbHDCvbkQpzsxY6fJiyRyf07DB5ye2In2JJWH0KLK47aBiI212DDv6SCB9cYcW
mwHoZmu/1t3+tVNl6Oijqw==
`protect END_PROTECTED
