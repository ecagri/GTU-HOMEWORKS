`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6o+VNaloghGhK1RAyPuukC6ffDJNEruOUOEN7bIoq10PxR7y0EYLcD2/BNjiV7gS
o83LxvpFcCVduNeI9XESMaWi1n6B1UTGWyq1sYuI4kb2eqgGLNUEw9Kq9d/GOmQq
RXE1ekbNsUYjoxg4WUEkCoWtxinjcIfAWq0m2SmkoKTDxXGnB97iqBSx2t4QtrRK
7RQQUAnWkUIabZ0qmB3dlHjsnhW9lLh7j0TCrCE4/Fq7OfQcxHZ74zMTbnMkruWs
fluYjsczbtg6ML+a/Kfyh0S924mN8qp5KSKtcfUb5yx4ZiDiEQ99FDFY9v9Z6Izn
MZ2OMU9jUwtFUdF9a0Vd13Xx1v+qoA4thPbC1gPl740XLGq/bDGD59uQVAL2HONW
1K8/xarSpX77A5YilBPH2v0mxCT01rYbj1uQEc3l6iggJ23T0+aXnP2/sm2KI5T1
j0ixPlmBPmlQ+tGizTvZVMu+tLmPk6spZMniZBORaEHyweb/UaBAyp1dIQauZG/h
uj53K49/AhVg82BQmooISaOlDu/3M4E/gxBA31agfxrvAGpxlab4LIVpwPnO/wqe
sGR9RrBIAjxqeIBisfCMYQkce5+p4+qPx58R6Cd9FmEBOTgTeIe622+sqasbsAx0
EL3YcBoT67wI3YywNqV7zUsJiJNJXpBEtAzietD/ONgFPr91HS9T0/Kuolyy3wkN
b7tL8hWsPOnQA1RQ84lsXWiTDxpRfowUQUK4MXbkaAwCB68yP7m1Dmq5uookDSS1
ZQqdED6SZ8wQszDt0WUZJA==
`protect END_PROTECTED
