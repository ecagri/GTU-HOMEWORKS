`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5nyboho+rUUofpNVmRXtAV47DSm2hapuGBEqaCKU+PkdiKW3Pl2TZJdfSD8dppBf
YgV0ZM56BtBXp4sZhW4ltQgWQDbGsYFqvWb7uDJmDBDcfzexrquhRn/hwDQ/WMMO
eur/b9J6UChyLUCfx11TPwEmMBM+twWajmwlIP4b4AOOVeAL+YruYonMvF7V8FdF
edzjnM0OMaIJiZfcvDfdLjuphoD6gqgty9nBcdEoPSTt7aP/41k622JYqOo06d2B
9ZRIAZ9Dtc6nMS+uOgg9YzFyWlNIFDqm6Ofw3N3DBRUclOSWUKYgA4qbVmAghdC/
tefhlILIS+W0prcaFVQ5Vr+2ysDsujE5ucF+Vk+D5qIwuG5Py3PgqEuSt0QVbY2a
6u8v80YqDVUmgu9Y8LrX+97i9v8VhWkUBJ0L2c1/5qrZUY5cuQLcsAGEDSh5PmeW
ag965ZNQXqezQsgKUIIrSWuK+h5A8fEpDsRun+xLjmNf/TAc9q34svtmmL+CTBvJ
0jJgDB59EeevA5UiNPN8RUxfI3/JJvWXTN+ZO485Fi0V6rRru6zppLbH2yyeYd45
MB608u2IzMMoXQfXyJ0p21nvdw0TyEBhSs/RM3Lffcg359BBmLEDvHTQui8bdzKJ
a0dxANcV7DVwRFrX+RbCPweTDIaNf7DGGl5dX6xvJaagymPlAfFJiZ6eVgxrrFp4
P7oviQSgf9AlYilP9PlXuzynVx0suymq6J7+NHZV1ECYxTnmJLTzd/9abQzx8xqP
/KB7FObFLmWfXEvacOd3VBYOREbdD77buJHiRsWqkfxKHFXOc1YmID2sEiLS+0pR
JGP2QvmaltarX2BuI9e7Tdswvw9mnM74s3LB0i39EwQqOQrFurLsYvRHIVKBUHY1
eQ7laWQz94T85bZatxzhzp3hIxruIWepiOD7wCKAvOcoFRYwEQxo3lIRJKcsas1z
iQHvWkiqTDwlbD/LLsfhvHbPPX6DbRg4HjHVNnhw4Rhc9xQS5K5fwsbda+Iz9GQ6
kLHJ3mO6Rjsscr9YzcjgLfXJw/Gf/K+OJLUFp07aVixeZ6mYZf9ghRysKNT2DxLB
Hf6nV+7uARgQzMxxUNVF5o5yCrRLU+665dO49Msaf8tLD1Qm7HqkKbwyLhNrClEe
nMfWFlyoP7GF0tJfMFR/FvpoZYMjFW9CUkfoRxlS4ipplO+XfbDsJVhND3ZmwXhR
tTjSw0bqWw4ywivPEtIomSEO+NMsKDJYY8lgXXdqSsktCHftJ25lts+SWPK5flHJ
lwi5dmrFN78d4b3nPUI6vg==
`protect END_PROTECTED
