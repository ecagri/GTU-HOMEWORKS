`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tfys7nQXbpe87syTtxixQHMIA5Gmn7X49MCNR8D8Kqx7Ozr5zY1SGW4kqbPaz5c+
Kh2JV8tHZAC4yuvuFrG9+fwNx8beTgCxYweMHhDcQN8dtnLJlEfugWafVJ01Bfm8
mR3ZPRzevrA2YmP8eSMk+8FZMKryiWTe3z4at+ssZGzc77vZSpicihIVrLlonNoT
63rY1kJgZu0GJGiYNnydjHO/dnUEg/BX2Au54b8HwbEKx7grR1zgGE74khyGLsYA
sfvvgtkpPtGKresSSEa+33Mm6Rx+J9EXYRRsxRhoDXmTnSsnKfGcffiQ6zTpjThp
NObVkRnsldYsiV/28lpwCvYarof5ctLeavrbdmU50NINAp2wYys73vpYRb0AHtx8
n0xMXK2Jg+Rcy3SIbEeEhUWy44rIAHI97eIJt2JX7uJV3Em5iyH2V+TiBIPH2VRa
pY6iS/AxDR+nAl3AOmIzYaE6NxwAQrk3jaZMBvuQUv9WsqdekW2Jq/Mi55dAxSnK
c8rkDAzUhoce8qwPSx635u7Z1tDRO5RTeoL4xaqJtxPW+cCqdZdLf+iGkG8jdUL1
rUV5qdkrrDV0ptFN8lfrtlfPLCpdCmgevPmE9N+IsnofcoIFJLwqitlxt2OqGjAy
L34J6ElInzYknM0ycA7rrRu70UF38txLhpHX+a+54PnLcG4gpB6Ma4wBEal0E1IV
z9UXy5O80RZ/PMFBHkJL6pjnE4N9jjgKYwh6BjYUZotemIeehqqBKd+u6ptKoOwc
/BLfzhnZq7xB2QIV//z7mwLg9sCcTZaEkHRBWi38FBDWgPMIlfiU8/nnkBfAzMLn
saYr23/V7rtCK0rGHmfgwkRkVe2w/pskEPyFaaGpwtq9KCdjpeJzlEgoP5rHvUNt
MunPNDdTQNvt5LBqHKimkmxMecoAeE0GrJ8Ghj6IBNfIq407ujHffBBKyB4hxlKA
u/0z2Nlrcx11GhDZ2KYciHLKG/d7om+7bWUkCHIOMVQHhZVqs3bGnlGMJbkqi7qM
Pum8Z5mX0bx16mKGllXx1MaLJ1+75jjN0bdEX2t7Qlt/hgDPnQoy4c1ptiNIMxhU
qc4GRog6iq9PUXzFwI1swOPGho3Tt1NssMOjSgDjsocKVnFgFMMwkAvhG3CDDOAI
kjJT2ChE1PgrTq6HZBdlxYgI/aLHtayuNkAn7F/YK37JzlPIegYP3EzBWnVDUdH3
6fQeqKls4SzvOqD5vESzIA==
`protect END_PROTECTED
