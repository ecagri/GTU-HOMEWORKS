`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3S6jIEY9gxQCJTkgUs7Os0o9TZzx7ePmI2b4j2ZlTd0ExPITnRlwBGj23S4KR4Un
Z0rsp3LOf/es/5FNwMh/dxlP8qO3b843JsIzbPOMPYnWcG+XSsBFqMWYqdISL1eP
bVUfdouDUbSV4bCWyXvCH0F9I7Ds87wm1CIiEE4zxuOhh/cfNTa2HzfCLKM85S/d
ybPwaPrfKhpQ/PxYCPoR2Vf892rzUHO5u4ehKQ4BAWFiH6cWtXGQxH/i4q2cG1XG
XLk9QirvgpCk89RXFRK9aQD9q/U3R2SKXtpv3W496so7SvPyfjRBZXQiwMoua06P
dVWRimnfxzYncqm0H7CclB2d0zBtva9QSbP9528C0dy9KSA9h/TqK9eKiB0BdOsS
bMpOs8Tu1IxnB/zUk7mpVxq/Nz3V7VXv2Cf3gTmrhsBCzf2Q6BG9yzg8SE0KJSWk
HkhztW0CGHj8cobzbY9XH6jx3o430C8VLhPfukig7ZwRpap6OanbY08ku+Rk3UnP
PxZUkCXInZK1bAnb3Mkxc3Ihw4rsy7ALSrmDNjE7ShKiXyJQ1Tm6kPDBUCalBlfy
NSJ1kiHdwW1c17KB5lhbWwmc7kpkKs2MuOIVWgA7EqzFGT9O+dD/gnUR+m5CmsyL
Yp8zSqSCEnnWe5gbxNwJTEvkDTosYvVeSVDSuhxK25NW9hWk232f57QTiyeDELiO
RVRiO9slHNKbEES/4OtMZMrFWQBZqD0R4TtyZ23R2ARYpPQSmwX2tCip58kV+ceD
kWDRdE/y+ZPUXfmVeO56osL28WRHtUih8Uuwn7tohOqhczWsOVgIrHeXH7AkL5Lo
YcNsZPkn6uRvmyJC9Nb8tLqW/5WmwMevqaQqxGWYS6nG4Hc4+c+5PgVfbIXCYHeU
oh5GEVkA0TBr6uAvmLg6Bt1IoWMet59Od95oqSuCG1h3oHwhdi0EMUOhXWz1pG+t
Vu/FR8T6LLgNlVF2mKoqPQ/A8hT4kO4YRiP7fZa0G/5o+9Wqbzk2vFimMd8ZBMyP
r2dKanioSI1f5bnZnCRAR2HaH7G/uHz/pbEuGg0VeKcHt6ViY6aDjdJLBrfAGQFQ
rDFgJ0EFl2SHAem0z+kY/54YZYtJ6zuTEQta2rVsvUIcwemlszuH0icuUPESPXBG
LQGDgkyhTBytd8MC5x8OPqaBN6yquxRUZePVeO8GTShJIBGkrKvbIwND0+iIpovG
3JjhY03gEohYRDN6bMgTe7dBKIeXyWb10f0r/GBfRbVWJ8r54DUNPNzjh9udzNB/
cX5FMTE0/8+Npw4C3mdoPYUXr13uKkuqAYXkJCvEBmcu+5LXZxHwHCc//Y8GDYXy
flOjGg6dAI7m832bk1tt7gRHOcLsBVzkvPWZfMTla0sISNK6e8TZktYlWteZCADd
yQYm0iNx+Zr9+sjE/mMYBL5poQaQsATxu+YFdEjGe/sXzXuzThKL6/MG8pM3yuJ6
wUsviLgo2HN8FZaIcMJDAyciJyTxNk+ZTipDfS5l0LtKsNJmbfNEHWfr+0rXscsh
oU2jHn/Q9A/CV3nXlOnkKg==
`protect END_PROTECTED
