`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oGty+qA4DvgX8XhhwKhPHuSrYfj6H/3+I5yz2rER4W2a3jSo3RFPzORiMDlkiu5p
uEej0daKJETgCgLsQ7nI2SbmyfCZ2p/sX7ReCe3E3eiBGFDWZl+FZfXGfVazqStO
xIF2A7zJO/pHCWkarTtvOuuHB+jcfr7sGd5XpAvRXEPUDi40yLgIe/hrAcEXSy7S
txsFeSwWjn8pYN6qe5lZX/lT4fVZrImqAEu7UAQcgqiI3nyUFDiQ73ffoeaYYH1O
6Ieb9ilwgTH0eVg8gYtMrMgAApGvheEIxMiIV83xG3ZSR3+h+49083lgwNZW5a0G
KrAmfrOYEeduq6RySxvsr0tiksKbFVAZ1ZUk/v+SPHDmKTjV2WhpIOQoB9+HSebQ
MGAmS/mSqkgjb43B8ExUEiAN9huRNVukuQYBVqktYkRQc0GhYiDAKWz/W94P3d5A
UtyWoL0fTjjtNJi0uu7jK7cunbYno5477A2+dQARmRubhKy5he4+4ur5T8E/pq8a
XWfJuH6VnJWRSAE/XvVvZQbWh49dc1WjFLRqp0nT07Z/mmVUoplBW+o7I5qe5Ma0
x4g15kw7bcDOUOX7t+HjePmYmLnC92wqiJ0+gtqKt/LedOR5oYS4aYw9lKZujeY5
qaNn1qLtLtWIa+6JsWtNBjvCD4zvL3RAwvk31PApkpXVd4F7XWIOchKXJBAgnWaa
8KVrgpSSLBg6ISRJ/bLCsojTI951yEyfVO3sojxo3j79SD9ZG8eVTqa9VYqZG/1o
k/xXzItM1pNgeBvXx1QGe3tMRzcUbYGNSoUrJtcWG7QFJefmbuufA76xKGWWGMFL
upb9JwrZFzJ7JMi6FtszVrf6aHTiQoq9NuwL/yhajubQva4n6nmxmEojYTIY6K+b
8LEfs3DUxTryydpaQ/uET8VNjuUIda2ngee7314aCzJ9q7J/yWA9hjwDqVAQRIFk
HwXmCAJ3k7HcC4E6YNb3wQw0/tdXSJhh3QC7S22mhoAYo0nyTAIN3YUbVjgufZp9
pK+GmWM/N4cWJZn/VaRQCiWJD2oNUtuu9YPh6Ao3A8h37GkJuBRepR7OoWpi9zhB
2elR+1h0m/G6gUtpNH4VXtCq5J5XxBV0Pzv5nAZIKs5V5HuGCSvZoP1bpmu/J6gM
jP/6yiD81oOdyhXGwpz4hbQjEsNiFI5jLcOZe4Q8KF1Y5fTmKg63YLXChf4PNw8X
X0KEZPVGMNHFH6vcg0CVcsyGk42WG1h1rp2+SdpOSX7fPn7WUt8jbtE3ahUqDMBs
1y4BbK1TUF0aA8lZOFc7wDUdIxxcY00s4TU5AuA+EqKQUcFUsp7qZNIuUFGfmmWU
alRr9hzPWQiY/lHre2pi+ibBgC4obbPEVGGWgvrTpZQ2nKccu7CwYEqolkfeoR6n
DC3WzuQBtoSJC2xaHR4lh18QUsmR3uD2V4BC332RWEoV71aAXBr6SP2wwK6TMQx2
W8Gnr1mFdgtO86g8Mu96TXKlaLWRATdwLIu0QAwh+Y/cxRMozPIV3TSxHIp1W+nH
S9IzLkIB1uOBl/3hgruVybzGLfNTA9vEvA9I9FUiAnw/ton28uLAJ70GUwrdCVM7
iBQiFYYhoTS6R+rGqGlY1YnJBbSDDhvCja70Ep6GUBiG37aqwtQxyDnD1qx95nOl
bRx6T9PW7bPQD0O11sZIjiH5YREndyfRyDhyf5U16Wls5rmktLaJfkoQHIwmgH4n
9tcin8WLUl4YKvFShgRgVO6XyvXsnqVO22axk2yRX3BVUBjiqo4s1OPenVlAgmGd
OuBXfBRTE+WELMYScalpWxA34itZNIGecfzzhqEvlR9Wi3X2DovUdEtU0mBXH2SW
3/C/GcuqeZ0WYENFYSJSs26XKeJ1v0oj6kzC83kPnhhmIKiCYhFONjb4yn/XDQH/
SBjTbeeWrYXgxHYe6pFEMdMrHlKVhotLcYE7GKVnbt9A0o6g3QelOni7dbD5bzW+
rk9TSC1ZNh3/JO3Xf1hHfEoFk3HeTytoU6vXj5/ITrwX6EgNPQISzxWX2eBJt1Ug
AzP5gP6bCLro4jZ3LVjVZo4lX0b/8sBL7Om98jtmKB97nZWIByF4B6A7bUbr459X
+emewOavM6cRfwXnWIIBz/zu2qzc6Xkka/7hd4YWHm2gM2rJ6cT+sOTD7i+RINoh
0z9sd9XMzgMV1Ty0Bd+Rt/eH0uRmxUblc6/01ThFWCeTE6WGF2ONwIHAxZGyosF1
WuJHPmMtE7H+rlAdkDTc/KG3P19iTB6wwmf5pnOXuNtaTwtAfzTuVuNA/gDqEGzK
dbXCXNV+2NE2DeHk1pu1Pk/Q4aQ6Ar/cQ+tlBfU4CAOzXNbwL+REjX1CsdfJQSCi
9IobcW7+cIzmvKropImxXgRJf/ccsTYenUriR4AaSL+jvQyXVnezi4QTCUCKfYUM
SUPwIPXElZ6t3NdudAemZ+WSRx4osG4js/x7iRPbCofxhD2tbG0ESxNj5/5Vk77q
CJEZCywWFv7egd8sZji4cihp2U7N4KfTb1qdlhZMLtLqiI/nvkR8VrEFYiZ6JiMi
n/8f60eRvXhW3FENh8zOf1MCGYDytpAcKfBt6p3eY0DDlEioQed/gmXrlVKfZvMH
am22RoHvL8LC+E2H8CVknTj4PucPGJlDid3NiuvFp2RSICHM4UH1Y4olr8oUlcNI
p3uu2QKrHYluyiNdDEoBjoc7M96KWhk8vDqLtwpDV+fdJGErekVW2atGuAcmoexr
RF61299G63KVweOv3ytma4N1PlUB0mfBI2osQjCETtqS7YJMaLSpO61RPjBNYtIp
JQYDbBHQJklxA7XuV9h8WSiB1XRDQvt0BBul00E+bE14rYJZpiqPOkV6AZ5Obl4K
bnodxQyAJ7TJCahWnuTW/81b0jXcDhcekZl3FCx6rObDrJXRV9SzHEmoirCxpakc
8iUD4yXCycS3L0edeu2gNlWy+SJRxTGvx7+L+2iX60Ulu9WKYdWSpeUs6urXWAbY
XiinPi4hhgCdAUAKfS3FEo62CfqISgFRMMBy8uZ3QhG9x1YgCh7jOdI6GxCe5wtl
msZ3cyeHYXYOJ2so/D5XWuLTj0FqUhKMxf5+xkQru28k49Ac3VWGXHgYGOvOr72m
aWwmcqcpAbe0J4avhCcWF/U8brUf+fBsUhTF66IWF1nl+WdLLgLEIcRgjMQquOHg
Hz81mXQg1NVE3a4FuyKxrnnhIAYIBt/mxe0AfqGtBtdBfwcgFZkIEB0d0FErYUmC
FaJ0CXW1B1aWVQPi6xqoxmgj/hwbkyA5AcIPSdOkMfwLZlKNpcfw+ZXW7a+ppFEO
EcAQDElu96VVWYTt4eRYuqxOJoVm7ch2aDVW0f2PYjxng0Dywbs1qhGDEs2Q7P60
eTT8f54lm3M6eDxgniI31ejXxefGMif57RdsYoCv+lhCKD+2scoJSBJq81pNbeVp
xAiPHXSdbljV8MrZ3BgX186X1Hrc1Zp8k2oshIgAD4R9SSC9FBjPhRx/BL++s53C
PRBJciI9eBKmi/24VZ8OWyl4FNfS5kIPSxpn8hAlKBqDJHVCGdRpKZVKzG1LYOq8
yxgw2eQc1KuOq/oHYRR6JhFUTOitPUjvZLSS2kaRYYM6+uV0K2C1jbEZ6xLifn9v
R8L2Db1XgdprhsGqHtCsA1Sxvk6eF2zumHAACHazy9bLiYbx8j1K75ouLbqtiMVu
jwXwm26OP4xSAt6X5Fgko+N/ArYLcGsgMPUi2IDlqU0LCoAwfc06/vnZzh4zCO9n
mYRxvF6nfULparimfhL03nrwRT2Jn4iFc6/Ef5ydlj+5J+SaZCXrpjXBdQNI1m7m
eNwAQnC77kvlOl1fJLI/pgaaWw04Avl43ic0fslqBVT+fyRmm+sZjxy9HwHO0f3o
3HFqwU81yhVwK2oTLRxTu4vmBsH6YPJJy6WoWBNYCqUfN1avTH12sRtNGE84Fy8I
MZfSlO66RHZk0V2bbSYaT6uPZhEFsZ9V43qzZzHMdXqHm166WalxOQPJUzy29IuF
zidIWaPOfSq+e3KiecIAJuP79rzM+mYgNKRFihmwTfjZNTBEa91rLLq45EJOl+zd
lWbhpHoPca06eB+ERLAmc66w6Aw7LvLREUeNXgEJrdtwnpEnypQA9euvoB6NbmzM
Xa03ef1IJ+PezhlLrIv5Y0hlTXx+OzyKIoOFoULYW6PubaMymHu6NZ54+70jy6GD
`protect END_PROTECTED
