`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lqrBsIk7vSgUx+2f65KUwJJMm7xQ+OYJHLyHHZz9tZ/5lG1F1SCy95FNqqDlFQpI
lNKtqP60OzicopXXwWWv5RSPnvr5c68QfpUSLcKuTeevrcjU8Q8YktI7TqCW6k8X
kVIXYEXGi69y+cQ25Wafs1ZnNNo0Tc90El9llY5+PWbpMyzZksCIPXrFQfDeCS6c
2Q71gk+s6j1l4DcblX7B5Ff7udarpbijRoU52X8uCPn6f9pQA4uvjCntrWqUKSGd
D4Hw91bcci0SZjQFJvvu+s0r+Ze8FymSt29d9vmgDRNK8P1suiimatVOD3Y9cT9C
c/Bw4mproNEJ9AIX6byH4nWFoqIiTSdvNaxMg77TndgH/pQRtUQOjBZfCqU82u1u
Y9dgdn7Xg0Cx/8oUBcWse4anY3TJOFL3g5DXwXKKyeZQR/tehquv+2ZwV/SxYYer
PWwNmTlaycNfXArQ6IqsrOn6L8oIOvp26ObjEy20EECuZlu+YCU2cLjRBQ0IXt7E
++ciE6ZcsAQgxy5gVI+/VyTUzdagMgrYmSAAgXOCO7efFjenrQKHkTEXA/uw2Uup
eDOzgf8IpKM3k2dryzdVCUopQguisByBZPTrZDd7takdTAoWDypdJNRsHj99wVgG
COqFF7lW0teRGWxWJHdQDw==
`protect END_PROTECTED
