`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
heZjTEu2TPGDA/8oT9qvsuKU6LsT6xZKHrleGzY0phb+pm+hYnBDKjHpj4TPe7VO
sGH+MI7QtmVxfVOXakITGz1LSFtgHGpebeEaxxakex1Bh7lOFdwrbZbXspDsJhcK
xFBEn0r1ahaujx7cTgZENX7C9vJyEHn6bX3vbvbYuGm40SeRq+GSRsppIj//1T1J
gQuAoUNqkXaa+HxG87vWNXACrSlUzsCZ76EpMc5P1WMhqiAL7otVrVN3kpZlHzy2
pDMVO/em5m8qaP75ftbytFKtgaxl1DCO6KGM5i0v+Afeo4+0LtAdCB2gcQEgUrYN
/ZL9NNsFpOTWy5FZYkHO+W6dIRWAHZMoJbxy3rdF9RiA37LJsSE0P/VfyrwXQ2X7
UTSTzFcqqJQC1HdcEfLMdstdp+p2pEIaDOoXfFgkC05O+Xl3TCexSoRsh0pFNzKv
nX6CYY8PSJ/CBy+8d/k6/sDgNW5ZxCnSdG9UKT3TbU0vW7Xg8Mdr4pcpbTfjAy1o
qn/UTrFR/ASGu654BZsK9JOVTNjBHFPN08F0XP5t1tqPMlk+c2gYs7FPzv4U1mfJ
i+y5P8167mKEe0XUuNdnontKBINv6E43Nh2ZbzFDaoEWB1ExjbaveVHeTf1ARHqS
GL8zC4uYa06pF1yFO565luN81noDOdYjNTv58VS056F9pja9VfthdfIrc4y/BvMN
le7ITyWlWpeBwC8SvKgqWI1LQy3Q4Be298jEnf3z/avitNgu6zxKr9Z7/Uu5ixv7
A081Zawov1n5i9cNqqNItCPgx9P93D3QN81ZgU2vctp+bmEfMviX824upGAGcyol
DjhvcvXzfm+8aV1MZVr4WdNPnco+f7Z4vk1PwhE/R9RNlV1AcfjLRn7YHEOjP9aW
muM5OyC+zcFCbWEWFS9mqMzIWzubzhQfsp4Q+uhc1qfZIRxWK/2Ov+TBG77nNAmb
kaR1++0kOoramcPUCcj+lSI/0VfioBl8kz/1qGA9hX1ciLdmCckZ+6DlybuMQZdH
ca5RIeKQ12gz3AdlKURDTE5LHjzqRvz5HS+JGgwxFtqHbWbzQQsBW7F2usni59Ol
b4FN/Pcf9NlQ7tOT0y2y+R+xqoQKaM2fW/XftsGNiGrhcb+cGlZoZcR8h+aZvqb5
ho7Ojb7dOm4T1Pz9MCK1I2iz5rVyjvrOji5YY5mn2S/KCikOxgL1aeZh6makX9jf
6bUxgcnSFHr6/dSaNorEayvXODZq8U2Hg+BplEniAsatt56QJTNhZ0O4Pz2CpZyv
NT9KYx7tYyMvNd04GvWesTDVJxHhVXddGrlSujqIqzS668lhjxh4JfiyZUvT/0ni
XzO7UhS0Vq2gZmeQyQjiiY2V+ZsbMi4kmMuDxibhgWsHi81h8fBSQm+CQU6G2Ocn
grQmO6flYRePaRtQDHw6bazKrt07h/6F5VUzZr6dF2xtj5Sy9NKxvkRHqMoqlj3V
DjWrwmfWTlyP6J92Ftu44DnM3OmyXWpwTUuX1n2phz9eQhLbLa7dhRVe/BhaHGRj
ny5UanZQjEZ4NsA1cjRDKRSYRK43J0atVCyptZWAifGoF2Z4xm08HiwUu9eARlsO
luyti0eA0INntM1INwT/YzQwsnvygkIn11erKsxHOPXvt/wEn3SQ/uu+ffmaalzt
hw+qIjW8sK/CQkj+Jhs9uw==
`protect END_PROTECTED
