`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YFV3pIfH7CFexltf4UYXDBAEaEq5PPMVenAVjVPLVU+mdUcLXuTExFxgb4OMvWap
vhTXfKXFUenlT31BJyzjb03+npqLmwaFiKyifrP0OA7mvF1c5H+PQRvk5XJS6aMW
NujSaurcxjLUhNIP5RLHlmMDEDbIGDh3ZNRrEA0Dx+sDKdSZYSs0wbMGJihfCcre
+bfmwpSNWQ4pvm6rPMfXSFiHR7WYJpC4axL2KRVaLxGFRxyVI1mUBRFt1juvrEps
9ro72notQ99/OMjvLrIQLYLgTQ1oq84gjuU83iwUN+GaSExL+aRqQSvPRrVB82Pw
41F/6GCWlCQnj+K9L8zkp35lQAxG0XqGWFGjUFfG3Qk8E1wpOHcNmG7SRwC4FPit
`protect END_PROTECTED
