`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z9e1yZbJQzNR4slfwNE+/l40epAAD0S/FKeBAQMihJZLs/byQQ2RdImx2diESOnI
CvNqMQ81ulFSpHKySsIrbFxNjBWhhJnPm1A5kZvjiekLUgYhd+Hbn2QjhdeNrRKm
vnO13RUjTLOpV76OQ9eiJbbtAABcWzbeKC4tFhUwy4mUiNpJlMt9yi5vLFQ7zu8Z
EOrrdHlkdOMfT7PPE0i6MNSoYPY0B86SNo9gzNmD0A7TZnG+XDpZ6UAldMsJTBQ5
BkBo6JrBPkQ84KgUcEBEG+0vM9cNwINivcM+eZgyNm8IsHsZDuRnYAfgwCdrteqT
4fgDb3h+2Tk3irIxNW5HxzPPsGheLZMw1wHmB+CuA6IlJNFKOTypCNXjPXzBNcJp
COUzxKyzu25R1OphkuFnK+TlW0DDOepIA2tguRE4ENzyrXEaJBz/uHmpOJO7Jcmu
dVXGRBcBqrHB22MesH8EZFwhftJr9KH4WOkyyJy7TE438rARJhDiyMxiBOnk9435
fbleq+QhXznLgtcWtfFWFiLMiVUiQoH2g6rDmZvspW/z7xeEkQ8RHAPJFZjmmaOH
W6idZKdQKIPNbtHYk79qbKfQ+TjWxkvgOByo0SwgpQwpa6cBAKAmTsyziQIXPZdG
SW9bdL1s+qnA1HSLMBpuaUsgEe61SxZ924F8d21s93rCbNvQeqI0p1DWmx5dfPV1
oPmX5MpAbPndof7vgnpcs6c5ffIGi3OHTjbfPhEz3tzeeqkI9sWqjyZl65SrYMRw
vOxwXrNBjPWQDVeVjGPYsX7JuRR+y07h3a3DL3u0hN5Xb2SDehrI3s9rEFwfiNLF
zuEsNM0xUS3RmX2Krvov7QLQFWLFVhFsC0iNY7LxXwYOuXNLDitf4az6va2yzwir
VpGtOCV8XnytBIl4BUJZBcyeOsj2gXer4O0DWo1uUzYje99GI0ONT3WnbKedu9e6
v64gGHjnSJ+FMDENDDgkpEsqVnFUIJIKZZkHVmutvbR0M0YEAU8tY9VQw6MJMcRv
uav0X389zHkRNNxosWkTbS57Taxbu/4HYtFTt9a1h6e9PcJwc1oH3WzHsDrDsbHf
PBOSIXgIkPly825RaUifeV5ixrbuP210i1al5v39wp/EpZfeNzaX9BWS4IriEpEi
ihJh79QZBXbAyH58FVQuuud9G5YuI0C3ugVdx+CaK5c2BFBv5XnMEKEIoPA0Fwx6
g1f7cJmT7zrtOnjMN735URdaxQEWAMP6F/QnZhkDXrxzzKS3wtsFV+NmJrCiufob
T/r7ryilTZ/tYLMHw8EoDdBodeGcdY0y8tWHYyF9z2RIYihigYqcdD9TCeBdlAIt
N7+LxKQsIreqrPxaCh67LvkG1N2IxTM1JMhn5jwa4+2kAYFS/TV7Y6UhV5mYQth6
exebgvGWOH20k2kIGnsrK+/NtjbY9iIXb4Yel5EcQOFxGFcBjwqfR2fIjZAl131z
5sYt4Ef8iD618SVYGTn4qUUUnSX1CDrZqGt1X9rQJxVdIdU7CZ8DSSEV9eb6+fBE
t1G6eeCL28JPKOImDEHoqST3nuTaljkenjpm6ivGATcFVhbUvccZgFtytXkL8b6e
rQri4gyzsmS5vPu9KurIf03O8yZMS7So+fTbGp4mq8fdYIbaAq+D0HeBeXPo+F+O
l/0+dHACPnGd2Zjgu+BqVk52YgvgSrFluexjkAatFUCPZnE7+87hOm1kJ//T5Mhr
8PGf5BwGBpWmwrbO/Kir05XYojfR0uQoqTDdqaN1OJZzi3vtcZmjQUHWM0UCu6IG
gj98zGwiZXbzx0KcO9jLejrB6HnAL0j1AYjGBHw4TMWtrywZyeiedXu3FJbmi9TE
aN+bWmj1p0dro4+8clhur7+0Cvjnuyqf7qALxZAT5BljNxMj7slrGroaYeX94xq4
iqep1hA16XFF8lOy6/l+FqqD1HmekV1UYcwwsJoMQbMmMq78x0Wa2QqooBac+wLn
6l4OhSDEV6JZ+Uldgecu6w2X4rg8dx2yRzYajHGq2js1C3oJRkaJwygq4DPlHiZJ
gsErilpcoHleRo5TWqMHfoDNmKyCcsrMTTlue4VScpAKyM4RTSPM3WY0r35hS6vU
3iWzrPEEpc+ifs0PE9iD4XY/vHUc6QllBtrqN4H0FF8w1T5jCHD9l8JzizMVX6zw
HYq6PZq9CyW2ZYgAJFUFk6LpB38n3hUUVg+dieV4WSW2xSksx2kQzX2GEnP2MS4Q
8gYv76TblpJtm77cthZ36NNMSbN7ge/Io5Hd6aeKWfg2A1PC1xKzWl2pW+tZNKPA
KerZgmwGl3Q6s4VbbBBk/m2blFzhHDjSVasAWSvJkADYker3CsX7TGUHeNyu0Up1
lDZnarGteTGu3IdL7KlIeDdsigvXoeLTj8wDJF43QWZ3n9XA9xt6eyyIkEl0NXiK
cXMXM1MhVgN1JK2AcBZJwMVX1Iga76m5Rpjomx3xwwpdAY4awlRgtT8qQiBjvIas
HSjcB5K75feOQr6A6KVXYkzTibc1wM7oWY3FfPDhUZYK7Koq1KDThkqS3Zf1qjwD
dkvdCi1EQ44fuZVnqhneqXpU/tqIx1EntC30DA2v1NviZ03naXtXlT5v9Xty7YBd
xhkzynGH2TwmLsVDknfi+Y++t/UGo5jn0Rb8dJtJJ3qhT3TEc380Md05q4/+oJLF
+VsCsyiVUKac9nU8A7BvGX7IN6INFvKu4Rk4DgWWLj/5mqMJBGkE+wMnba/tWXDG
zk8B3mmihqWQHbIJnfxdFWcs16fBgI3euCTWwnFHSfOSoo4j9BLJLkRVLwLvYh/G
wPq0f34O3GomUJA6hJbuxqxDCwrs+HRMjolhsZ7tDHa04GCMTiNpAFDafkwjMmns
fRObrPUIGe3TZzHjv9Xq+bVXrlA7+OI380mNMj5T1G521XZ+s0PsBwgDGqUHGq2L
ldnaTmklCTI0FhNMXf0aVltKrcakAI6qUazTjaLulT67iYZYbADaWkwxzWs2qQ7q
Gz4GjNVclVy+i953UCcTjrvfeK6wR170kTIjEWlsfb0r/eAEQ+gKCdSKDaJ68mCy
M8bhFPsTDLzRbzbTYbTXI5Zr7LxCZqCWBDkEYERWBCp+yAuHLD977tYia5Y2GnU7
VOi5bXSZlb0WBTd56CHXv+jKs0zGEmekAqkniMuxpAixNxMI4ojRwByb/ShnylT7
Ru53yV2qIj7XtuLGqVhPvKERgX15xRsxufLtZWyW4p3d6HyAwVN1g+8JAdjU/j1Y
DnicBDtgml7bE8NnDFHX+g==
`protect END_PROTECTED
