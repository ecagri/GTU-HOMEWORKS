`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6tbs6tJlB2KX6GkxPlDTQ/LP4mTTEPOBphg1oc2d4lvhA/uYnOGJBp5eOeHeuVBJ
dfIhUbRMWKEV8QAoTiXsdZ3HUCjt+zFc6gQDhiuDIY9wVhwn3+yMbfhZS/M8HCsn
JNAsakQqsvtofOJ2SdVdX8GiTIThMWJjzqlvr+tTCqMpCXINTavWTUEPh0toDgSM
KSW83auyU+HJjsTy8Z1rRJYKTlZ/k0tWamSVIuegoqSR7TcTh3N79W09+sYhetvL
zNsVB0U6jQ956haX2PoaZx/Ln8vV+MNA086rQP5JUiHKzcjakcK6VITyAsfCw4wW
/hKt8bW2ivq3n4H+ZMxgd/N9kMwssisi7dcGlzkaFrQ7YKoP/v9pK4olbhdUxLoc
kQXh4cPPgQhgHERvdHVPFFJWkp8KSCWMs2h0Ub6kVN+BPV+2TLNDaVVyJCh/nYf1
MHfbOhwuaclHTOA6ZDXJBA9oJvL5vlXurB7FsZX+TrD1vLTATVnQcy+9nx3iwO3q
yyMWdpvBROkgFWyQib1KaUCZEXyqGG06ewrvO0tyN0aBeQJuHIR2jWidbN0nPWR0
6wr0sW9U1dM0XCEtIYUIwGc1by1k936kjgKYCjznkccwgMufHpQgjTbCUXu0QNQ2
uzq4HB4o6YIq7Brmm0dGghV197xTmc2UOP5jVxY6dt7wTFp3wUi4TnhhfpeY9MGv
+g+9N18RVIRzOWjaRQxLap7pru1eHJ2RpibjULnaklF06T9ipIkdpaDlu7iMkhzL
Clh1m1C0MhfkTCGQuHlGpb380TucN+kJixmX5htwnmnGiE1l3H7mKJndK0/QUobf
KD7jhUhlw6jdBNNEtwRDiJH/UhwKqkfB+iAFEh9Es3ZMiuAKOFxdCgq/SRHlEknx
dO7SPHO0wlvOZBfcMhcLTsMNGWFaZnTyvdY/tb+F/Vy/x79FiJew78Y2SjHTDmsf
NnTtxnhxPwVACwcj+pmer1Tl6nrK6L31z0BXHfsVBDe2csAA/KUe9LsvRihfbkqm
15A89LYLczhRlDeB+gl5uBZZpGCM/dy/UVoGx8B9AWnW8F6d5qRQhWkGksFcx+Kg
mMwtK3FAE945b7JK/EoEF85ZSWhoPD+AJ/0Nn37UB4m1BkvJBYssGdn/DzdkVSzS
by6zSyFsnugxcn6aTnNnPEvPET9ouNUEtOGIpYiX94sTsH5vxLPwu1EAihQbZ5ap
nzEB30o/DmY0c45r6tNWg890rNn/p8XocgA7BnN/2KUCOcBnsONthJOL9RVueiDS
f9UlBda2TXiPf9EFQHIm78vtc78X8PQuqnWi3jCehh7MxMaa2fI9xPh1oAYIePN8
uqdNr0Yl+TSRADfFuqSrL4vX08caTrtBE3JwSvt0117PgO1AATTCDYVrUIUrFPo1
KDxVtjJv2+JoiGRsjLy1Xf/0CzwqafiQ1WbKlXUeLQnYwG0BbwOdhLG4gRffoVom
p19bnT8KQHgDkVpL6Cst9ZE4CPVvBklMJtvLl5G7RsiQpp3MeF+e9xQNpYlao8yH
HGNDP1/mHnT5Y5+m5MlPYa2Q2rnOnMFbukzVL+BIq5huMx2lMrNGpB0doHMTwVsH
ySnsc63kpM71Ww5rQILd+SpKJ1dqKn2P+jhwsilsSq85e4etv9gzqZL9Eqk2U9kl
b5UIhW6AHE1mCl1vAT2mEjFPV9nh4bqLwnnEzNwuHeM7CktQ4cccNQ5flbEmvyXC
nHaa0k8FFSnJG3KXaWmrZZVQRD05A5cXefE6+8HdmSOalAxRkbUIniLlDl4Ox1d6
d6h5mc7bpLayd7UBO/fMSssH4J9zFbq/AyfxNRox9yTF3G9vSgOEelkgEu69rcn1
WAaBi3wpkOPqLAcNwbKAKHp26v/mRSdMF2uyK3WPuvW1AsyF/jI8nYFwewSmwDEW
fW/rvpD010ezbmfTlW4CeAskD8I7yb+ALtcZgEzWOCC/+ZJtifXc92JCxNn7dGct
L1g9J5KDjD9PtAvYZ8L5PANksCwgYvbgQ5eJBzdAk+/S5qe4KH4I6KpeWHOpwQCA
QqkGSZfgbeVj4LBn9GBZK8GfwAzF9eOtI8PY5wke6jnFYZOjC+xdH1P2xWCNv7Gf
a0Bpl6bztlbj3iZ0VzV4dzh1NtrMTYUGI3Vu2Ql6wZ2h+klyN5hLGwNc3e1H/MxB
FmgoRB9V/cmyIb7Af6xlTM2MWoDojZaXzmve9pBWPPZFuIR+yVUHKKEYjySPUKNg
y2JjVU1FFToYfVh9ekKzUQJ4xh9ow2/6w2JZ9PZIqaGf2DE6T1Q2ydKQrbZB6CiD
0MvHEaLgsJKYOfgM+mgYlzBWAF/mLlq9jDAZ69w5K4oAWHN+imlM6Yomwi6autoH
28NtAOjwXUkhrRrCZuCNeWK9Xr6eFpbf3mC25xjGIlvVvghpg8KiiNg6VTQV4zdJ
cczoJEwxF3dnyd+8Le2FoW21aWkrVPEL+r6Jz5X2bKdzRSkLfNdBCAOjmkbucXee
YzdHA17YNIIbrYtM7mh9vHrja/x5ZYlDDnG/wOKCHQp5BFO078VVplHHaCYELR5F
qyBewFXNiQpgm32j45JE1QxpV7SBikYNDGbFgrNwtM/fekCLCdhbj7dHG/xr604L
x2+V3V0dYzie5zY5WFdx2IDZudzV6LvIzRqFtGzThG4f8Vp+J+t4NJ9WPnhCP/gG
rit/m32liP4jgLEs7zLrRDoX0ptfVaHiXJLZVEZ0wP8kNJJv75m/nOYr33x8AFOq
0zKzgCw+0hvw6c7QOCDTnPuK/JMWepBmdkbtGTTSeHl3ZG9g6I3R20gJcRd8bn8+
NJMkEBhGwaNH2JQthnTAK6QTqYfgjy7ziO3lke286ytfbeIyTF617tzPvfUAlyau
6w9wWuA9MrdVimuxT9b/A17fGiMrrBGC2aLKSPRGlqoJfdzQ7Ookjz/Tn0PwFhc/
VYMLMA/EhTM204pmB24M8sDv6wMzv73Fl+CfrqpuPmTqADNV/3XqG0KtC/X5zBPB
mbTIFZcpGqA7tIktrwVxLyqg5DVpsUYwpzA+yXp59Ni2j1R2jjjpHkI+7sHVfs6U
hU24XI69UspF7lXaziFoylclX6gHL+dkDPhhuske//w4utbMlKQai4e+8EnczTL1
IcrkG3de1O0k6XD8oAw3LyPlobKc21RLYuFslgBsyjW/2fcQRozSRoCuxLIwxwkr
Y6XZvaZ5/MulApuEcpBZENsAXELVWdXxVmek8tC2RMM09Eu8lOiIJORKPBIW1OAF
iykstNG+P/w4ZFkunD4m+I83B0G3PtuzfTq/4KsDGegpEFeJp8GRYPRdQU8NA5xU
osJw0VP/HVAnAt7soB9WiBDQzpnqKepDPkBNiPDaFvrKl4YoapjIS/5eLLchKKiA
825/8MiqiPUmHTiBuxNFlUg3s/WfphdsrawnC8aeBF+wd88H/u5mppQ2ihcwv3PF
gYF10Su0+xB0e1JgXZqvsfB1fhi6qWm65EOOW+N/eKuVtQ9d7aa1Rl2RKkIrWXH0
xkicD+TWc3c1E0jpuh3Xhcwv4+KzmSgkielKf9Ow+UIHFWoQkBsgXYUnMSTfpDDP
whjxjmEI06xGcSjyZ6ZH/88+fUsJAE5SZQZkqJviI7+rSuhLY/rz9eqy08VpTXKf
Not9M+O1ehsK6mJjh3BQs0bIegVDwrpGDkMnArYlGZqTKZKBeq1hHdIYq/wTJHm7
WPVNqGuvyRbDEtIPgnYKWNcj8Z2JPRhFMAQAMkdipY/2DIIGR94R6Nxun5aeXUix
PyYwhi6JV2pIKHma/LANOAk7wWlubPUShyvjxL7cVkqWuw1IX5IQFZqxOpxY3dOT
kYYTgYeIRKeUv92w5BSXRMZYF49BtZ9cYl/3RZbucx2jNCpi20+/VJfNSYRNCj1w
bw5ENUZK48+XHNkOs/uqi/5LL8zWFzbIoihUi/0X/cGT1z3w8zdmWdL364jEraOm
7d7hLCdoroIjP7LdcbLWBz/kvybeop+UU9sMIwnvDq1dDQKEQLRv6ViJZgnfl/xY
IoUYqbAWnMiXsQNljAJVqga4mrVo25hWiLq7Dc5cjVJfufwbfvLI/x+iVhNRNEAn
3BbGd/hOY5nPREdst0JrQ6hy/CUzuCe89TvagoRnVBZ8aUkuSpJFNwt81ZcEoVW5
bd/bSWt77pkeGraWbLxaD1o2FSfy5FRtzD0uOPXl4z/hc93vAI5ahpC/W2W2bEsF
NW6889+QE07DK95uG1Vnujw35zWZQQLfQColJ9tmRXC9Du2kJXHJ7TdoanPFlpsS
56VCaLJ/hpwRA2/tKeJ9LK0Dfd90etbrBoqgdwMjTJ57JZw3qofHfBsNzIkClZNU
ZpeTlTMF1ALyALi8dQEMq5E2dOfnh81vtPlfQKeqQFzpmdHD/7axhKD0wzASnLpA
XR3ZanXvoaxCUOwjsWsNtoLtEY83YRO8okyiO1YYiWeGGUs7ayQxcChbvCudkIkF
aZBfmAqwJ28X/mjfX5E1eXw7BipyGmhs5kOxdKXzTaUS9RMnY/pxBDASYdkZ2geg
3/gr96BZRWUD6BRjRCaiBabL0Y/WlcyGzgwpntJHNd2RFc3SAm9r0LTPopMkioio
wqJa5Wri+WDAq3qbMXEA6ANUvx9tBl3rbrciC6/10JY2nCQS5nv5FUzXd1tM3omf
OrCj5a8lBrxRDSF+ZfTAz5d9IU4/ws8AQhVEo2TtbSo5d/FiVTXp3BtL8MCJd4TD
UsQDJreZD/Cdf3zPmXVdYiCqr5+f8DKdTCEOyh6YPYj2iCMY23ajW1spxKX/LDa8
R80nvoTR3z7lgUf0jNowhScTxZN4HV2k/XJGfotPEvxKgbzNh/qJmj861lvA+0QQ
/zeLscGftgkQBtGcTziJhIvzSpd1DF2zfvfW3UJ5Jpnr4xHHy/hnUJd/Ift8VHJz
B3IgEBqKt2m/isBRPZCgMvA0k1aXRqJr2RLRWhDNVkmuhUmf1O5c4VFMFCszFk3K
CaT9MoZUm9OQolxREJHTvw8IxzNT4oYPkkB0mENIDbNyPtbNuVUXW3pun6wttogG
o8Fy6BKY0LNW1I1HvFpZMFEWv1RFGIBDVOtF/qp0Le7J2YSRwSQUGvT/qTFiodML
ceEpTodp5hf5AMyvfTcV40nM5F/giZYPxby8mOZdvS+FFkPzEtg+1cbN/eJE1ohm
T03jmzmqviRgTepfk9ay02A2KGe83fNeXuP6Q0vAaXH6JQqHf28QCrPtEfXrjIXq
GyMpZ++h964d4bsoMDYjD9EEBPwrkjbgrWgxMTCZaKky98nLDEqxYe+/RjC6Gq5O
UdOeg0c1OHrNvLVIGolVW549KGso6fZ9gyxnE6uK1qZx3SihXvT/BMXKaM3q/JxT
FDl4Q1DRLvrb+NLlcvJA7YkxE10VDEL3bn2POYJU2M2DDqvqSRGaxsC83N90D8LU
IM8BG1JnKZSe+wCap/LSlim77WB4IVfDXmYLW/DzhAbPvm/QBOBqekB/Hs2wQh1v
5U3/n8CUk9Vq0pXl5duNkCXzLuFFWzP1tPn3qGEaBrpUo1ZS1OMP6v5QAZMrBd0l
8CK4ZQNT/WnIBsJAgUL1HusuXHGD7oVJVnGXS2Xg1T6OL1rNdcjU4cCxJHDJizhz
w40Kd5xrKX05H390sMQdQYXW38qpQQ46fQ1WfIjAY++VuCT2+GAoqr8AKvrkpCks
9fUE03TKwDfSHriu1VUOrB4uDVI0HPrAMcRX3o2//sB+BJvnXtZEzP4c31Uv3j6H
xM0LfjxTTc2x90a5HLuuxso3UUqdc4JsL4zBERDOD5K5WXMgOc5F0dMkbESpSt6B
45V6fRNW7q2m1/QB7GEunAjOgIVeMTwgEphoMOS8iUKnGUWBA1fiWmS1aRpTnM+y
QqEnZW9g99xMEgDOKu7pNuZUuVu4Vf+jdVg/d4qa/940iQrpRxH+4ouRc2CR111N
NkQP766KX0++IDQbzAI6BM0m1WJ0b0ypl20fof96/PLnOaanuozhL09jR9T9bvKd
b+03DTAPgXgi+hL0p8hS2vE9r88UpazMzIlkcd4qzo9rzsgOTqP9Zs61rutLBQus
EMs3Cgn+u3H1VrLeE/J5i0mZfm6Tn+CZEWjo+1VLcOr0U7WfwS60XOxJ81irsrom
x61TbEC4IJjNuCrTRcbWDrxj7QlJo+B6aVj7y9xrwphu9sNwHdQYoKA1HA3TOeKv
YCFjKr44/D2MuUmRw4JQUE3fa4xATQ9qOvsDHa9vuu1H+wzEWAuLgeiOGl4sh6ul
268Cfwovf+q8S878FZ7nLll/sPtEpL3LjIzdVLpxP2YI8cskIe/6H6S8ynFeGL1u
WT+o1SYCKGKUpD/1Qpi3cAZDmCdXb2KwarXk4vBPSOzzkwH+B8puOkSaQRxmOhDa
xmxb389c1zIUg09yxaxZlWqKxiYXzB54yAjnPyDYMuJsdzDRB5aYD/y2csQEPMP2
fHAqOa3/a0s5wgFX1TNsvzo7DfKPnSKRG6qz1kwS8AWMhqSGefDIN8KFjT+Gx9lV
Rot2djoXMogYyDUBsOEBXo2XHt5YkXuStueE2lSk3uvY1GecgpXAK9XimsxTIO4b
pbDZrRu7lZKOp+rVZibfMbg89A6ZvZb1jd7inHjLlDOg0pysCfix+P/eCPsFmFqJ
IORkkGFeTMixhNg8gCQSKUuotEECGMneWDUZ+lxs0qeMw/azhmQCM8NFHgrNcfNi
XAoeA/VvW1WTF+cdTo+oiBF4PW8PcE08k4m9MKZkg+/seCfKWTCRftzr3gJYcEx5
skhs0amjbhWzGTJTPVdPxl3p4db/NLkFK7msXVcHkNE1KDmxmnR824dElA+zKB5h
gO+Z/0Mn0lVmlsgwef6me5+HWNYMgEmGR89Wts1av8grpfVUws+PWrdCLNG+8PAT
uH9cI5HRSmATy323JkNPuGXYAelDhPsLX7taiSgv8ncDTgiLm1+eCu18wpN0+KUI
zW61vHKkIHmG0oWklglQi46VIJLbwiHdw3HZOilxPXZRLpI9fB8xL4XFP2mVjIk6
KPAW0TmphV95ymQMd6usDiziNaVZAnI+oK/YS/skcngRa2C7uNZhmLC40RTitgMx
CT/n6rZs3Z32xbSa0UtC75OMzCWDBzQCRIao/kvyL740nMqu8IuGixf9uzzmClIb
AGhseJDtA6MzH6MSEDg8oCJ3dS7catOyI3SjuIFyzzrI95fMBriM3RBIE2Hetv+m
836BhQJfHVOjs7nOdrq0YxxsFaskdNlmpqfZ0RLZMLSNE1tiVTwnFhc6pe/kLBLD
rIUWeLXX3pDTe+FDdDFlFP+rX7P9+e/YcHoUEjet2DAE0S7KMdxMvzBUo9g3ONJV
gbP2oa3Y6+M6rqnjxGqbkLxHnYPagqVhuwTTyUOfSTDCw4Beyx3PfPKZgeR11Wl1
H1jKi0SysOq+gpj/hQUmkk5fJd5I2d22aNAKdbuzJoBICDbCPDJ4lmpT8wr85alw
jX7cqGrMByo+9n0zd24ZmV0ApxUT9xIJs5f9PbREJWoC8Rw5+uOghWaY+C+rRQFk
nnwrcauC8a2VE8svhDNiwSCwp/blSwfij9e1GXhnUtvTgucy+KO8SFYHfiZmVB85
Dc7eWx/BrSZQkFKvu5tiiBPDS/fDHbuxsab9egiTtua/+vWVhcSaKwXZKAZXJ/ag
AeE9RjOTvco6KLKpkU7P6sj+8Ua99Hiej5rHcnQPXsS0FDlJ1s24BR6JI2N/T5GR
mPsBoJL4RlsO8ZqGDyz6my3OnxISFxelAb4uNEvpFrM0wAU2bzsaVURgnmB9ooNY
OYQd8bzb6p9kSuyw0nNOQJmjwsAJxtwmZLrKX2JI6S8lxSqH9j22D8tT8zpT4E60
xYmuv7NpJG8EjZBZKs1s0trA7aq4iLfksJ8MNMNFB0WMWwcZ/beNV2AYsVmpJDUf
UjWOnshL82GrCaj3Nc9tJ+kTudj8PfjFAs3b4fpfpNfp9Mtb9HiakvuDLSEOXWtd
vF8O+agAy+rneU5CmDq17cB1pWt7/Fc87bCWwWWwR1248NewiS7PWZfjA4DuTmSt
4r5McfMx+UP2A39hUP1y/1YXE/lRXJGSm/jVLmqCyB7XLPTsUhYl1B/VyXRkvzyp
VXsjBW7JXI2WebXk2HtvuLHZnpSjsTfFq0WROugnENgouzao/LfI9Z2u9vrUEOiq
NIOqahZCrWzUu5+jLEv0AIm03GHD62RmlByxgtXdrNsvvBMQDik7sHLFtJRqdVM2
hJqfLpHDDajPFiYNqqMZ9joAx0r5blAiqQ2LA0qlZuTZpfQFI9OIn2Tu+DxF4P7L
7mKZ4STVm4nXCBNt5PiU6tYiTEqlPOFA5RpiaVv6duc4wU3gnHS34nbSnGZOXkgY
9yib/RoqMKEkqk1nt7ZoNRcVt/sBTky+6oNrQWeT7qK49VrYpieRke+S4Z4qzYe/
/zS/yDyYxcgFaWGwvHZ4cwbtzj899aJKVBilspMrBaQt0UHQ3IIQ410nhlQGG+Dp
xuE1jGgd4WT1EPVl2JwI+mk4lbRW1HXWtYtjY+79tNVfcvcAVi6zYsXbiw5zT7bI
/LyWyMNli4fcfxN6EHtFK96H6cPnXqLfUPaJ5sVyvg2n8ijf3A+1eRsbma5J97U9
G4whdIac4UPCKNu0yyfKPUAcXIFrwD+1WtfRgM27XwFuuNbHJDXs/DilwFOxldqe
IwNOTmI96E+E/aa6a6+AdOtP0B7Jnoy/4WfAC+jEudhcgn6YoeiieBSHBB4E9tPw
wQ2wUl5g3qegWuSQD9C6u/lvxkc89/5N9dkDxoxjHKVfyrDTFVuq/fT0U2ODNoA0
fOHTa++11oOsdvmi7uP/ch7hYRLS+T21JSCIsx6vKz0aKS1dYJdAKYsji6DMb4nd
Efx6f0qf9DnA6JA4ORioRqVdi15JRt0/WuGAPRhF0/2Mu/npmBhtlwAVje7dqitt
7OGqWw9PkhTTrIssWbLIfXZyKuFL3kbtazNHwdyMpVlvJiQctdxSE9eWOj2eImWd
SvhhcwJeaoZL1obkKbYNBVgxCCl4HBoLaqvzp03nq3993bNNbpbv69k79IG/g9MI
F9SWOld+j+I8z4zmINar72L/Xhw69Qap9NIv1mxUBrP1C0tMDkYjN8DXRMEkCzqd
GqrDsfqcQu9yJHnO38DSkcTEtn8cBCZ3glKeoP412MRMysdcW5DN1EPTJsQQC4DR
xNj8Hwf5bdkVYUxOHneUp8zzVHRsywGHFAi2IR/RtvTu4NopSE3OIeBlOPsN7xod
yUhtPVKlv79HV7tpH0CBTqEnWNogXFPt27eRYGi6q3Q6usXTlSh4z+CTcGyXF1H+
0zgVEQXe4VaxsO9aWhgsGC42YGt6b6wgqG4/qFX7Gz+doqtojXHRTbKy0JsY61FP
GtqF3YPxec6ILwKiOeSQGiFJ1uVLvRsYrnKLcuqyfCO9ROV16lkuLCqU8aeKckuk
mDYi2e5gih/OZB0bbR0kFGTKIrDRfSfIbzslVl10o8Ho33T4ZSokKztvWLldSRAY
H2G+WS7VNCDvehOQo8CEcpJsgI+QMD13wV88PtFb9AxK3KI3mCKuE9Sv8f7eFiOY
fhuX4GBXxgbodttLocamUQNEJ2r2uPdZEyAvOQQ1DmFEsd6JLGiqfwYyAUqtd3XP
hB/7Ks6N0i0y8lj77OqxChnnVnt9Qrl7cSL9zbdb0UeLtvkQYJot96miKy+b9Hlo
s+dq+W++Rq00+riRzfm+aLf5aHDVJErxEKL0OGLyUyUnUdHtb2JZTdCUYxU24FD7
9BMoFV5060BDEIlbU2OuZnxgg8sYBoMx+spKCBwQKF3BIEBso5jUu5HUiUL+8J5L
4xcSygok9JdfW90E0b93YAIVrRWN5dosw9bT0dTSen+ojHhgn5uYqayY08DqiGaU
sinDE8yBDiHuNMk2Ir01edo2xXgAvfH47WdjaIM+q8dz8ihdctX92fFsNNAyfug+
L95YgdDQDAgFhMi+heB+XVq+Xj9MIn7p8zhaAdoxYTyabhkBBCZQdQ9bNHQahN4O
tef7pfheSwfMg1LDe1cwJnGdHZY+dltbu1QwNq/HJcBesX4dSyqAVaO5/HXUwkiV
CvW3tadw1bw24Mn8RiXKojJ219aGVu1pZU7enoye002cMXVoeGJVIC29gAWWZGa7
lmMohk0Ea0IIh0zQ/T1bdPkN2zTngMQT1H72Lszbatw1e4bjRvftfeY7yNT6uIti
FxdMsLds4oSGaRXxtWM5kVmWvbD5AcwobjdMThQXbHWtzuyK3ZdYNXCs8qLROqtI
7tNbullw5SeUZ1kTxeUOKmtYVTao1BvuWeD0MNkz7jSMZQntPfpYH3JR9DGWj6I+
YzgyfDqd571et9ZH+6k5sbtplqGQU4a0VYNC3+A3jzF2Md7O0SPddDJhMR4MbM7A
A36yvn8Tl4DHe6Q4qmJA7a+AbDnvzK1yeN5pWC9ys/iMDqu7R5cGYSkFBOXPkPRS
oVlfJWTttc51zMb/n3qZJ06u+W5s92mtzI7O3YhsHfLAwVYECAAypQiXk5puMU3Y
FspQO3+YucPVisiJmH3W34Qpv5x3GiYrDaGKaRVNM4ARwkEcGrvlczQ0XI3Zp/Lj
OWHT/dVddkyxxxLC2W6xq5TsH5kjuLMPGKmVBl1n7YIrCDZTK1VX2WjZoouLP2aY
pFVkX34Whi7Mva2Caaqxn8Z9dWm1VMJiI6qa1IEGzB2XVeT230Z0oDdvS6nUl+M7
lVfID4Q3lrvWmsWdqNjgdHAW1o2i2UwequxbNcX1cmPlsx7UykJOvRQrzBNKV6S3
dXRcLK1zH0/8ONnZMVk+V2kD32urotf3LG27kp9oFTdvBHQSUCJZmipxOQ8hryiE
o97q57mXV/AEyc4w4Y2zMUQ//qnkiso7JJdI3cbvQLwhLHmGl2IvBbfuEVLIcz4k
LC7GKuxmoV1ivazaSAavS2jr1OMwK40KEj3EAg+Y+t/xyAL/7vuRfo7lFm4pvtp8
Kb4rOHxpzg+Q2neuJVIlLXGtLKgg2J/wwhUxzDBZLl/iXN3cB0gkvA2/zZ2J/jR5
4hfN2b819hvoBs+NW/ESJQ4tOZmxoRddCTr0uO+oNRc7g+bYOBaRkRhZft3IVS0T
xFr5/JzD94iYAAGUnfywKsSkQPs43MDnj+JtL9+onH0uuqcakb1EXvQzvbaiuAKL
u5d95Q+RS0PkwYUycvZePtNpN5QNnJLRLZIi/gbMD2uvl1oRJZ2fEP8O858b1wxN
H8akCrd8b6e8yJAVgYBBbWhw2wTRv1XO9Vy3E8Pr/arPQsTkynJrGB3G6us9I2IJ
ekWq3RgbNhWtErafHAzZ/1LExuSuGPgbHGNfCo9aNd0DJym+MYxQ+tNYXZg6kF7h
eXlsE97TAo2R2vvF+R77Nw9tbY/B4VvVrjlh+anyr99RwStz8VYJfPte7YWOsQ+y
6uPE3IO321V+H80JJLYA3Dw9UiER/BZnYykyuHwDTsSzlNRWTs1Q/wMLT+CZpI7F
OBtUbrR8oToknwMnkMVqc+l24g55+sWavwTtmd/BVKUrINy5D0c2yod3meQOtTtc
9aCcJaQkXd/V2D/hL1Ld31A4vHLCHVby4VR27NYVC6CWKr000J4Sb4ZaZpjfYj2N
aJTTHRg+hj4FuN8TgYAfnwjjq86CXWjY93oOTv6Q0klCkQlW53CTruSnATZl1DI1
+pmKhQ2RIcy5BInlDbH3ZGoMP/b/X7+gmCozEkIGnxzrbrvJnoQDaHn88UuPq3zK
c9e2166K/UThoP1PZrpvs4h+qFFV0SIi1Zj92HfxFNl5djI4+LD+nemhQeS9LHqS
csUuypLmvZvqUsbHQdqRhRdnD/WikWthRJAL5o2QNzG1N7+AG/nVEQBgYZv95TeK
5EjpuhSzcLqyPWt+Sz8h5CJ1+8c1woNKp140EQsB3rTGMGE8qRmYaV+8gvXC1/aZ
VgvzSntWT7Kt9VY4Ls4DX8srSzKy2Hm1ClXy7c/NHcSuHpD4IQJ8tNudJFvQXz2L
JAgbG+fZsbdTPr58t9BDnjuSnx0cnhnyqf/4k3/TVZ2UAdL3JbwbnmPn/Q16RcI5
EWj1IOtZeoDf94Naur4K7lygnSMtkz4BawH/8isOlF+7nNtDd4YSNdHRF2vmt37E
VXqTe1N/2fgzPuHdzLYN9YV47TWqrpI6m9Isa3GDJ8MhEuEU+ZzIK0WFRMjPR1Zc
tb9m3Qlc4YUrJKEmShgsWEAn9GChUShI2pQC0ozvJLOTIItn2Zw1ierYmRXAFZaB
8Dlrn4/rIzTD+vFfLdF7y7mIbsoLdb8CT63f5DL6vpXHIV48LWi4XFu7sAwmc4g4
Ew/TB+yAN/b28RPWdyK1D5zVNQRv9HGDm63YMFpagjkqZ3/CGZdYYUkdoYqlFAnY
65hVk7rjaGeB2/7G6pcU84ATd6SF6l6Aby/yFz4hFHZy7KziCWoCx8xqWIjkzd+1
M7JNKW15Xfzu1cTWMv1otnY57QTEEQjK8kQLL7J1Tu2VP7mzyIePP/uI+ySV64XS
r7GdoBGh3XA/cAo97qjSfYhBeNElScEMgefcATChqXQh1wddfLwR7BBd06WniZsX
Dq+42wo1TAXeRB5vrHRG99hxKE2RtPU2foauqoJ85WT3uZzOKh5eIfWz3NCsA2su
cfVzANNd7W1QuwkGEI6fjg==
`protect END_PROTECTED
