`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CEohTjE9tzCeq8uaUaOIgi8yJWt8q2WCDoPg8t7GOfILSHhei1BKdKiPhc3BBR1H
m2k5ARf3VUa2P0nl0yQFwE1llUqavHGoTdpbNOrZdihe4FASriIVw0drSYqKCDVu
OB8lVG1ehC3aXztVGoIEPcC/dQRG2L29MGVOt3H/9I3fi9zhnWyDGi3F6GFO31Py
Zg/0hWeGLsrXQ7R/Sq5KC1yXpQu3tIZ9Bafi7w6Sq9KlpkEywkeet0oT+BF9x9fN
LH7GmcogXTw6dsZvRMo85UTupIGbQlKJUX3HoTG19v//KHlQq1Xvdgi21R/FaER6
0HhuAuPFFYBRDU0z13UpNyqndmt2cQgeumGCQaSdldpJmXH406S8dql/okFTKzQb
iFxEXkcDJ9cOTstdRWWlDzu2cmL1gKIjHSxozyW1d7IqjnBre0SC5Va0SjvyKHaI
fbOV7WvgzJEH0/LfI6lPnlk8KxNs3cdRTDVaF1oMUvFQhPrEUYA36AnPxjXcQQTA
5hNTqKRDbvF/4rYSgn6NpRQ8maxmML9HXxa4p+ataEyAyovJkBG2FCIpNhLkDn13
U9wOGro/7Gb5Kb48swTse29mqiDYRxyck3oumDK6bzMOrBf2fsVQRpv9W5YYeOSZ
xyzH79r+S2CHRzm09/6OdoQ+6B9/seu2ZXDkGm+VwSSoUgH0FX8sNzdJOfPQDAjw
n2yD2I49Jyc17sZM/1SIZa/bTboQuXCtS6H8uzFQQuN/3cfT3voc0CTlBhaMK7+U
rE9QQVsVi0l5zErHFM3LSZJ5L26suzvWJItwL776P3epdbg6zmeu+U3NGuL8Vx92
OSQ69N2LZAyLGXccweTK7+2Fl/O1ZLz/Q6Lx1bHxPx0UyjYcdfc51ACk2uigViK0
XDCGmNUzsYx70MfSA/NE3rRgxvtI/+Mx4Exk9bz0dateFirgQUKhYL0TP+nsUYDb
dyKtD8i51je7qv1SFOWtf1rFUN+4MheXzwaSVvXCMEgfAQz6NJ1D+luyDdsyCCTp
ixYVbZ3a0CTsgx4cX+eA8kHyq9WZ1ByOgqaT9eVGi43kt3UP2znq4YneD+h/gDfL
98ZClr0PZhEg3cBzt9fSelhmu+Lb+qj9RUmbtIAslfAsyL4Y17B5aRAeW+a3gwCK
KIjQvOuS0geAJhQFwfkmRF8Y8X84oMQWKwcssD+oKcyP1UoJKqb4N7EsomlmJg6K
uwYo+gCIU46adVkylj3F8Tk6Gc7mQuwb9QDvfCUAgeyA3IjUT7JUhmYKVNzMTRi6
CekK36A6nSkW3dmZZd9erUU0N4zVNhPg5XUocf06yGL3hLJGbNRncfy/stE2w71c
L624tcFD7RhxPgcIn4oUW114w/u14MB3PCXqtpEJByOyl6Qvth9Sg+VBJgUbREjG
Y48JF7modt/dvXSvAHnxcjdcb8tcjpx5sbjS7rdEYeBu4vY99TOvKAFaQ3MM1jP9
PJNRVHKmgVe8dAoleWw8GpPFHxXIrkupcXfZ81VRV7kDgR7suLVHAcdOSqyaLF4M
4dK49PAObBWfH5qPugjIAwrBaojjRcoRikNlf4SHKIcKCNSjwwoInNUMBnibnF2L
lxSdWVUW0qopCOi3t27HnMa9AkZD1P2aIRNxnZh2p7q0KD26MfMkwrhmWA8QtcNJ
VOoA1iVXJppH9zZMN9PPzzRN/nvejC4Q5IIe0JCSwSQ/D5E/Hw6fcHdENUzuW0eV
q7MdVpO6ejPFF4WRKIMX8I4ta2lHm+0ep46RnowPT5vqOO303Y6ZNMJ3tCiWU09J
THQqvTBm0tkV9e5gYG9jAINulYCaGkcwb4Wc8vfgf3KBlN8HjdAhd84btUttQGQc
7j8x0OcohwREFkT8/IKqriyZiCM/W9MdPbYYbTZR3TFWCnC9HtakEeUsvDJ225eH
kZm9AcinX1pdXiGwxntgKQ==
`protect END_PROTECTED
