`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fVT0lIJSgg3maXP/KCHOgiHoIiDfe/l7Xa4h8lfHClrAAOCAHOCV6Q1ok011fiOV
EaWOjR04zs7SbQuyZ+AXNFDdV3giardU8ZuNjFwmxomrQOzeKiUrhpsZAqc7nL0K
WshNKYGHFeR0UqZW2Yd5bn8N1k6bp0N9C9sjl1Kc+UYgmD5Vf6ry5QAOdWjT1KKV
qlKwJCNWzuMF5irIs/RSLe4CpI351B4aFLt3NQA0ZNya8RPnnEPJDqxwXN3+//jx
Jby6XqHCfuMOcxNvtdV2bIxwBG5x6arqtXte6MJN/Aw/hmGiBlsskZ8TIRJJi+CC
UxUbzXGGBJAx81tiOiV5cRmv1ecC/4T0DGDMFyciUiHUTUKKpV+Ga/MwQlPdsRr3
/+w7NCZYQ1MX7bEn0VQ1azXO+D8Id2pyof2sl4GQlUbC1ogsO+3fhD1FFX+c5XYy
unQBhWZM2OhgdjeHbM6JpYdN7JDfnyKkWo0Y45ctxZbq34wEiXWHA0S3btm+SJLg
hMzaalD7jeYkRseCmOIHbcwMpmNd4Hp6WgD/3W9e2C15zsf8mDkR9DUj11BCrWGy
XUrPNARCeSH/WFTxhT0BJn5bz1enKJDb4wylptZKIcVPi9iHP1KqPjPbu/dM6txm
9j0BXmKsOy6pv8TpvEo1cWdksk7LU/GneKn0bIYAXA0uvqQxcYg/8nqegZy+1oy6
zE1stnr+Vlmh9BsOB6a9qvGF/lp/dEpebAtUYjP4y7AojiLuEOYFaNEgLihaCnpG
csTz4vsZOchYgjR9drt3CUCAXePTdoB0dns/tk5O95UrpgpXbsXBIaJDrfvjhz2Q
q6oXf1wcsBz3GeUEu5YlQoPX+On+Bx8K3pBGv7v+54Rt7TUXD4cczLVUs+oPb725
Ht576PC2hCtfRln52vfVjK3qGAhcHf8ub61WWzKxqfShK3D+NAA2t8ppFgXLdjzu
q6V/9hpkjI9jcrkv3q7rEoNv6iq3K8oLC6VN5PzlAGbV7xlj/P6dGkwTFjgeRF08
VX1tiDiNYjsrcQcVDHIkMv7PlUtkbhHgFZNuSaaVAtUOu2QD+1uXPY5DNfX8mTlR
MhF+n9/vwrp1eGXWSqDJsA6vOMcfsTSjwxD3wcIcvRG/ib6zBa3zClecrSGbGqJE
hZAVxe91QTVNnT+DVGf/+g1RTF7mfvR4+1Sj1hMNlWwsCDQD6I0jRWoVdxTutlDz
n73VyJK3gAb4g8f4d+DjLYa4p6jNhYUBEERECbSUmTriBa/GsQeWt8/B2Ji0Rbh8
grN1WdKufy+YiNky9Xbf0pP+ZrH8Qs+BJldNXivPukO+V9eCUn0x85D/mv7OIjZl
bRr+uoOYV4orn/8kaXgC/+09BZjnqIARX0vhFJ0+O5K+ShX6khLMOzVMsLvDRxp9
Z5Syx3bp+sl9bN9giO8r3bLQuQJhN65yE8bsaK3E2yXdMrgBrNVLs0Y0UBDmXiyy
RBqOodKc2ZytGXJD9J4SyfBh4rZ+V2ciXThI+TfmVYA=
`protect END_PROTECTED
