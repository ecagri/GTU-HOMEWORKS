`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R+kbKWK0WU1oTm78NCwP1QyNBEg0oc5ft4lxifUhHo6T8W7SnyhxktMVcdYk6s88
27KkUYbbxutjSq4X9NRluM0euYQil/dK0gwVXbu9+2MGhDmRWNZq5VSswSVxCyTh
4J+Tn5PukAZQ1VuTwfoG6OQF18kp+vbqWCOkxVl+ZC9scwSIerOcY8ImXOhJdmgP
NkU+Qa27lU4m8mpwXlP/z7QxYBlC3Mx+Qdnm/LOlVDOVr9n1Q2G1oRUY34TvyqQO
eDgX/Gcz6l0FFz0+g25tqJ/NlMd3idwFJ7YKcrWPpMjqSsT0KBiIwSUjPYKBCeLM
5PM6eQuzi8kxmizl149Lr1OAHOWVsZDwj9nm6xNQVlSNohDK3eTfSwBTGEMzwaZ9
DeptyKeSpGsR4F2OG13D96aQNwZhPbHys2/3FwW+P2YRUT5B9VWF8e/TA39FsxZD
YFvAMdUmXh9JhzIHUJT0nnaHAquNZ4Pb+WVWCtpiG7MP2pDxWAvS7PJJoB1NkDo+
8AdzliFcybLIfqGW13R/GztzYpC5EhFyJmhRgYytNg/G0nLtFzRKDczGwUyBiXH8
wzRI8RCy7svx+eIm4j0DFrrsuqGj2wWs5Gnza1NDgio1U8RfDM4XbRKfPbi5kNpG
3F2lhyEDtscfa2R1htrJ5Lx8slZjlNumoMyQk9X5Re64kcFZS6bgrj/VQiA1X/Km
E4J3TmAXkMMlemYdS8rbYYpjwYoN4lgil8XO2SjPEshkho7olZlOBInJYO6CaXR9
HV+BRjY3AvdHrdgkpnjaJF4dBB9wjRkgyZHyja2szVoC59GVwmDtrgXA50mzoHSZ
jnrd5bkz3MB2fD+fju3fEB1yHNyrDvM1TUG3tB7HfhZtUUtbJ7RZty7alNnFxleS
B7hq3f0cKr4hJKJrMe4LVcjhnplkhXqDkdxNrhV7AQoVsBbSM8wdIYI+fmH6jt+9
nuEXxzE0zWSSG862gLX3GfA1/HOIpJC1JzK+8FRMbWoNwGMvzaox8lD3AcJXQmd1
/AfKCf04YeJODg58a77CdBD6uSzthGLgMzKeaPNqs2X5M8YIX8bZ3TnixhSijyrL
NrQ7moOtBnX0MIJK9/qyWmSdW3KqDeBTPBTj0mOAYL1Cr0bkwjgW6ypPDhe7Rk9r
acVRiWCiJSrC01Enfbos1UskqvD7AvVFAlvU18PE8wz6mMIuaIaNXvH2CULB4vrt
+u7mxUj7h6QFPwH9PyO1wU9+xrWyAoaJCXTU8s5WR3OEkYuCiV9Ot6eakC06FLXF
DY/aaTN9qeGQ3L4IzmeY3oU+clGDFfGEB0hDgaTKPL6b11hwI2OLrL5kG3sMNF7d
PTT/3+1MUndpvaAfxZWVEIvGi6bbD/sK8XmWct6e6ZIIA/swIT8VS+unQjxBy8/f
CUC9QDZH8qq4EtslrFu0HM9KNvnknL1UXvsJyIVkb/zEoY2zIY3/N3kFWzrZLhf9
wPsATPPsith+nNqARptaJj8e28vDifUJ5rQQbNrzkJPkT8HerjoalGD3GTAiBrc1
ygATN9J85Zt2oRRHdLGCxrxS39IzkplcaBrJuPa61wGhzHnC1bcNpGWzTNnszBMR
hWU1m6T7qkYbvxUm5pyREpD1vQVUHpkHGy53ARQ/8kVScR5bjkUnTIGE3Ov/aBW5
mD4EgMg4PY+r9T/BhMth6kCNGz6a9b8Q+NLE3rbqQ/q8sRraUGqGDHUhppdVDFxQ
DvHAZHBYCSHnP/VONQ89Ag+19vcKfs1qrJjue2oDuRnjSHV5juAsYQjudXyI7tis
xpDFpAhBmUk5Fls6JRVuxk8G9LhFuxaIA0fQX3ldLgXKkTehRma8RrqKEPQXgtu1
z9inwceu0y/O084ChqaD1Fl/izPfWRewAi5w+XNCV2GIh2AMD7DgniHBwChuFrBQ
G2oYx9DQ464RkyNlJG0o1FqYlM4VYwm7hEhsSY8fzNaVMcJMbuNLSJP7IPzZlG07
w8H7Zvk2Z2d8X+7fa1iQXwK3CgvA/aTU7KJtOaxZi0HS5NzpTn/1R1fdeAUKNW/M
3AZOvtnF6rpK0Ui8xNq89gtTzU8WrWVn3tOhKR+C6bKAjWWiFgASrjLuH+aqrYJJ
hZQOTWAhIaL4fVpmzNJSj5PoS3eYLa0r3d3GHm6Js45s30Hkv1Cf2pB2FoVwsTE4
E+ctVawDS+x6CmE/nJR/mJ7FyGCIsoBko967pjLbWa32uOI5oJ0ak5PESc6fmAtb
nW1LKAnC+9pqFGcshv/KapazE04RlwsFYLwbPZU+2yOPHXTJpMBw/2opN/t2tfZZ
9MvlZrEjtj1JOecVneBK6cAaFtRlhP314f2RYYYP5WH2dzjU8lWVpi7DBp2ELbah
jFf+4lhJEDQKZyfbR+lYx7T8mCWLv3oaqXEDG9ZoCQPLOVEiyNGBsJo2Rpmu6fyH
qFMz3C/IEa6Vw+PRsTsRyx92IqVLklVfY13ZqrdF7MapCflfjUu1fpm2gqx//ZtN
C5OjesLSniUjqXFCBSaGVYaaQcHVxAXNEkFTt79FRCRZ/Wl0QVcC216PZ08l95VP
wqIuiFyVdtVlKRtK2WnzozqXwLhGTKNtr2lO7dgV8JVrbE/pCXJfeDwvz4eSFuxX
bDP22MIok/e/w+ZIxicZ236BSMdSYlh4p9rcPDdy+BIcaU7WbkbdeueE8mtpOpFa
3tVg292nBsYzUdkA5dzO2+SwIWrGeHRU+TwhsRALlrsyGMYgJA1wg66Tb66/7y81
I0kgDyN2hO8Mnfr7+MmdBO365/dVdJnBVl+5BtRNpZyvHAfEke+maC++GN6cFFuH
RqCQjxE4iguiEQMbb+t/VuhhKU2Ic6a3jV1u8fYbBXHgSQrnpX3ZB1qcNGH3FDWU
+HLjAGAWgbxdAORAbsOU85qhazqbn97ONhUC7pW97wli+u1SplQ9ST+A3Jgo9eVX
TBvajbItxgSInG3CyKBysaeAx7r/DJ2hN+Eb4rRzKHHqRjrpk3jmulxOlwZSNSni
EZV6vJduhn6HYpGYOeZ9kMPNVQ4OBYCojwA16hYiUtoy0Xoh0ROCa48wRVJRdmZl
D96gDN09fx78/CSLQODJ7Pdt9WTt0QilCM7vJrwjjVJTBN2pqANwzFViw3Bsc0hj
LzvURbh/pLms8q8YafK8IP2eOufd/t7aHXEUH2rLU7858sh7hixpMdXneMFlkXmM
yxRyiKic+ET0VaA2PBm3vUhTGdcAlnszpOJ3Agq4iVuHttP/VBWl6h5W1YS+UvWN
8soY3eeEbcYU3VzF1k28wMEd+hFb0dqm7EaG39TbUwCkJ/W3o4wwcHroTt13+eUl
Y+JDT3Qt5CxhwoT+8uIDTLsmWQ3pqS4Z8HE9oePOIpGcJ6wmIgxHtelOE2XMeey1
/nn8oDsiBx0pzxez3iANp93NptMeGdyMZrst00T00DZj7HXgbh1uLbW2VdK+2mcv
d2oJxLLlhsi/hCXQjqfX36+dLEWJY9/cYX/Fbh6rh3zfEBg7Ft3vY3ouUoMb12ug
jgjSsR2dS0PIkbXqm8PiNatcZkvjUucN8hzkuFKwJ8NmeVZWE183zjYybIxCIzHJ
Fw08Z+rcAYyQHrxLAEjPwwP0N1enT18C9nwHhJMkUlSEUXa6FlkTtyzVSPHxDdnF
5LNOLjoAMRqzl3XQllXR86hPUwxZT9WcyVMOOeYYFDTLj4JReN0fcC+3ApC3RsrG
YUsmcrbpzCWmHHSF3xLsEkqVvkLyPt6Etg+Cb784Xftm5rUfkTtVDzfscmmuz6Lg
yKSSrOXV97iqBIrTyZqzNjj6QLUq+Kr9IUGMPz0t/YyVm6gG5yjNJ9Hh9ai71e/b
414eS0Z42GxAP2iHLyajyw==
`protect END_PROTECTED
