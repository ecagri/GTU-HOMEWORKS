`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4x2747QXEuTW/vgaSM5tJaAN32TbTsqb19CR4b6jZlHxI/5tCMl8LBNGD6LQ3T3P
iU1rJ9TsDlQA98ZsYCTjWMoH467Hlkdm06b/9piVsf34dUdnvrrxZrz1LLX8tI/8
4lVB2GuEDfYDd762IezdYB6FwSUvBpnbhTZiyvDhzDKIxiGhBc2s5IxUEbPbIKrH
Yy6mDkNn2NqpVA5w8+bmT+Am9ESAvOnnMw9hOX2/bQLgB9oR+pDPUxJ+hvowfQQE
i09ZiHL4LcuCyDScaMHCikYnVKRDRXIe5KCGzIqHHdacwQdxMbMn8bh0Ntb5QWaG
w8oRMyySBNB8BuhR5YP7N4KrAheFWz+yZMpqotYyZZhDPVlpwwOY7MfwbRQKqs4T
51Uq5/m8+JIn3zhCcT02h4HisE31t5L+cniMjjxlJpIiAh7XRiBBP9hxoDTleNrD
HwM+Twd/9Xcdcaz+9mhTZpffYXAcRQAi+H0oJukpMVER94tNQB/pBWmGTaZPVm2e
f2UZuvwdQ4PdpsBSd+dkg3FR9hRTc8Vi6JTPlPILqVFS79UHCz507Dg1dGLWYU4G
ZjmnFlDMiDdMYTIO8UkTwyQAr6rGSVMKU6IxYBxEB8RZM45Wj7iWO3+u3holXiyy
GfkUOIUtn34o7tQZ+KNRfXdHs89+u9EarcWalmbsn9ELfyEUkAHuBjzBzmwDm7Cm
Oxf3ZtS+Zv4GwU2kog6L/Id4/q3e3FKQ/SzY49Lh8ApB7mnNxS96ERxmdZJ1xYOS
pjm49AVhXpCT6TfELwI3apG8bJqCsGfkWamGOq/Pgu+LlmErNecCBcreWm4pBRf8
gIN/9AOMYNcruLenlPo9K6vquu/xzdK5AVgU3E5/AM1kEDwUECZWwYTn9ncFaYpa
iyjhPy419FpnKcgMjY//L5nGny87454+res3XIbtu/fwUSAK3x6vuXlaBigZEdGk
jFlu7IUXKK/kFm3ojz4zyuicMmOczn0r37dhk88aeo4z/b/b5aa/ci3g74GwCj1p
fXbikZI3K/aG+rii9TZbXnYfkLDcc8iNql44vvlA23md/bS8C98soLyFgNKhvLC+
QOEz4gmEDyo9wGMrd4z7UAY+Uuun7N0K1QGfixvcp23jsrw4aCMNLn1xTPiATcJj
0UBk/m8HG/thvOG0pAz//8eK/EBCxatoAtrem0T7d/1BC7ac5XQJ7j8+PQX5XdXN
RIKfVylnPpA/9goJNKPRGYjPliVtoZvNT/Vzug2HPUVCjj34vDpbkSMwWUqIG/hV
/UarX4FoBhMAdPJleM7i+AuhV74OFKWWBK4tIQow0NggiqKFZuODut4UlC0FYgTF
doOFujghS6liiog0lCePZEKpe4YhMoCQ2/1GlNdSnInT2/eGuZP69BVggLMKLH1D
yAB9L3Sao9arFBerr8RQ6J0TagYeMGiJsYaneGKjTbpEEWNXv/LKf6/9l0VdSmyL
INpMCfnvx3T6noTX37nkPYfXbdn8I1t3ZfRoOhcm5/r9OKswA2g/O+q3nFIwF3/E
HmXxWRNVqQ9XK5ry94wifFu3IIilMP/xXbWkjWX3uxtSYKBboY51Ypz/c9qqs7Ha
uiBn9k+h1r3WsNwxRzZ0CWVksKtxFcZIWFsdicT36iyXckJcYzy/k7LREp76+G2W
6gyaoS7AVC7RacxQfRSypryn4kngAk3fv4IArEOrmEhOBHDK8n9d/d44XRcwjtFB
EVURGkKuqQ7pSpknCZr9qDclA8SzBhq7Nv8egWBn6xgE1lggPI4CDqZpc9PPF1ae
JbQucgV4v2em7TzmykcYZicPjxqLEQWI6MXOud1DDek=
`protect END_PROTECTED
