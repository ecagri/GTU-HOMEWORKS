`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ce8yvw3OVs6BhH2cB86wQlLo5st0Cc2qr0cRPvzkhQbjNCMYS1uwukfv5r9sTksL
Zkjvrst+3RD8aZhsZHNLDCWcmopJGUx2HstpHImfxcvXhi8Yae6L1WteCBE3swLT
8Z6jo0kNbDGnVhsaildc3q5b3OTZIkXbdhXlAXQEgy1yH5kAj6e/wA05t+gND9m3
g3XboYRSS8dy3ooiS447u/31nqnxWKQ1t1+sjyd4OtlBcFqF58X8lWcszK68HldC
tM5reuFbHML2SymMnXh+Sdyfrc/A8/6H4+aa0tLmEyn8Bt10p1pmpeIecb3YgnSm
tv8pXWZMuCXQm4LMMxIHx2mUKRlSd6gd5XT1fcUWrq19C8A6GWECLJZJCgK78iX3
j0v+UN6L30TJpiG71oMC8YALaUqd+syQDb4aiNXiFgE19L2gKkPyjiTmiPgg+U33
sKVkQIBYyVD9qm4jX8ycmifFHdxeBh/ogurue7p7xYZXxLRpqxMxxiC9w09z1PrY
004SqABgnEeGA2DzHojbBjh30dMT6T3H0dZxaoipaP14KWIqOQIjPS1/AS1vsPIz
1jsr9/xeKNpZULaG0Lum8qeOyMz+WXV9XLSp/rj7YQcIHxMbNomv/gMEkHhXcZg+
FdI5asm5kHbxBfMkC72L5irNalSJWn4D6Ge1+Lke2s+Ei3lQS9d9/Q+ecaV8WIUq
8ByENaYYAR1PCSYXR9HbZU0t7aMd0k29EXDtQ7isoHeJosHZHxjpSfhdbbgYZCdt
awTqLb9D6GDYS7xPAzcuEMRcgNudy0WaDCZR0kh6qfe5UGWZUkX65Bn8gLaAsl1p
Wsd9JY87J89uuLVlKpMn/Cqr8dLrQRuhPskYwqU45gjfhrc9fbJMDVEEH4Pjc/qA
zTyHovs2kO8gSguGnurLfXEsVEZf1ucMWiq3mmpd3CjX4Ndc0t/+Lmj7Wjx9fMRD
ThZJ61EgPxO5y4cLaiuTM/r9fN/vkficN9FtT1SJDRhOKwXkVyA6RW+1VKt8yS3s
4QaM4RyNsj7A8d1MFzsl3Pj/ZgEUD4gJXqkDwAmrGefwlPuT5NlUmT3eP9DylM+c
oNCakWj4zW26w/NVBLJCdxD+8fAwegtJ/5UzXZ0kMp8PncEjs3Ky4Xh3gHQ5nYFj
O+Sj2BHLevQW+CEW72pWgw==
`protect END_PROTECTED
