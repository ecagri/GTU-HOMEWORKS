`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4SmRVHE2wuJiL1tKkIP7PNGWiiVy5oP+1xkTjfof+FizplIkQ2pa2pWhdypOjsvk
2JqEIr1dKDlLXrIJWS3Pd44Xqj8/VYh5R4teCJMq2NaJxU9aPlMQNxcIWl8H0/P1
apJg4tEid2wiMu05R77QGobQLX093iIwpKXZBUq6AW9m+AJx/ZiPbR9wxzVg6r0P
DKTGIh7dHhmGT8PM61RAG3UTBnYC0AXVvMkSLHb2Qy8AeSi/veU9r2jqDpaLx57b
VhdMZ/ZnXf9TjmwZBv7AZWEUHQByGs3BoGcOon6wF47w31oN12D68MR4Rp60Adc1
0NIXL0NXCn+QABZVT/fDkyUa81ES1avYMvINCJUbqTnYy8r5HlGqznvUWTsz2AMJ
hOojXjKHzzNXriejyywDLjEsuMGITMyIjSCnMJZMF+QTngg7C0qnIJKnlIfWQT1L
zfZMQeYzPbt1wmUrnLs3j0xdBM+qs7uoIArK1f8juTEUg+nnCRrX34FZEklsXdMo
MTl4P9312+YlsT1lc2mMVpHlK2dPsbMVLERXEvFzjzoWNsvGBYG5oPaxU94lycVV
HSm5gvBefwlmd6nDrELlzC5EJFXjScEwh8bHI6LuEAKuixiKHshXM3F2HSR+qDi/
`protect END_PROTECTED
