`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
17JpGF6bVUG+2syiNzh01BzHjpaqU40xvlXutvmvfqvGABJdz7ZHtkmH0UHUh0Aw
3I0jLn8W+gTbUHrbunWpj8zaaN9gBWhVf8AbU9UR9382NAum8hiID6KYVhwjA4rf
42PC87IJfp0R1mctqbTzBGE7s+WzoaIrDHpZDcdZE2svLHsoLGw/ctZSrgoUZhkL
ardU6knUGJF11kmBOVsPqubC59MD75zfPriqhdyFZ5qPvdITnR1DXmX5lV6mPixd
aQQLZy/m5v7q0Kn+C/GJ3gn4qvR45sv+4X5F9jEKkSpi9E0YoUIjbzEwNc3FQDaK
PgVUM88Nzp7qPVmPKyIYNgRpvlJUhIDKWw7iOI1GR2T1Kd0xShdlq8uF6lwGZPyi
WmRyN/lbkFsWfu2NJXoS1bZwVfjqvnRD80g+9TMStFzNembN1jLUBEy6LYlbnU0p
n9yeRdAMg2/gzWwuILiL4amHOTk1qCF6adrdyuFqqmangkAP1/aCg+DR/jI8EOAj
SBhZV8vwi+tS9MCY5wBO8oqIYsThguYRipxr9xZgPrxoCQtncbTDbWZQyM7Lw92u
ZjUte6oD4UgLVj41E8AUVzFt5Uh819PUm+7ynknyJrMWJJViJFyMh/D7U9OuB+jr
DX5r1saHkrO2f2ueEvL5vChrCA4HZ/Msm9ldfbrTy59KtIekHKvHwWeRDESyVXp6
CgoPyIxl87aEXW66o/AT0alCIEzJH/b/puho/2a7TY8vvXBwy/ZAlN75HqtR23ms
c66BQ5me6R/A1B6TrqWwVhTC9OcNuEAfkaNUBUp9trMxa1nM5tRoqsJoNDBXTfTh
NaswG0+1LS2W7+og9TH7HaD7zFSJnhava2B9VFDG83UgqFkx9DEeSiQzO0qGg/In
SLnshv/TJp6l84kxL0r47dijsavhdqKsyM/MiuUTKrpFDEWDVa+gAdoWag+lps5P
LbZa7rsxT3DLk7y2O9gCcUrFGFv4G20Nvh30qzAzd6fPo09DUWJ/lu1bu3c2dszQ
KhJUxRHROtB1rB5tXi4+5U3Rno1HuCB3RkkKJiQRoCSdr9HMeUFoQyFsndDOk9eS
N+N30VP1I3WfM6A8U4o3KhQvUNRY3gLgOPe4eYCshZ2d1LOVPj5DOmlBDIp+AEpM
EMPZebFOsyHeYtnceWXLbHsvNw+bJ0EHlf1e8mjvW/iko4RoF3WFXLhiPtAgxt4H
4LKURf0ttFxK/3pRah/PX4annBptqNd9Gt+gBgezC+CAHBqExcsN8tbKHjauNCmc
LY/QEilDRhm5+oORjYq9KX5cFQGq90eYNGxrILTR7aeJ8ZkNpNeLsNl7Rm7YDpfm
n71TBZuhbLY6bfHHYjHCSORVknYbvLxF9InOaBk3xdrlYuBMNnbi7fp2DrGVI2zW
igenH/GXFfKamwphvlFJjWzdRKOi/ubtGJHhColLbYzTuTY7kK5YllBlHy+/0ZEM
5zmtpFk5Vv7fVru/Fe4rqWt9iERYimYeIHwusvsYAzlzoe6u4xER4jmM4u5sXfhG
Zf0I+yDMPw/u+dwRjuLtoeJ1PK+kIhr05xb3wkb6o1/p6JnRDFh/okHVzgimCKDS
ohvC+b+6hbp9uGWw/tGcV0ULGZz9ZWQt83zhcGuUFWIo4OlzNeIMYqiYuKeFc0Xs
c2LNqk3dIutf1n/rVidwttnRKiFK3+2jIowQIRr27jJfzoZRBN1cdt37VrAoK+b7
26aMhCjIGgc9or1HBRiftT3A9pKIqgJk/y3mE0BuMO0=
`protect END_PROTECTED
