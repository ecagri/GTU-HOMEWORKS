`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WSl64Dzg9fQFCAkiC0Ml0KTgArJevjBLQPS+K/Y0GirvXJkEjHzDXBG30V+5w6BL
VFP1WgmnZXNm6SrGAI2/GKk+epSOURC+6DVQfGLV1qeDB8wMivF4ydEsTCCAGD/h
nS1VszGZFa2L5ZbeMTuSfJyNPNwNdNzhXIggyQv5t6D9rOF63kC3gpIOMNoj6C2A
6HuInnV7PF0uY6VojaBlmNbUAUJ4E5cSxevAE13vtJX3WkmbjUI97mBp0/LCq15K
fGapYswnUkCuUIP//vjSc8O+WHehTSxisu0su40026N+GIQAGhCSRKtbSKqbhURG
OHc1J0R7I4juO8a51UcmVgNfLdZ6EAuWyPP+FIWLxFqD2y5JTx7Si9WCL76CZf3H
BgpBHIwvseALTxTPGfsBNA8yx2HimDgNGw/4UFOOwccdeSJITtcVGwCBI70zyhwr
0OyRSiJQRrN6bG+ZxnKa47tZ86l5X0buxJEm/d6Wb3xzdVAxP9K7QNyPCTtt9X1v
wLF7rhBYKg957dvXYtmeft9JO0VPSmIenqSQU0dxs0FhLXbrd91qu45NbvvhOleX
vEGDI5V9vGF0R/4oybLLaOwzAcvRKyHvjlMg5ty6OhQ/kOCv0Wrb5STxMHjkiG1v
MfZqomWsoAmLFgI4GDFIgdd4LyyXSd4O0L8Mp0uUM8R3zMQ01ymd+VLk7iIjwyGO
qc7UfzO6fds08UxDiM5KLh6zTeRM2PwWGCH6qIBrCUlyv/QkAG2lTxCDeopO27+S
wqVvr3wfe5etkusQhmUSxNpa4wj/301+bkhChBoNB0uKJ2ISDbhLG8e+Gqx38Y60
h/KgQx997V20puNYEP+p8jcFDK/VIVORktJ1MLjt44kNw41qdo52YT+9PmdLdocU
w4wYf4UU32otpGO7UiN1OcIxHByNCUPxp+c08wH71kA=
`protect END_PROTECTED
