`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1m9PU0bEzIhsSuxax1h8gUkk/4vegptgenXdePzxlOK67VowjFNVRQachbev3WAs
Osavj+hZzBLQEhi8mXmAphTFGnQLEbcQthmmbBgjnOxwp5CAE7d1bm9gOddQisFw
eKxQ0a3722crpvktr9DcWJMh7asdMafl20IsTIcR1k/VX029rjZJ9tu6GSDfKBzW
aHGd6G/IegEJDQbDLf8rst2Pc/fN54TZfpgIflamQs6BYdzIlv7dDeASDSTR7WH7
4wTqHgb33SssSls50OrgjzHZ3o54Xb6NmCDThfEu6nTBm1Mka+68GR+6awyN5g3X
BJv5NfIwGKoyHL9XxlUo99S7Ra34GWyOq3RVklOpTq1oCHRIa6w0EqzeiLV7dXPW
Ons6S8mmwLxH4XgPM//tyXTpI2lV47oQs5Z4Fo0vEsKuCa2tHQGrfeh0fBz+Wco5
kzhkDp5+v5EKNEo4st5VbJHpNv0esRQT4dQLvLySsw3waD0C3zNOKEomrpA/A3QJ
jS/MKP5Ud8G5371hY2StoFdRwdrI/BnsPl1R5WJrY6gvs7cMOXYBbm943U50XKZL
373UZqIJO+AuC1iYoJqHK6V6gZlk+GbQWpDY1hjNLra8wF4VUtMb4MqpGBgzRS21
W+3Lwvo1qu3UtiMGQw2oK7jqqSVCtBU+1GaKEI/2yBJOfrkAJ7kFg/b3QjNdDRKf
plJidcgoRXVtfloag1Kovpz5yZ+ylOy31iyFmzgxIZgx0ddErNgSebFwJiBp78HP
wsZ4BmiC2GG4BiZuIUGDaS0Q18v9y67d51Zyl/PMho0epGx0brwmEtZYB7yX4Vly
o69MnYWpsglUuEyPE8YfSCZZv0U1c5lbEVEtiaa03DH6MERP5yG/nFCgH5mgR85D
eh5jPMiS2fd2daql34wuHfox12vObA8mGxIEo5+Orh4JyMZBAq4ABe1lYRDDzMtx
6+VQznc7vkqDDxp2k2/ETWS5mfCpQ+CIFckDqCv+IHzS5bowOll8v7t7jymaEKzc
FZHLqrOi2F6avI0dHc6NmKfo5VAyeyDXaLx4qz6nHzh14BU4E06V4BCNCnU4jAuj
BpfpFVxtW82R+LfAMtDw2qbUW2EXrpDM+oskl8cI3ny6czoAUc8WQoJ2yXAU883A
/aOqKUed1QvkalhLL3zy9mxaASXOX5/C+fNQmVdB3sd3YsspRQ99AsMqsZlIUdJg
Vd9FOo8jY7F4xiM/t2K1hEPxky+tJlWwA11KFMeu9PQeT2z8aRSDHpM8ePCDfx4M
x7qgZT2k9WjwRhbYItEDjkEaFsIr8El1UzqDJx6xjbNO48b/suyX5bpigX6CbsrN
MRITDHYw0GuoobulN/UID5hPW7oy41bbQ+wr+gKxcciF75MV3NTSsixQhO30D7Ff
17/rcM1IZ7mCC9bwwBnPdjr4viC+JGz18j/uTcdAeWTIDKcVvXPaei7LzE03FOR8
Ek5Y2MRFWCBrA62ySJAOx6fw4Q96WUrryjFF492eR+iM+Oayf/PSakX+IXs3BF5r
UHZBw9rATjYsZNpi2sTBRdbYI/G+wXGkCIQAyy1yGSMZvOcnizwVLFoZFnwQ8wgU
Ok/DYa6CqLcCvZH9jQ8IGWPz9Cllk4D9tr8VuJpPqGi/dicOGBZIOz0EHS4YMQ+q
exNnvm35kP+sAtQm0q4GQMfCTXYm7YjPvlrUsW9ndaB+LkfVd/RKMfIMDC56pPXH
6nxPUdBY/7o1FfknmEnSJxdCAU3jRhdGf0UsP6xKxp9pgZkStzOuiMiEjnigU/V+
RCNHDFpXjVa1yPyMAKyhy8zkbfyz3Hsb1WZKymYmRnsKuiawaMFVR9pCAQkNLrDk
aOq5Fq/WqQ8mvrB2udKWyzrUMzdidKTMt6eC5DRFQuDb8LSmnObkXIe4PmtXlsuV
fjYHBkqupt0OqZw/Rij5BtQr9W21t52rAtaP9GZ1fCuMBvSkLU3rnLetcKIQeDrN
tl92zqk/K4VQyTDGHWQPvW5H7cj3etEFNjh7SgCCVU3qqO/2lxTswX0YWVSzC3Rz
nsgZ4UuMHow+oD6w5AMVMx8kjR2x7gECPtOCBk3AtIrjA9SAVkgzAEMzDqQ/sDqz
sWbwjo+QLJ9AT+Y8sY7uoeRSOtrx0xoIJ6wUaXEfu/Ng5EJb/fR8EsktGoWQBcE0
l/1NLz99BaqJsv/QMIrhxoDothTPkt4cvlsVOyOoKkWDH8ltitlDQUZeEq1oLsrg
Bz7Kahl7T/fLePpU9gvm6hW50SWtWTmjrxhGElZ9O7rcn7NvjHHZ1iJNlCy2NZ3h
RpRu3L/2dbJZGCg5GyaJIvtoTPblWwVSiuMQ+mVvzvZyb++Q7VOob5IL8c8+VUHl
Ti8fs69gtV1Ivh/CYlaG2zqnyQb8pGZgT+pCOmdAA3yFeU0GFoOnsiGbOL2RUT2l
sBPp9oktgNN3TmJRyidOiGGGEdHTX7qme5VBgXn4gnGQpLxprxZNCgeL+OVbmzfK
wXQawfKSxArn5uDQpeUkrvFQWqD/eiH0Qz7gOa1p3ydaH4AHjx3vTpdUvfsK2cKu
Ju9OFzr1hw8OSf5Z3rHcHHGWZGeWQqJmAZE47gsZOmfrrm8uOT+ZMy2La0fykDGz
1L3AIej5k0NyKonC/EFcMI+MMw6difVGz+bPeflCr1Vexi1ElQV2YztggwNzJut0
DoU8LZL2XrnyaYez/5SsXlE23GfWorT1Le9gv7zPl++F9Kxn0FYBRrR9NS5QTu1J
CYvj/tlYnhmbKhBVr5qhHJG4AbCNy7+LqfyFBkLhG54x7w9YLBVipDNHNeUEjNZk
CiDuEAIlDgLvNLJEUFSCqKNoD0zWZoLHHuWPOV/YQ1KVUU+bUf02sEZZbHVv/H29
INS080lzjbSHGQnUMAhNn/mJw9tbuP1GaVN5WuTU7trmTSgIrfGbvYpii9L6bYxD
ZqQSMGQUoGR2c9/FWlzSShSRGoKYW9kKG7drxqr+4i8cvikcsP0IxzmwUCLtDdi6
KpVqsfcFGTwJcCguJPXMGR+k2nCGydkcmrcCxUCOhbveZmhIpRL8tNF5H0dhwNa0
oqbsBFxGz9Mbm+uE7TJ9VdENLBFhdhWyMJhu7WLVdLI+GDMghEoJI0vAgIrRwuoA
Gpy8jl3gercKkT4oy17VasB7bKdnxY/2W9owNQUa01XmqHGa16J8bQzGUKG0I2wJ
cmAGPB3CthmNBdTwi556ITt3uNyZJAxdeCyQHwf4rEi766ywvMvK+OyANXxujLCa
uWuREu/niWIxeEqGK313QU7jw+zKZLodgJdOjH/tTxwFm0Er0+3b/DI9Z1eRmgAV
hFH2dsCvQcElLtMYqImZE2brnQy75RopB72LTQRwb5yTFBO9LY+l71VaNK1yzpRm
sBQ5v9N0F8yPJfyQnh7PLwbdMrSADiyh5PSExIjQuzDYo+HG4q77mKfpPtwmCuCO
fgt0Yyqqq2ue0b68mQRoaJ2hh7QFq8pfIfCa8++9DdbbxUpvrGYcyzZxuJUKpuvI
pJp8lWniBoqe0K6JrcPQeZRnUsf0iWbJehL6YbEYie1tQO9TQFLdZeX39b+Be1lw
1oE9f9VidjlQDJkhyGTqDAlNSVK1WC5Yf6vKCy62bUBUlMbDs3WdmObCbnDexNpQ
AnccRTJnmnOtTc7I4MFtNFDZtLlJXvDIP6Ukoke+3xXahodK1yvQS85Q8xUd37mn
NNvR98Eme7DW35pCduZ7Msjtp0gtCW2ag5yyLrU1g+WD2n6hUXx7dN1BugjqUxIp
SUgqdeFko5UEYfgkkYHeFI960I6Au1Yyw1qDcWa0E8oeP2f/HcpLGO+o/BzVNupC
ZXDtzcUr7TVmo4OHVLF19nN6hrHfwvVCG2zJzbApWYBcwoh8x4yVHQAQHur7xheh
cw8uscgTTbtsLAPbYu9+iPmQrqv+zogEDjg4D/VrLIpH5iesO9/wZOksid1ySPvN
dzMvOt/GZu8ixIvcnp8cPRTeTRo54rwtPaUFuEl+/rqiXRG1FWL8RiT5YWMKotBQ
WpplRbHE/2A9bRt3wDjh+ZBDd8zGPteUkjhzMLup3RbWERIDHb5g6ekwtWwbQPou
OjDUM8CljwwHo55kNEH6qwl399yMJahg1LJCQLEKcDhJPxdTAnXNJxIuqkfSWqbL
Vki6B7nVSC4Nzvm+fINzAOevgp2kFtFb4OTXalbibtcHc6t98vbn5rA/O2XBimed
1PoDC81FkjmQSaqPE59m0oK35QFh63lDCjkgijHW5LGfO3Qe/UZKP2GD/lqHBb8h
svZTLX9mOE9u/dptypXQ/MTVHBM54aEhGQtObB9jEsNgkcCtgimQOwc+NZiPhe96
2Z88AdeeCSZFxjHLHyFzFfVi4ZxDnTM1/VrHAqC22sIlldIWaoyOPkdDQ9tKGf6g
GmGCeG1vNLm1rCVhGWd5FrLANGgZQHyDCdrEN+ePmWwDHcUok2o4SqC8DsK5tbaK
c1HUkK64tCptrNfwMylmxdIOTcqyOshBaUHjN992WpOrMzISJUf6Es8+cZQKimmZ
CivucYB3yOi85hFCd6PBcgKJtOzUAnjwWSUH2FELL7Pwd56wttK5z7/+0C1i2QKe
wGOgwKvf3vke/aHYHh0YqJ5Z5/Q2ZapWKpX1vv6mTrpCWbPvtY3fJmX/W6Xh44ka
20BeGcfaxf9HWSB8eQAjh6neqY6DajS2uahZp9G1lR67a0yLiXiiPZQ/JIo2s/GA
J7nxIg/gK4LSss9tTc+sLdKQVWZHfkf+f6E0kwxzEQwEq/M/U7pJIFbp9SkXsOad
AjNJttSK7osKwwfnxQePxQhH80nL357IbvpcnZpReEoOUI7n0qj+VpiLMPxMDyr4
uB9O4wxP1SGC2g/z0gOH30smKOOc5R3F0xD3BW7Xh8XeVL2GuayugO1Gmcx8VUw8
17gb1Gf0N6klpTdatrdGUr/jfGYaurrJ57PvdS6tW0LWzZuQC1dj2YE/qdVscady
JOBnjt/6lkZMC4haIO9iSep+T8hFDSA3XEiunv7Is5FV71TOKItMzanPOQB3PDFz
hd43Ru+X1K/4vJSWhLYjcYLxm+XTNDhLE5oUqznqAgkxRabLljauppP0Jf7HXF9B
ClJwmHKDM4Gc7is4aiMPuxWu/Yk69gmQeoasFyOfySWoPq+VJCv2NZKGFoalzAs6
6roQkOB/UVwhqG+HUoNaUKKaqLS7LVZuN2mENWDw/z5dIdYVYtwXMKFqGb/LyTY/
SAk1xfAf/fBbKsMB9fUU/FQ+exCZXiJ3pfMbNgyW4kbaMM9IoCHjjRPTJrBuMsaU
D06icToVBm/KhyAbPMaOyQFC04krU/pr/ac8uiuk7nUg+vUoff+wpth+xyizewCJ
UlOIBCYAjKzMeR6rQ3VCp1bL+OC919iE/5+TVGBztJCncDNnw7lkTnxob6rL6x0u
QZuH4IcsuCc4OJla5iorpVmF5e/R0v8rqqRxJigo2bFZw8BitpkySNSDxxqFggZJ
gimEyzqyn4TaEtNPRGcTs6NWfn0QiwOUZMjBerCxNX95n/HbJDdvVupfW3hbNb8y
2tFZiGz3i38IvmJdCva9CdgXxHgTdFOQ1vsI1QTgTZxv60NVajG0ybvZkJGapGHB
7ITsKh07ICZ52cpnwrEi1S0OH8QerMsfskcLJitZqP2jztm7/NvROLKewZhm2PEW
AMG0y+GT2qk1QBhoQg02eo+Rm2JaylyyKl3TIm4vUo18SXYsCHvEhV+TdIbbOUmU
1qBefunHx/YcNEQ3URZfKR8j8ZF8217AF4a7nWvhip6tONiw7L4TGMMS2jvBP1Ba
pudN/nSlW+U/vs/Cpme/AKlbkvb7EgVbKfYxc7uEd20dXD/E97AFYcKx24ZL86tV
f72/zJfMrEYyCAGsYA65SHGt7fCXZdqfRy6mHqsGbA1vpe6EBQqXl4odP/R24Mv/
gQ35zjZBAG6V7DbHr6Dx8NsrMTcoDA3p+klcYe6ri3D45kAkezonHTqjQ6ZuMblO
XbZwAfhxFkC44XXl+g/eI8AwG3c/MfHdRMm7KJBFpT1eb3Nkl/zBt+QXGQ+VK2m0
HbMAJ/GaPvbiFi5om2MAVOjT+9aQ1KNziKi8c5NVflJ1KH3pkNIxzdV7v4S+s8G4
S6v204gkKEjm93nJbrHJ/Kp0rZh5RcAFBK3E8ZNAIWBItWtNg6S7olmJxoI2BS2A
VT7DIONEYDwizfUoZrNCaaqrDbftwVmUumQn+bycf/e2e89zI7ggKo+r8+5zT1K+
w/KGszgq5BZfnQV7anY09q7+DKJviTLSq+2WRBd6H+XpEfvpvwILgHnJyy5VwfOE
mZR/UR0BdDO0gWCHYdCAqPP5CpFZYSFRQiteZtT68+wy590rpQsWwQK+QPKM1c2F
6VhA1soYDg/9j//kWeGMbVF8+24XaEk7UeIT4lRQjJvmssle4tKorEAKupVUyxuz
/Y1ljuPyM4j9AuiysiUvqm+7yYwFSMNCt4oAd1kasxwgu7wPSsqNJbb22ZKW7jnx
l+4iUt5eoo2onqqWwKT1YdjyQqEADrybTsUsT+O2JkZx8xwJ3oT0xu46rRyg0S4r
VztvoSp19+1rij8m5GYEubSzGAxWkdA5eFpwPmW8Vals/++MlF6fYg0drqarwcms
X5CNodnJ0dJKfyzQQ1aX6ZMhPWOVLGphHnljaYjS1wrycLpciMTDoeSA0wUzKgo2
I20wqFv0KPm5ZfKdRNf3xXTwm+c66F7jIzQxyv2mJAaBPSdy+9SQUdbX2n80D6ii
c0EESuldo4GeotCSBeUolspwfNfCBNCO/szw5jjJpTD+S1uaSuboapb2iUg4f6F6
mDTeiggeTMdgDTAlSIlxp2h3w9kfYlRbWj7ng0agCnmSrdciN7og2OfXI7t1tUPl
9Ysi7jtavM4irxpPMYtIa1zwNlPpM+5tVD1gMREvgECCZV8TYT98Yk7cZ0WR0xFQ
ccXgi05OokImbb9r0iGEyTrjmoY16KpX4b1caH4w8bzPDZwTcTKiN+2lnqShr2ZF
Ma/9JJHbD19UgBj/ADY1VZrZKiTIBqKrzSMdTSBMTE1zagBxICGgpu9ZIzl/CbWY
E5W53acjKfKdyS3/fb/AMcT7k9hSWmp1e1wOWrcM0gKJZqNxzV/mAWDCLdcOTHpV
YSqWCkLxuDNNZ0QmhFGEWFS34xlUqvNKMcfi0d+XPqAAdbD8WOx/X8z7XWbDkflo
8GsDXHzuf+/1lVzvt+Q37cvTN4gCZdAXxjoleWWh/2Vr116z4bJERDXEvYWvfQwr
nu1MOwHC6HhlQsVe9oZanvaaGq0YdhgFkV6A8LtWdbk7NF1Uz00nEgfq28bkVqbm
6USO3mhgpee8Si3Ky/3WBU+3qU7hkC8yllBCmp9YQQtHuOcDwCmW48elX8PkDBYB
8Ok0FlvgiVb/4AsFqWslg9OMwBtozNtkMjVyfvKCCi5zIGMps32k5o7DEf201FTA
E50cWaJZEwm5UWlN6mztyrTL4NqLocbx2XmtTtJOG3MyaZ+BQq5B4aGuwvbrRkhw
qmiyAlQAQR3HhOjoRfaD3a38M94m7ajLRYI9+PAu/tAeKAMjx/f+hVYeok9BJdQE
shhf/fiffPC93adfyaEdU3URjrupLLSRjfcCpcG/U7ewbI6odOKOoycrth+yA+PL
r7KiMhs2jTv/szo2oxIdnt94VbBY1HG0134IUkozj/VRyiHBrGyPkLtz53K91d8U
Eqaq1SQMJfB2IbYNYZawUVUviWgo5on5doqEeb7yshcge8PpViUB13IRP1T0o0RS
vaduuucpAaW8ST+1uhulh9Jn8l/9DpprmgbAGvoXLToOnUrosD3rLIrx7QGbSa39
03bwLmlB/sOveLrkwzPZaKy9BBQtOBNiTp3qdEK+Q66wmRG2hDA47ucpn330jl6J
cpsa0VxcruMIA3b3fWolFd62/LjjUI3DUU1MQUbZc1Bdhsw9AwU2eaB88vP93gA/
NaHPp810lB8JJ0iRfNeen3Qmsw3KDfwNr+bIgA5rXbSyFjMc5g0p7QAAw3eGZ7xA
j+OcDSx9i2sMSNFKQjOEKqdZnddoCxvX3DqmhD7XoDYxcSOPHor2OazFNkzu6pYe
f1xqP3uq4xyNKrYMzkSxPT8HMyIyLXA2AwHkjD7f+0K7ix7lzjqBWT18OcBonN55
vicfqWBJVKC5rBUip0ILUgE8Mzpo4hDBuEQuagor5LoGTmE6pgSdnKwNTsyg9iW+
K6aVV+cNEAAzJo159EnwAi67yMpRFMDYtntQ7YDjFtw/VoX7Po5wRu8+RQ3sj4T1
tmq+4Fz1zVyQZt1pZTCgVRXfnwOEUjd7MLearH0h4HJTqVXzVF2/VvbnXszKySYI
PN2Uor4Vu/mWjVTYWvhRL+vx3CVQINUFqraixCnvi9DJhgOKuQGRk+lbGHcdy+OA
1UnGode74fQCT04JFudj2cmA3bYH5d3G2+T7jKncRvdPRZDzBAWRQhRNJZJYTdN7
y2Bao1j2md5RcW/OJx7Hwzz150pyySVgrlkeey33NBlU9hbQCnS/ixZvGkBPoYEB
0zRDl1SftJeOu/Aonp+1lpKUJmPCA7ncGGjr4vhAJaw4HyYXayvwW54D0MRVgD+x
nRVevGwC8Zdi5h5YWAbVbGQzBJ9+heIAjrqAt1M2Eu4VeA2ADz7wkTAT3ysQITvc
G3i+MlXKrAN++jmyKPdysEaP2+T08z6lGIsZLuWb4oO9xKqbbqG2t4uGBOD18Aqi
Qd0fU6tqkjWpZ/gqnG5Iab7hNDUbPvdACfGeBcwprjgl36LEPE7nn85JSjohG0in
985JPo22GNyP11uaCYOfj/IiN3dJq3UG6gJaGFWSXMUZt7uk5dSLqkopHgTrRjDh
JcK/efv1QwRFdXlFibkwm1wymYOjo5/zpmV1n3TBI1W5Vg8YUTjk5adgMuL9CRyO
lDnm6taJj2saRd/3vJg7v6/R539Kb3lhAXCJWDecA8ZqXrB5gUSgE8Eiv2didqQ4
uKFo/T8jGOkrhvsc/bY8fA+4WvadWqrBBa0XDg2kaRhfZ4WHxLpqaCzb32hS7aNz
50OZOCz6ksno5wv0iw0qs5vNIeaI/LBAFXaaXOI8MSEkOObe+rgGrYCwsBZQEusX
kN+z3frKjp4kxZPQtFGLR4/9UKh+6C0HWdceJ1k5Zu3hBeownEWkgeOvLZjH0aZL
sIBTrY+Zjwv8sLZX03tmMNt+ASTAW7avNgGapcaaGchdsMjesZnxDxldicaXfSRy
M6pU9LgvNetdrjqCUI7Meei4s8d+EtlyT6dhGq9K+jTglE8S1xt8UG0UMrYV/HrR
STyX0ES4Fzjm2FYvamM28Khy47xdo6sQUnKbQWGtj8p/2h+f1CsHj0JoX3xGv28A
hRm4yz0xyYQD0U6Khs4gkZOfluNKrLzyvkuv6daMe1GfEvTQfyJNxOpOmPKsd2N5
oG4TxGh9qtI4J6cPgovQ5JvD7GEKOU8apK/O/Yh4WSYTEhjT6OOXcbH+ZAwXfIdL
1BL9g0pIYI1aJq1ag9idGFS+4ji9K6MreG75hNSIxtZB42Bqv2yzwTfwtDhUn3uB
9DN0Qw0PVfx4qJIiCBJFi1JuhzLxSswLndJndomZa7Tsmb57SF/qiBfxMmsO3laQ
2teJbWLWb0JVGMDWsVNmnN9qnfdCKkmVEt3EquPrw9cDxUxqqpeHnpe5bRtRZIcR
P7+s0Aj0bPbgEkmTEMiYAJzJFwfGbZPqlpifnnvzxmHL8RPQnHIqbg2l71EjltEA
3BuuhFzgEr2L8KYxTTheOLq2y6LmFkrAolxilXdRnFStBJl9JeOEjzFl4Kpzza+9
8BehNhO2e/xGW+kR/2USAVHM17rAtWuqve8y9l7NE7HvYFOAVed2XtFnhuVo1SA6
v5W80zwzWefJycYQ2LtlHcBjtau9NIdnp86nlZdXw0n+kgA4Hba3L9zCTeo1Bizx
erVnqI3o3yglvdKG2E45SX6vQgIxzeFTmxJ3lRPLOIWTtI5xOUMGD/Z6WslpN+sv
rn2zwmp9PgxPosl7J8Bo+aEF43d4849y1Wgx73mUs8sxkk7D3mY8UbDoveX0Slz0
0Tu7Ivw8nO6og5TCoIv8cJKa4CWUWTb694JiSFTAxLG98rYlPiHyQDZP/4xYMURL
iViESfXKsiSHDFYpN/Gb4XKoac9f2bzmzS8NCljQQuhzhZH+Gg1wUCQHcL3KmX/n
p7ltEbsgd0pHaGj2IW8Ee+yG4My3YirWI2FjKwLwYMTXFFPrfQRtO/jJatUqTKeG
V2iVhhwIRdK3WsiBSpvPUlLoCRoxuJVHgc01ZAaU7h1LLBQJAvbPAaQuIQUAd/MP
wMAgvTDvNoSCtFVVLNSBGuYRG2hLrF17VmgcAMRHFCkOu9Zbb6CPFXMlm1i5eHjR
EayvgBuxzRkZf9H4ulgOen4gRnqIekrVPjWzENUNbMh2f4A7m3U2auwaTpic9sYq
r4p09ETADXSDH/KzJAqM+KcE22PDxJ110c6UKNgqXL4G2p9Us1i9NLbN7T1vUDw2
k1Wy1+0SFTxMXyWbeFQkqMRNM6J80QhYszwBw93SjkLd0SXUt5Z4A9Wn4tgmziUj
iumcpgeDaa1g83CiAJSLozBgRbkH5HeLLzkz+aBJU1sY6SUf5h/uJ/9U3YPaCrUZ
na6mRpth7zriTGTj81Suo4HcIqMjtAo0tSy7Nva5U9PvJgIRN276ET5LznxXSYmP
7jY1+GbVk9DqM2b7vHgBLVAXueYgtFVNmfv3LKZxIu27/iTlvQAz5v4fuosRSlg7
kqWX7G5ZkIpFdCzceOIJVame1OdiWc8S6MP+W93QYUnslPCJ2/z4STvHP108Ch+D
nN6nD3PAW/qhEFUwcV2ZnrPgAxyCDfJSugpRvuZDuidfMFKr7IfqQEO//oqNB14b
z6MGavYdCReHKQC7q7eVAwAMCW9yfuQGfl7zRGW9L3Sgy8rqJ41KUEVHKdvVm3Rq
1pOb6WUlIKj75naA+DEfCEHV31T1G69ga3sgZv2mOc9AvX5TM4IfG6c8AYX0np/k
fwLoF7Z/FlsITsdcj0FNYrkfio/ww5OderhGcgIRnPIn/XORceIg6ecyVjgRtKyY
h4SOdhpzmZfH9s1DZpjcqDOl2KR2hy6OFtyoEmduM1rT3mn/AnqDCERybBCnCGPm
Mp/8NDEFjqdXwWYm8oYXAzXVXmOJIOTBZiQ+eQCaPoHbyl7fkrFtVEd65JoG4rFY
HGcQcM/XhI0LWK2cW7OLrE/9owIDw0Zh/5luIh5XX+XIwqG8I/mt3qSaYhSe7sUG
gCd8WxBcIk1yX1g8xWhLeFmHHyvzp0fQgOj8hO0Yaa1eWsfGPrdYBdhD0aYkiCEK
qCuZlB8OSZJyiCrXAEyKLQM70gLznyR3RuOVMr1vfFo2l8NUzeFZi48tR8ZktMxu
2fkypR7NGnTU7XHazq6hbAGihKMHRyh7norFk1sZ3LnHzVSx4p48XzbzNnaEEeFp
7z08Zq0uxneQSRKov78f+ZzCS4+mhNzpQH76lKJ/jeX3qiA+DJiuwEMhzqNvOlPt
FL+MBMesqQ4Obeg2NEQHLORH2p6o/mXO96KFgvm746x1i9o4ZhpND9avJQpGnJR+
9wfCejK5WGmGnwywZJwr3KM1xvghbsMyaF28Dh31Ha47/9gv4XqnBafGAWYjlDrc
xmqgQ5Hj7tXKuMPkozP0spT2RC01JZy9s4qhA9GSr84/jFGH7t432djsffu1/ZOf
3NfeBvxuRvqiNWwLydvoO5YSkA2aW0j90qmTWubyZgTd78Sgiq42MiQOiDkZjp13
notMeywS9hsVjmcd5P/rBVO8chM7wYxvHPsMvAIiNoc0BRubwWj+Lunrzm9Oy7jH
LprAt9pYJWMCEl6wSdTCVF7H9GQoFynggMugsHK6jPJ/TQlrXWJeE68dUTD8I1FQ
dASTElgHSOR1pn5yj3a5IZM/kvWhZ/H+HwCicVxhgpsqd9mSYlFjS7spM3UsxI6F
Hl1h6ChwY8+aSTeGGfY+WszC9ekIG8487Esmic8Y9NGcyv5vPwziOrVgXaWlPdhE
LBvgoz1dXI7+H7fY/kyfD3/Dgxa+xzIhzfx5bksO7flVSkzKBLyylUVCQ34ApEuS
pwcuBqibMsywqr3NbuEKDHZRDyH/UldrRIahpY7IIAyBRWSGbcEEY/hQZHRbEebC
QwTjK0u5DetsURWmDLXp0rS4sJwYHLftfR/fWTWRtCGBdiE1Q6TxUZAefXFBPEyL
Ne4bZiI8AsoXcwEx27Z6Z1dl3Jt5iKN4ivTYe+3OeZsw0iewKQxPseH3a5BbwowG
EcfY4BP8jefDCcNdAljmC+6+STBXsYf2z6fBkOxFVd8Af7FT55a4XDYpLg9oCI2O
E12duqJdUmmAZt6gPJiaVTeV4mm4i2Usdahr4D0Ih90qp6hSmtgAn/Xd7Da5KPIC
pa1QbdGnM3dvZfvZakoUKC2zOpsF2y79N9Y4kuiY13r6LJQrHwMjQCfBcxjAa6H9
abCgYYwLlwL4kHzNRJABBInO1UD649cTKuYI0leswS97tAud8TyOVDau8VnAI32x
3hjw/IeYSm72kz64EtuAq+tiT1WmbOxypUY/F/7LAC8SWLVxmda2QXlgYmnsmg9F
4EL+4oGqs/yXyOshTyxsz7MpQXcit3NB/E8KwSBvUuUeQSYFytfaanmQLQsw5zwL
X88jwwIk2JOxPJVKKKdRp43H8/kWPkGTGEEGoiZ2i6jE287Ih47946miTY1V4qRD
LpYa1MMGzLyLu6+7pPjZXoHIzUUG/2eOKOgWtVF0HoJaiE0aP9ewt3F0p4W/QZjp
xVU6KUJmYd7kbrMyzPgFZrEVJUIuJFuHhBwvX767BCz77Wq2/vy0+az97wohoDz1
HZrXBWQgnLLr35BK7qmL1nGT8JRT6j1LJ4PLZbGMLs2DZhibLTphUy3NptZ4OEuR
Iz8Rd9KicCgS+P25gpB036KiissZSUaRilvMxDxD1kB0ofOfUa/LzSsuI33ZYKK3
buPKtRTiawQCAnYDfwqFF6ZyKOIbS1L8XRdn6kz2hN43E4KpMRfC9PqccRBFlv85
jJED1qSQhyLe8gnqbLUsCDBZxXhW/2EbPOp5UKZSqlW2WQ3hJo9An5UB0boyieeU
w+4t+GL3+H12gJ3Ft3KIx90Ho88NktsomXE/u9tgKj95sdDe5j6KIWacP6Jr8q9w
FCY7qNQp5M/0mXZqm1BTyCiATglH7Is2kIbogEL6qKk1+zeR0/tJ25CYFGTNAaL1
htrIzfJ4RrvIUvRaUW1A3L3v5muB8kf7tnyqK1MM1kFlovNVv3gGRy9tXfh9wx4a
lukrWwTBa7iy1YeOHt4YO8qrQYsL3nSe31HVYa/XfRXcybqZCxCKhyN3BWT8iCKs
wg4f3j0z7TRj09YHeJistThZnM8CkFQ8n9rBEO4djnpt+oUts9XYceoXhLzVB076
LtEw5J0zUVtam1dlEoS/O9IH6XPemHlRVdxMRTr18BTE8bdbz56JETsBV+BbNbSh
XJc7qaTiEZYZElelDmh39Z6P+fwb8GRrNBZyuydwkB/vAMaADjzRkeCtSnY5/NYi
0851UDLQvpt4p+8Wv5a9AywVwerhu3c/BaF3EUsrLWRjUTfcOgGawewPea0KW3sl
6Blt63TNpNCSGErJEZgbybkPjufbuUEavsX0teBJxP+l7NlytoyevUSN8IaH+Sqe
F2tOqIC7u7jpVPru3qFZCyK0H51eBXrRx4vcfkWfoh7EDcLxPqH33qAA6wZkW87S
K51IO28dcXXO6Y8VGHQroiUm+q+typIyOBPAeb6PBJ2vpeUgszC5Cp1IDsprbaI+
8NNXvX+cLu2kSXcGDDjF39mvR1SPZEF00nlecdd7QjNYHaWtmQygAIiduEmUyN5R
WtMJRLBCJEtHAHUgYX/ktsYrvs6GE+IpUVvElnwiE7C2OSxeS+mKL4xFdVB9HAup
CQFC1FSqKAsO54967GYqRSVD99myHj9f76V3Yzj+Syz6zfJDMmLiuO6ElSWUnwZj
NUQpuVSp3rujqZ1QOlagUErwC0nUJweYZ3Isb6tpGWLqUFxKsdgyUxpKn96AfGHv
8FkRfEtEsRstVNuC7ZWIwEvENK23p/MgdJpL5GAoffv3nkSZwXhsFKt1FgqADLkz
Z1ZCy1+pq0Y7m7sZQfbIDSvrO6kWwNSCjJgIPciuE9IitRBxiZbMSHBqpGjgK+YB
aTZ4t6gL2ZAFRaD5BC6tZ1TozFh5sCnHGIbpU7jfHb/NETRbpcK/bkKEYaSd/ek6
t7H0iHGXrmCPsB2nqbK0iy685ttdvpKYJh9KoJBhYC0x+5blE8i6CKgBhJRsaiSr
5W9uzybBdlK2Rn58zoY+b4bYWMin6tnx6o8QLaKmzfO0h/5Bt2ZZ6y1I4UAkF+bD
WaUHWbll1NO5UD5Yqh7cv+V4oQnPVoLu5uD1nuVE6XtCBYzoQ9w8MtE6ytPKlAkD
kWaaiAC9vrP1XAENRY6N5gjsgp+z+JuSJ+aofVZ6suaS7zrjP0g0XV2rfQ64PV8M
FKkOvIqChnXHF72ru18PXb0KTrhHGtqNgH8opHTcUWLLsBDxEMKzxZHfJj4V7vuy
YQSCx6p2Gxy+82ddcokek//fXk4fVtfvO5YlH/HFfqY/pv6v36l/nBCifhknNNrw
5moSTKb2Fz8PqWzRjz4KCQqGm25fntQVPbEo9ihlUc0EC61oacX6HUVolegnaRvB
KMI0yN+ppn61lxGw+KKHH2UrsKcczyjd893xw3Q6h7qjL1VRTlhHpEHo1XaHZwff
/DS7sjNREwfTPUa0Z8/cLYVn5rxvGA622SSz7U+mLRzeWh6W25lFZj9BJkonjZTc
EXEir2Tn2AerlgBJ/1cibEYGoetgWhQpN87PQYqotwDguTgE8G1rQFj82UmBTM8Q
x1WrPsq0x/7/vhCMfvgdL+4MM3M/rnAp+y9wEGAE5M4sst3ZGrR41+PcpRWpSc6B
//I3+fnxXuKVI1QzneQDpYLZgCEOEKRyMJRmueBvP5YDjfgv5UvK4sdWlplB/STY
d63mS4MUSVVgXpxnbD5oNZVMuR000MSbcwSI0lMizIsVyQahmt1Mkjrh1s5pzaEe
G1ZR/uA54duI1zQhCHu2Z/aNMA+H2vFZpBEf61jaCKzxj0HkwY6M4pKa8PllEJ2i
QIdzOIdXaghP1ZQEtuFWQlIugVGkHcoc/Hlb6zvmQtgfHX1LlT/M1QGVaRfMvpp9
ttacmmH3psL2acqFe0VcugO/N0PitBdZmmPxc5Fh4R6Er/oJEka3Chj7xeCNQ38y
E0UU+gVgsU/qG1zOcjuA473OWnVka3c5fEsHnZ8Lt8gfLD6aJDFeWoBBFeOqw9ec
z/nyDXjfafIt6+5IzT7jvtucpXIm6CUeyupERh/vmYdApSh5OKm8+HYDBfviNM7O
bycUt/eMX/YGjnaeMI5c8XxeZe4v/y9SYvTzx1kdHhwVMYHHiPkCyrr4A74YQQ73
IvZNYosW615U7gVh7kJRL3q95O7kGdYabp++0uOHtMMIarfzScOngANzpMOdee4p
ekkWtjiLSuqQFQHrY/TUoqztiYVBG07ge0f34Nj18YRupyJvRfhF0ltDyJZPOd3u
oXWfaO6PSjX29kpLx65KPYBYMkGpnqGFu3vs7KUfLy9t7t83GCbt3xmpsPKx7Gkh
fEHspY1zKuJykmBBcBVit5erQMSiVheUrj7RPR/Jv1z2ae8Y4+JPdFlEsikMZUW8
vfBDvM+fRjTwk6fhuEavQKaz0nQRATVcwpk7IVg+h282EhnoYAv+wuJhmV+Q7Qsm
eEE8R0fSP90Qu1nwusf/B0kx6+audaVPA+NOWOqPFXFNa+ETDF3fSYP6z3e7zMgM
XDbL0IB+cbmVrW1isw4MDxp0bEY82IEZjDy0YB/YGwDVzBSW/6kBxb04gmoBGL2T
WdIMCVcfzgoev7R6/Exq7r1OQoNfnSYHXul0CWY1qlCACmV+olY7Sm3lvOlFeUOl
hkXpteQpkXBu+SodPFSCek9/7MPO75eBc5WiPRVjuE6dl2Zwnw+uzP7JWcZjGhhV
OknOO84z1EdT7A1eOvu2VPrfPD6FS+26ocyfrbDOtETqTDsbk3jE7M2+Clwq56a1
/wd9uRqtGfJE/QVMB0j9cofef7EovmJ5zUMsKTQrUMSYxXnTtBpY/5a4Wdy0dZWy
Gv5Vzn4IMVq3U16xkVsZrAdtA/U13upio13dJq2SFlF/2aNFtmxyUe3iNWhi9Knn
+mXx4WW8XwgvSmnMG0ODxpO9ahJWoMHTBeBt++iAWmJQe5LtVGXsDCvTBr9H2hgF
5z28d6l9GaqFi7+bys+jw++UHizyjlffEw5B40QaSZMM3+KvpYqabC6EQajmOybO
mBV+SnzXfM0UTYuzXjMK0E+fAdHtL+zs5AFTmAXjYt/he+QsFixP3JTO6NlRX2oE
9IoR+TAUMKNefg/4ujmTuKUqPtufRWB4ucChqcSlsP/LUrRn59MkBR5MeArx2Y6O
77qbYnwbqiYgahEozIHjf72UxqcyX/H11tvDdFwPWP9+iU9Ui0gH2rFMGf3pOaiO
lPsCUYGb6+wTJSYouJDjktTaxcqIg1ITnfWLZKQb5ONPdK94rgLaX1AF4xK+Kbw3
/y08+u54pPGWm8ug+zLgoBgaEQvupmOVpjmZMzHDJA7C/1NUnMmER1A3p6zkylPu
m7nUn7m2UqdcbTsQwbH/UBFeGd8SiAW2Xb8+CGXvEJPlhU/fbaKBXSQbEnqxzl9F
WF+Yez5GWtxcr2Ms9c+jDckX912g3PXD5Oj6JT8w1bIP7R6riTMZ0x54d5aMSYPc
0a2fyskZ9c365l//ERXNssa3hAjrYs+qdisqCf0EaT0QKsD9wnyv3/PIMHyGCGWE
m4Y09yPHsh9M+hWRdkz63V81FNHpI7SjB6vz1hH+56vpn+W9QOs3eUCyuGE0JW9j
peB3nFnTOOZxpxXDB3dmDkM2gvfJecJNorzWK6Q05dVtmt55I9q9DXTgTIcRHoVp
wmFvswkcD6XISct3iGVLBymsid8adUsGk4aNcc5eqEP/yRwNykDqPPdp2l+kuu//
0QifxwrWzTCEfmFonkpkzcsKNd5lHQA4FOw8RVG/ihuq+lNlAW41Z5GfSA4/MyjX
/3Unfk2+ASQOGdi/78js8hqLPSDdaejKegkphi6J6vKEiIJmAbnrO/FNQ61wg7xt
qOhS0L6TBxrZ3Ij4Z+qv5936BJVYhvudNDX0BbCtOqDvaeqvisK7rEU2rNK9Dwyz
UK2IF/WNF9axahb2fU88v2V6Ix7nbgg5oQzLZsmonAl/wErM8MkB0nw03YqgoBbo
yGTv0Nm5v4zBiuoUDaKOvjL1sc6bPk0ny+9ncSLbZeGieP7lGNPyN5j7cHh+OVr8
R0Op9aLHaSzrpIi7Dy3CYgjlKFDYKRpDVfLolfVKAS85CbIMH1ydFuD+B/JMvju2
5r4Qp3sbPFvKL4NgxdcHh8WEJgb6ilzudqX9gXrHXwkm2FAGtV1i1Nbs/KjdGpZI
1FMZ5pA8WRa1ZOtl2vcqGCQ06TyMkD+k+RWSgdIp8yacRuOsLq6WKFP/0ZKdH96H
F/sBe6WgdA+UmT4xQabe024ncYefnBaUckJz8pgtZldjNMXAphrO1qfD7cynO6xE
3CHkarbZunLKMWyulaXApw2DDd9By5tuUYcGXGGErTelm1z1ZLbB+HFfSpPsREYT
GTOHvgpCLEpvshvOV9lmojSq5X/UynUcvBLTSeAqJfdx+z4xuxNL0bIKXSStjrBC
Wt0SciHzOQ0w8bFr6SIBoKrHfz3Ak27aZeMHtklgoXdaq2BCXnSfWL8a+eLbK1cP
QpB8Wj/zJ9iH57tBH4Zt4GxMQQYeoS2xogCF6yuqU7C6nxj70SzzDh35mJzXN7tG
vAbcGtc9eKUIg3kDn6bmpp5AbW6Di1+wUsgaHRIoUUQqkldebhijf4RIr4KlZ1RT
nQ+1eI0F0SNOabnxgSmfBt+2UPAXMJ5BwHNtLrwTQjmUjnl1lNEs3zBCwmGIDQHi
MQd+Gnw4XgjN9ruSTrykWIIXi8CbbgAU7XWAf95lHDorNZbH8rF1LP/g+vKzLCfs
JtCYME7XYY5wnFfrvNf70fjpHMWqJ3jRvXNiko1uqPHEndDTJK6+1bnl4Zp1V21P
YqrqDJU+9ivAFwbJnPKXkp0sm59ljiqWldEHhy5fekEZXRvs8+F+dQpu5FkOyCZ+
UJUxkw3uMFsQ0D01TqcZUaDesOYTFOvjvv7Rg0OPDausntGaO6Gr3gBkytEV2iPo
Qr2SP24ublaN7obK4eqw0S8UbxZjs4KDAhVw4+ZpXUUSkJ1MYd7V78Yjvo/DSeFG
Sw3CsONqQ7N5MeswAvqqGU1uhPNt7JK3MaURdkeNFjF1nqJnUHQKTI+fQKvP1VIl
1R1zwkh7h6D/hgzA4EEqJBJZy58193cTdT/yIRnm1SLZCCy5qbFgi0FaZwjnNd7W
wmjfEY5j1m6KJUY9/MF73Pr64stPNNbrNN6MqZVO/gqtGePb3neses77tMaLjCPs
wdGXhly25MM57u2Wrfkv1Ecqkf79/RZMKjBC8+EjTFXj0iIhhkimCpf84pbMTUdW
3E2qMLt1fo8wO9Nmr+9MGPXQUk47yMHsJz5XAacUbCCxGmrGQ+e+Vv4pvnvNv5e3
feLEvrvG/O90smMvfGBrrXUVf3TzRiXdim1M++VLMrjknmUt6k6i/BqRb+q854Q0
+S1FJff16//GMwWXE4EVY2yPhEjLtiILR1uLqOwDct6qZGYUUaOogMLjQfaj9r2D
voynYu2ijKwwt+TIBi62MzA2k/HahwBkkA+rv9w4G+5W06x6CpxTLeB3APk3uGA6
KdBsUyHXXRNhJzrexgV7d3YERh7UlKBqjFh715XVJshKysyLCvei6TQQIEUgj6Jq
7aLPF9+p2tMmK1ppkSrV8sTXcuA5MmiTDpEolUBtFNki1Nd40M1D7sm46cpnWWxS
B6DzXXPRqOmgj6gq81aWbckdc4AMdfCOi0ELeC5VdcS34k0Imkgrd5oA7WIL566x
8zrjx8Sc5tXZTO8BErADiG3mPwwboP+IYospW2B25oRsbQQHkrLKlOpSY3GyMZSu
pKoEY6vZwVmW2Nx/dZt534/BpvJTmmiejO4am8ZwWF1R8Sp+4JTJYFgWsnS/GHvP
TcDYkYric2jEGwJ9LeTeiZEQbVdJPLAENRGGsl55qXWgS6G+sdx2ttVqHcULb3Fb
NTm066+TxHYAMSdzXp7EmAowbf3g5C/Zl930fYGxp5fb4YMGqh9AK1IKe9R0kixc
K20QOildFyIo8Q8+KZylnC9BjjHDwDcdB/xhh1UY1yWCzKKIwCee6ZSVXNkvImC5
OmLTJNEJAi5rUlBKEBKOVCkXyvEuORJIcHjz8LQy1/Vfcozf5RZqgeDJkk0z2FVG
oBUj7yx8l6Jp0EEz5UQ9I2IoEZgTiv654M5ffHCENUhUkoCXwK+LNgMTEbS+ZBAK
HlLrN5IG6zl9mF1ktodUOc05OS1nm+kdc275MXAQ3Y1pT5YWjwxFoCXrT92ZM28x
IH8iZ4R8KJem+bylRCjhOY1L4EdfMWs8Pti2o4biL0yWUv9wFuMotGQ7IuoV4nOP
9VgSKeJURZg4TQlNdPCzZttdkUe+hheYfUAdeGHGBVfYWqhc0aTJqa47fmGecZQb
6c8Kjebd7Wb9VbzRS5ITVxM1W6qpIixs/roRPPuab+wltoCF6LIGRg54sWvMpsGc
DtGa/cnMA2vFm734w7k3IkljF3RDDmgVOX7gTbMcp1DxT2Zv6JHVMSwc8tBlUG5o
pT+pc1ZBh0mtn+KMlKFBN1EYwEHEzagEIk1pO8mJJxSoWbai6sXszU9vaG664kFS
gRJOWyx2lRMe1J7227RJakI1QdTKqml3HZh3ZK5Dm6epSibJr2zosZG+YDPgX0PV
a5UzyN6UikPlXr8cDj1nA34qXVSbGO3Cldo7MUIG/C857cdWtyBjN08rdW74uUhI
QajLz4n1BMdEI3gHZMMD5+ZRBzP9bh3vv/uAmdkt+e8zW02z9wkIhs4K7uzpX1TR
yTOmNG9Ax1iJkJTRQtWW6u3Vh/SQy202jCXkyGR2CbieA66hcOmGIoHKRVeBtPQB
Hxt24Rf8seUMZdAYeklA3fbLTn+0q9fpUUeBhwaVC1FJ3OAF/raM26LBulfBgIuF
dbRFn9q71iIeECpnMmpCBCYyRayb6zL5PHOzod6Kwqd4ozkQr9qMWvS1UKKf1I55
cZYuWtCvH8ABzyqYiG0+zpKm6KAP5C74eTxQ1IhBy2F1y74CYAemsvPFX74Fl3Ks
jxM2DBC9jKAgMPhwrbpLJ5uRs89Q/mF+NWw9axxklxw1Ik+LzrPBwbkhhxD1sfuD
Su3Ncuz58xZcIJ/Tqw6GIWPLYyMIdqVSU8gVULzLVoK1czkiHuMPKm84VnS9HC3I
tr+1SIwRjU03TSHIyz0e0/wIm+eSx7uhp20rGCl8lzgBafTTkPXOK3EMdr9IC83i
H0rjngvrSbK/3rXvShF/0j1E4Sin0IA7z7bRu2UkWfeoCHPlB2P9BrxiNnXVVwaq
GM5arOkZF9Gb7TyF0atl4DyKrv1K7Mx39yr5dhG+KEFrymUuQbThV4oDlgHqXnJJ
CKPF7DrLrTUWOp/KYyEKj7S6Imlh9A06e4NpdDGl1zZaSCHrI1SWLMffRrlVONoF
McIaKHppnqmeakp7RbTBxc89peHSKolgxsLXShM/X4yZ3lJWdLwQ6hZzgKRMb+HB
Evw5M4At4pJ/rvcnAu0uv4/ZRaCapYZJuB9UPzhVAq91lJMzaGqzCSJkt6SYGO0m
2VOhySZSt6i6Gp0LVWhwky6HNG1E8R9srW3WNV54tKHiYa+m0ZRxzVOxzQvcxlxE
aTCeM31I4sajsxu9pdYLqPMPl3vsV/yHgj+Xm1SXljw+G3KaUTf9CGQdzNkoAUDV
xqvM3j+EJKboD2/F/a5aROWR3T1lsSd6mFW+FVG5D2IGF7oONnKqO3hSHgOEZ7lT
l1rdYHR6YOKaWn6C+ACwZR3nowZQoUapOUQ9xJPO8D1ofdz8kWKFU5eQxIG+VHTy
2k6Lf1S+ifeLmsfGSDleRulSuHGm2rHcFcNXnVBtlh4GRNMlj98O2IK+3qbdhiQz
Y0cQ8EQO6r7weE0uuywwwDqdXVG74PTaUJQKnfjR/H1JVYATWlu+x2qIsqx1hWX2
MnMLhVv7+Efs7TwJFvQ7+lRs4IObzYYurlW03O/bzX/prlfEQ5yrDgwZ0exhg18+
87UfWYEGXTZT1nPBVDt9cEajY0orWQVifu/fevDIFCLzGT+nyBXr3XSKNUt8QXno
eyQY/hrZt9gZCP31YxtWlbI2HJ1J8SGEGKUojzIzodV+8i9pzuXd0SoM12jvdrTn
SxbaqIhIMB8vScun+LStvD4scg8F0H7Dy1SGn3tPINQIQw3Uv0B1UVUj8QzJcgMW
TvnrgiYH0JWhYCl7vjiJ8+u5nDpcMApY1+vC1nXGeRRVCrNLGnJ1u/BIfqDXkCvd
FkyPmRhOac4BWEnbLXYrxp+DCpPky5jY5XP5T7qJ6gIP+nihLT47YYo2WcVEQuGt
o+x2//JdKxml4swDY+p0OJA7D6bPbNWMPKhZRXyYqWKGUg24o5bOO4fHOlvrNDUr
CvK5EssKckW73nAxrfmShX80sJzJ0kqkRboV94Hcl8i+GT9nsIQL2i9y57ecp5Gt
tuNACckfH4eU7BUujP37AQFvtzl2XXLej+VMBGTRGfbKPOEIVOj/XcGJHDAYb5rF
4oj/UxGCZJUgiJGkRehvzhga4nSTWwfUK+EBgyVROCpHeskSl/0RjwJjZsm8BGM4
vsdWchTVfZzU0lvIAnFsr7yisw/3GdACHT79S+wDUL03fBV51MhoxeZAKDCUfXWS
nzSCZU/NQm2U+bpRJdV+5lbep0984XtLcXMHp7LIUgycQR68e9/9MbqPKMruMEwu
vu8XNHoH+ftuOs08rSo9X1NWXjIutABamYeXyUPWLopl+k22zcceiVRXwHPrHlu+
H+4vOkW9MFXoE7eAnSRqp78se5A/N5ZzKe7+ynsU0/ca4ZVQqVqRLVQMWPHSrNKw
Wx+x0yFBUDXxGzBqDrRJM30j6oIlB8lTCd+L8bdrXFM+FXMnF7w1PZvJp6cFoHtN
7Bdm/a2ubl2kZYhaQz8XBjUwogPAPfaMBFkkkzwODgfsL7rzThXHvlHz5D7rlIUy
iR1DlXh5G4eMjKlrmvLTQlFI5VIUX3VbtugOYU19VtjvOJP13/lXkfVqbNLyyurU
pqlwCdQboGr4X8ZIvU3Gn+QPLZfcbtb6479NvRePydWlGTi3DAVw2/QSjYJc+6Li
OEHDHKLY53Tq7a3gIAtjKW8ROlPNC/+cKYrjDV48cugk9lLNL4YvxiaIfguPm8wJ
VfWDTI/8VXdaeaLViCZJJ9MvCqV0ybTFNlP9LkFs2detxn5buAU2XSUtDXBtR8Ax
iKwWfqIZHaOeOdgFEAxMoJQiRId2xQ3URDR5UaE5sm43Y/nZsySrATHVtgPSB3LW
WIAILgNRFlBuz+CplcG/5v6OXV36VsYOh4vmoBNr1IK7YRDpznNdCIetmT2UtAiZ
/K5pN2CyCiG5w6GtfsxeVo+zoUncCyJO2B1fKkwKTTmetkDKOkjW5/Pg0JzyqJKw
3l8SfMKgQVACdsed3nj3aq9tUJ87xjNlSwUtele/otCDlyHtRnvZM+ndrbRhTxHu
zLfOTMXMM2z2aXCHQzOq9lzoT4jVMc0XOdFqOA+uUjFXS+nhMT0av0W1HvTNpKq/
/s9kZQ66h7G7RYfqMv0Mbq7uMcw4C4M9VKLSaGqsW+2IoRXZW0VgFEg9B5zj+imp
+Zj+hUSaSVASg4RzX2i4TXTbgo3Gh8M/71Vxdh5iJ7PZn6Rplc3bhvLsPiOeVOv7
yJ1CfUBiH2iH6xeySAs3kFI7WsnQZMG2QkP9CtUnbeIQLkz8NN+TyQMyyuqOj4kL
X4y3swZgmPYs61/JaaluXb8EMumR+OnJEBbY9u6+JVJIVyZTCiffPRAu89ms/GnB
MRLMy7JaxORDZxzyoaKKM4f26HIoGCntt6S1LSy7woZP/1nMg1Fix/s16jqxelC6
x1LcQaTvXcA3+Mu1hwy65es6vpuEzPzcC5TgoRD9cHx2OM1VqB6/+SfBlyiOiWUA
sbEr0kfWxR3T+QC63G6XyxbpWUQkrJLC+XnuTlhaOaHkf/J/cIW01MgAxzYaPiVi
frCnsvVcnOpe3pI5juw23UVJM6fRJft+EbdKHFIGV+CzO4mHtk8xWlE1oWHYTnH/
TZxQdvGAVuBdpKUcT7F+llGPKwXH5IJ4MOHgrjPU92gyD08NW0jIvxAmSFe9SJkn
MPO2uOQqv4KZQeRYlSvb5q0Ik1h+2OpROKEwjJeLLRvl4Z8NueaFxA9yafiwcRZd
fBUgzJmVj5KTRCCifT6T6LzVJRlnyqxKzdXqq87HgJyWJSK/DASIvsS4S0eDRxv1
UOLngHdmNX4tzFwyFlZnzBMdQXwlZ21sq1jNIAlWJtk276BPtgomWPTwpuBuUZ6p
okCGP4mCyBbu7DC2k4n1gFQuzSMBzNNVgCfzsvUDFM914gNfqrlk4+PHmSE2axj4
Cn3eveh0E6w80KkevDCB1jZmOXidTIONMb1XeZ52/YUP1SvBgMU6ugj42sW0ZoKF
LAltE9erP6OKFo5/wxNU3FNTstjNwekEhSWuafzV3flOlj1gyKl2KfsX0BszvNiZ
0kSFEXDfg112U5TfGD34URlzoP0YAA3JZPG00DHa1STjzmJ9CYvLfoPWE6VoKuXf
b53LpD0BnURGGvZZ+uYGqjCHMnAA9dKQL2JW+fMhQUDIlGxtoigDsFP+hWNqQv0F
WM5DiI1BerO3FaltfFPJ+yljSGAHtQFj310uSedayOJg1clFa7d2q6aAD1vvk5Uh
HlF23MAnqqk/05zQiaZRMNc7JI4SF8+QouNt+d4pIcwdZrJPyEkI0FbWn9JDk6Xv
u3ExA5wZ/9/arwAZ0NqcjHsairxszTy3XwrxYOMmHluxLGfvT3motd+auwhKfIPT
6YCzqy2SRhtcAR8N3vhEPDkqP/U1cHthWwcKfpH5tnwmlKbarf9wwyAxdLhvrVhc
GPV8MPDwIMvU0LFV3S5rVpwYkxcQ0q0waXDR74tHnitfZ/TYIeRV+4aN5JRbzXas
k5dEZr4TXh+ae+efTTzmtxRfC3F9HublTY9+pIEeY/PpOULOB1GcYJ1RcBva4x+s
1lOC+V6OsJnTj6mNxNbuRWuOYARvSniR5SAuJNW2evHQUPEDRXN6Udp2cJ4z2j++
AKGQnosjOdEJY8unnBDdW9MLpnOlL3fzH2ktgX4/nmRM9OvS2OhA3Y6Nvot8ByQ+
L2I+sLJ51JM8CyywsZOJjrB/O8R156kUqkuh9giR2k0HgC/LEpf1bzj8KFfFvJWX
WOt7JKgfgye52VV1XffKPG2nciPkfC0VJr+Bt81yJeYLHv4sL4hs84YhHp0bGW5k
QP3GK93CbPLiNyEU3TWzABlwG3yJyVaO0ots0QbkIPMPOTls+xYyYkW5vwwrg3Cj
CX5C1ONqHxvrgES7iU7+PpUnF7ZsWlzN7jY64rRSzR87Tp+fzrcG3RaKnRlGeSXt
5FiN7zhsn2RoujmCysa50AXRM99/PDPz9e1sd6XE3IgaDAReGoyrr45y8WOr4aPm
TNWk8GCp+hF6c7NN5tH3uhrxMpFYI0I1TurSJqrpnzMpQeU65OQGXKG6X7nAZHBe
IgXF4AAs1h7hBmMVIY5GMslUcJbLRpdE1hz9qbi7t+5rboDqk74d36g0O1KVdn4d
VWw/G7v6/deZsAHPvMm/fkxfDwQLJwFFjFU6pR95yk1lR+igyGpsfrWG3zvESN9s
8ptBcsgEQyi6uDnHbUqVcGlGzGcBRUiG5myzGKADXjrUALY4QhheyWwG7AR7Urnh
cE4p8isqO42oUHI+KiyNbAd0lhD9ubwD+qIYxfCngxvklw2Cc/grO8QlSRBmSZOs
InIRUGTkW6gSSUI9rfUG+RzdQWt+BICs+685XJ9mYc6sYoSJOx3LIrM9YYx3uKJE
7W8xwCxk2GchoU9Mch+fikiWIIqdrWiUlfloPdjVJCZRv3VsI4/RNbOc/076586M
mzoV/j/rPqumHhnse/C0V3FhqyEIB6wu7Xm1ygjfr6vtXKwFwjK/w0IL8B4vrrMd
ck37z39PThA+Ird7t6xaNBdUg7ZUwzxDO/t469swtruk0yDXfw5gPULnBo0LFh7Q
7Id5ouAKAdIgx1dFHbNSb7Wqyidf/uQbmWSezvyi4kmRAt4ztecKqw99KOqvL0GO
++EMXuY3iikqkHkeY63J4Xgc5At8FgJTBK6Xq0fDRxVgr5+V0DlrSysrpVLUPPRh
Pp5QBpU0NXT4r0TodHFMTls/Y1/G9BuWpUaBdUcDAugJOPEsU+GUWhFjY8PPfjCB
UP8Zipl0Q+RKLPdEKpWakyIfOHBPGBkSK8MxFqeHV79aWn4Itz22ddy17qUvTN+9
S9Ow8wZ8EjYlnElNdQZr8iJcROIVB++jfT/0GPhTVTmX2Kkmmln73kS0Xrvh9LIq
kh6WQbqvKxQbTjVH3WPWZWXbv4THJmz6q9Ts2Hw0tNSkuESugdWQ42UkxL6J+gk7
eXVHpjwNIZr9NOeP4CVT5De1wKXnUleWu5s595mTLq/xp1xizAJivPqih7bl934M
VBbT/G1w7LsDpnVjxKPh/EZYUifYV0snkilhijMQCcjtMM9j2uYUuMOThCy7IT+w
P2IDGyTM1qMEOYzsbbNY79SZoXssQo2HFzNSFbYFgivEVni/SrtSNpihiVV1yJfv
fEBow4N9ovvDfCXtdXITc/iVlCE9Xj5atqfciSpQGry3+SxShWoHWKE5QzCfSK6v
xQVo9U0ZM5VQ0HCyeU7IiB34AT/DOfV56Wvz2fdWXgSFhNLN1+b6sB1Z2hAeIIuY
+kM2MsMZUbeao/NXoTT7KKWlN1Ca+7YjNLxoBuQr0bURMGg+kw66fP8oDMm4gMM+
4GrVSsH9+5zuDYcqsKS6rtBfw7Q4KS8jKbtpEVaaSinbcf5Kp291fGIRNJHRVq+9
dZqmwDfC+TcJTVS2GMhl0Ia7Yta7JM5MovGrte5Am0qN2JN1mkoWv23xO8J3eUei
lHQ/dH9Y6OA74SfDJuO5TF/KLf3LbQagXP5Vs01Qo3o2ZdU/vpc7an7MJhmDUdAD
x5KB3J9zp/bepXiZTH86blWUcsb+AEmo+CE3lOYvLrQbAA+bMypTUwxMYtexW0Qg
wOVqILvAFHJUluJw11gPItB44RM8lb3Sp+6HufYvFvCxvuDPj0J/ZgH/ElgeYYpn
jVb904eNmgpahlSOHEt3Nhx2vZBdbPRF4mhICtkYKWH1tXh5aIAJrA7HpawhyQhZ
5/XA0p4k6AveHGE9VOpaIiZV6ZdJxTtyPKFEG8xMmAoAXmzDd/pbkPqL13LeJql1
OP9SF9C38orXGSBAQt6wBKCJ01vQ88rOByM8IELlSq6RISVpYXhrcP15pM8eMjvu
tceE6v1mDVyrhrg8Xpyc6ugBTZfeCPYUHa39sSoQdoWE85bshtPxKBSqV98gub4f
TiMzb2Jq6LFY9a4K9SeKQQq3Ujqwl5uSA4XEZTEtZmebOzdCrAUT8m3YNxSEnc0f
PFkZXfasWEbyfJ4yYVrbW7FPgzGHVQd6REigEw1tntXrsJ2WdxbjpjhZFjU7em54
PpckiyLD/YeBYwSLQet9/PVBlY7eVuI/5LEYX4qma2oeRBx6BonZSiuQncgKYvil
MY1esper66FeuRqvhauOEnZSvs4ohN2ElPaw8YbyEosectJ/6tlvZRymmf1OXLyc
885YQc763hbx0dQcEWjBYsGcBoBMd6VUKPldrj40As/GlpMRj++P6NU8lerEmhSf
9y4lMY4w/HaZHxKXugoqFjPZkn+EOtyct5IxARQvZsTmVzKwlnE9aLuAKk057ip/
PmftPL39ahQixetk0+E5bp4dzadrQD6Dj1ep/X+64zo4Y3AeyMeY3Bssp3oUngmf
nkaExZfbdocLqT9e3nox63aRJcI6GocAeOzw6xMUfwTYddt0MOIeJe3KOVpGPhn+
xq+0umgg743FPMf4HV5Ec793RO7itMuwwWcd3x58WLGCE1FqdVRka3CuHZyAATZz
+4ijWdBB75OR9O04ITlfacCgAAw+t6fbghxv18K7fwmWIWL/NmDcQe41v2d2KvCM
uOR8elQ4s1tANwCjpAk4TPCfhsz8XKPRIoXrKF7/Yd4Bo1ktnmUajxgFacxVhirG
EBZ51O5RbbW1GgXv7e8tANPETW7UuT9oLH97B9xQsHGnQDoZsdkrnjRr4DNS2QAv
OVkgGD+hccxnF9r/mdnivKXw3zaQd5Pkq6v7/AOeLSY10MGqeaa0D2HTAXO2sVRN
muDLaOWdaSK+awVhy7XS4juWXkyOcayTk3f7lWIs7UrMPC/6X0WsxFw5wvdrbhfl
B21EdXLLnoQ9wJ/Pj61IpEM7dbImtpbUNHI+1EhMjgK6h9tg9xkhUjuBf/6yHHYk
17AN+CyGT+yspc83vsKkJjjxAODZoy8n5oegfW3uDgfe3MKD9UnCeAHo7xLvxtjG
irENVLoH+KjCVtiEAoRJA6zjTrN0WsXLBffRE9earLYf/xPIJHSmQLbGT/jqc7hb
5CWTYX6xGJPzBvSr7kctctawsKBifKpKwmLGVrQnMvYgDC/TcBkTncPz8yVNtoJp
A6ASoDGrJyZMKbQ+Z5Zkjpb5vi2X6T3snjoXBu5FMUkq8rFDwLdJylRlKTrho+9Q
2HVh0rKhZCwMuGLZRPCJlIBDJflFupuD1hXyyqg2pJJYjKEY4Kl4ZxwUslus/RYB
zMlG4Orr4jtFxf0I07ot9k2/c93jnRcXZGRjiuomVBja6au7vsOSRXnawyGrTI7g
bC9b057dJ2gJXgSSfLj+HDayUg82s1naCCgk0T2cBElWz9uGVchXEGCmI25SpB7m
69V1g38KxqcKcow60ioVbI2OzMrJ6UA/vSHEoiX0R+wrAw/6C3NFsZrT+xZDX3bQ
dBv6W2LNFfY6GVa2f0cCnGT51V6R1dOmUXRC8hmfNQs6HL1KGBsQOVqe3l5gQ/R8
+HJ1NlN/iouX+Kzq6vzLvE5cUxqIDWBEtdalO0xk9t7X7GauNZkS7HplcGn5u3MH
0C5p9WeYJ+hjuz2K4QJMVYkIWS63pHixfzsZUiN/A30NfcK0D//H0k3fMQd6dC4Z
wJllRUnMszlTcKxsIAUx+9Z1uhaQ0jVr93QlFLJJ40xcyzqGbcUYxzQ/Kvgt8ea5
bCKE+Yc54Qr1gDvfs3ku3BFq6c5+74zu2iIQrPJhIgISqCcEZaj9qUwtaPnud/AY
tViXyP4DO6cn7BhWwXMYAs9SU95N928wbgHW6jXv65Ub076FK4NI0yVQUsJO5Zxp
G5nAAhuXxiYFpLYJt/H4PBxUyJmUVXxElfoMkTYPddnQKmxOJ8tmIUJm+fjrfPGN
Oy3IRGMbXqPPGlHKHnE+B2tyKpux8w/8JKKPfYrbSwOuVQHeZljORZUNqcJOnSFu
qEbeCtIZ1NWEvV0VIw1sP5kGeCkei6UJ1//sU+UW1S3QHjc+gUXjdY3ic7RS0tRQ
`protect END_PROTECTED
