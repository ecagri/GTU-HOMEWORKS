`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DbRSn0xHo4P/8xpjZIaDlmr2NZ9IlCQ2v3jxZO5jQXLuZUQin1ft5gURLxx8uJbe
/saxzRAJykKwClWSEDzs7L3jDO0TNwK8SmVr2wGvKqI3j2Tls808ygc0jm1/5p9b
U8tNGHvpE6ymWUHs8zPBvlz4fyM7Edhbz5s7kvQ6ruNyWnuSkbt9CLCYFDPyyfyk
dTSMIw0mvYaoZgwThf3YWER+Ensw2c0aaK4rsOQXp8vewlUXauPUSw9+1eYzyGWo
WF2IE93HE+RebKJJ5TKLfJLsKuyUJ0PQu/3QRnCekUvXaVuGs+1EsBUbtlMxoWR8
UzU9tQPEz3Jwr+ifZp5nZLnKoWPFYir2I5ZdsU+Hwnv8rQizNdntWVVMRDa9A7Jn
wIgG6K5nCbck2F5+OPdrLQDFP+LYXch9ktzvftww6lH7gaJUTY1hRyvlMT6UZKTR
7M2gAwFJRoK2C4AW4HommQbKW3fuCAoQywgCU9bGaQWwN4EekGfIPFJlVXnOvo0/
bsDyrAXYpPkAVUlq5N/CPTJamsJeBhELxqOF3QKAcoG9uH4XuUWgNZMCL9zLN4EC
21l1xS1BC18QQrLDdiyX3vCt/d12i5JhQIciAtw3Tijv8cO1qkmINumDiMw0IZcB
OemtONrqgncPA3iKm523SIgxKiN53rmqQUvJ5jikueowQFMTXbt8wwSxrSYmMmko
5BUmIOIx2ZjT67fHGbjzY4/bXIi9/0xMBj4t09EkyHqHnJuBJU+UtWbyRy2bMCIo
j4DrkXlEPpi7ialMVhgXVyKQxtFYWI6GB9A2QCWeh1wiSzKyVTmn5r5xAJvfMFM7
pKAvVurE1NdHxjp1mMW5hly+JNjykPiF8jxGrhAHCJWihXgyh1+efuDqrzMUAZ89
lu+bZ8Xcau4GT4Gcl6KXC6aYvy5JXuH32LGAoP0nDMzx476O9LXXKHB/jJ96/Kfi
IexO9Tyhyr/mC65WaFpbLsUBrLoAai4LKt5yLo7ssW+s0udUAz61Iwjj1nAxrVwh
KMzlMcb5EVslrAYf2dcdgshuBGhQsShekU6Hjk5XIRvwQImZ5xcTSdb2zn6EumwL
EEh7iqMN2DmnE/0Mmhiow5nXtnDLBO27eCr+uO7Dj6hXFTc/dLPfzP013IQkoYvA
pXEU9CRlDLqC9u50TbnIlnDY6FeZqCaMcbNQiQIQk5M4mwdB9J8Qa4+FDTKA5hjK
zp1e0pBaxvvf0BZdLbI1iVsLFTGuWk3RwRtH5mOA8pDrXIwcf5lo1mMm5/A3X/rf
rs8Y7QJH0aF7n33vf4yoE1hGJKP455CXywcdG6tJrwQ/WKOAgfrMwfxuohtET332
mZTSb4+iWQdiIoSzTjkQUuPmn9SgjR1aK34oOTI1y90Cxf8xIRtJ3w3gW6L6Hh2K
7QTsVR47PJkkRdZN9t3ZgSKehK58FKJTHBQlkb/JmmkmdVZM/UgeeaK4RSAYfWy3
Cz62OhodA9dRIRjFXTOfJeaRw/RSTry6h5GbunnLKuOXxlPK/winksUJMhuTB52e
sM138Tz/IXZTkBMNHehLMKplY2cIvD/HMcXKJIbpWVi/t9gmM6Kzb5vtwuRi2N1z
qXPB+IQ1Pme2Md5QhecQom4mKdn0tzXRpEXO6M6k1iqXU5+YTr6WgXTdtjsvA6pp
22h1UTVvhN7+AsccPE2MyI1cR+OF31whAAka7PGBi0jtRgKlNWpLjTrgx0c6Ff7T
/cBsLTgZsd8384T6PFQs+JyzwA6MS5UX60Hh1221ZqHyq2PawYhmbQfOh8ZbntIU
5h3xGSrNHVHLci4yX6IDUUoYQmhAXFxAtl2hkv+DrCeaA/B5cAP0LvqWERHCv3HY
ng1zD1RoAQ/R2Zku9wH3YVftVruSwpl/QkD4QDEA21WHo6FrksH4QUZ3KNNwiYra
JsZsH/BKlKqY0MTi2QKMpJG2oCRfbVbj3Hg2jipsWb3A1Q/8vmLzAi3gUQ8aj34F
dL9bKBrk5TT+vW1llivgDM3gQp25oiImZ6ZCcS5V5NEDreFm/pK11PEUdUqbs4ZA
vqHXno+0EYpIv2uC4nbSW9f0ELijZrpGBxmuJMTfiXrlwBryFU3vEZOypg9ghSXj
s59IR/ryEBc/eQ4/byfuZBCR7r6b0FB0qbcoyoaMPpPGMmCqHj08O/u16JtEh1xS
ESELeFY3721AKtr0nsA7Z6S2cfd3IPUvf6gqbuEWnvOnRZdlyTVhvWx5gcLTXQfU
JF++K0/62Vt3P+pwolBMuiLjGKXfmHT7GuUKhroxRAyyvDccB8/j6QPmO9HlQeDr
aaWoaU6Vsl8w8jWvE2FNA3YrLHDs5m+2GiYgL59nCtYEmLBT+orQlCccfUx1GrqX
BmpELV+dJBQvxqbeo78qv+hb8kE67z0S/FJiWxNQfWvjJwE6IccqUIaw2cC6uWRd
OwY5xvEg2DjG6/g5AlOhL0FvqfFEe87PbTEJnE7SDsZnJdMTXcnnhlt6ITAdUtxb
JPSz3rqfH/xNJ0y16GrJ8FUbBhreNHiq66mCpdffXmmfosu3MwHaeslwB4tNRBIZ
+Xo2QZh5XfmW9ocz8WnMo39Gj5I/scSxFb+19CUQoxOjljlNjSMxUVq+9qlOvc10
sEbNIbkGEIvsTcoGFgpwBPs/qyBOcd7jf3+V/sx4HCOC3XsE+ImRRORVBZ/d8/aQ
U7xxccT7R5OTPDabuvdmtwehSpkklQFWKex1Es7UrMRWuAwJk/j3m5kJOI6J4sFQ
NCzl4coKf6Cizr0cBJWZGBRTaKjEZlVGqvk7fAOM5+AtJ23aNvM3XOkGCtgAxzlh
iZe8nI3nL592saOp2IlpkJf5mKqCYFfp3yqVT3Uo02iy/LiHfftFhhEJF28bm2z4
aGU7nydJluuQoJspOf/Vc7cTvUa8n7pWO+HhRpW8hW+WR+tttS5SA1wsKLNtQJSh
K2IKEhiz/dMJMMCDYqi3JfCjnCOG/0OO1P7tN/IVW2gZccCJpiXhcA/VE+uFL3ZE
fQa4aU7qPyFpuvFVl59VXbQEQTaUhlIT5yOOhnYJ2T0pxNofJlmRYxvKqHpnmVHd
/17p6g2TIkIQE5Jqpp4icosuaH75XYwa98AzDMP2y8r20AsXT/nOzNfv8aCXbxty
HLH07FlS3WmTmcAERomH8cee9oZ0luaG3PMJzt/enwofeHyLvoWlKAgTVo0THcs3
TslTHQMy5sNMWtjQc+cpMb0aixvm/V2IXS4aFiacmApPq+8yiaKn/E4hbwiXRWS3
laz0+hUEwKtl4uktxbUCLaGpL8BVlED5Ad4WvPflnu2YTvuQZNjFpV98cJL9wSsu
1j9tG7cTgF5UWwp/usmXcExH2woPH8gn+pOR9L3tI06Kn9X8hyXhDvla41kec+Gn
yb6BQW4/QQFozzhEQF1m/CW/l3nzsm8miAaCYWAXGNthfgq5YBeJf/vpiuaXsUS3
0ofX0RjDcVFAhErQiVKhOHWloYJVTLRpPYTSbBS8+8WHTC/Jk4bcslh+Y/Ey227n
vFrl2fk44mI6uZ69cf45qmbKvOvk0aYnjlkq/4ceSA52d2Vo099LOMa41oKiAe3H
yFkjkzkKQXxpqZOSq22LwyEcEbZ/4mp7xAUb/qcpI6tQT7YNm7l4ayVKy7rFpRlG
l8+H7ZEbYEyvtLe472iLTTyOF1wHxH+kkmL3iLgFPwbJ5P45317UmMqgF9j8HlBj
iRE9N2VCb0zT7tyQoz2ImRRfVuaYoJf03MoUIAJbnL7m4YTOxwu9nVHc6FoK/quJ
n9+Qhfm4RLJZ58fboHlDXfZpBUIWRp8Hhm6+mBOPhA8MBVwp45bDZQEUnP2o4YGU
c2Xod6hZKx7cQoo+eHcNK+ALO7RMYB5XOoYuqok8Fy4NBMX8wLQICatiazuijewb
gqS5xHZhbUJEZG7imxC9wvvEgWzbuA/lOTNL/rkg1jDuy59cm1muxiSvxvSJiEMO
tY5v0WgnLAEDplXR8C3AoKTjeduAqFsK8yolauODj9GPIVaze6zherbZElh3b1Mj
zCCW9LcHcqI2oIhbN2zB8YpDbCfZ5LEgU+8ZiWZW1fvurazMDuDQZYn0MX02Rhgj
BAmT6V2He0RMeW0SArETvWdqpKnGbnS7XTe1wv+mJuZyQWgTk8I6gOG7ZdjabluQ
VsILZjJpiejVdzQ7NbVeKKTnXqG0KvW54q32SC8GibfzAb98KX+GIESkOIlq+N70
xH5AhAguPaJzLq2qn8UiUbsKa6L7Xl27auX/ceuwPct63yySAHM7Jy6mi+2Jq/QZ
Y77SiBiQQv3TFMv69vfqlrvA3ZiBrZo1Nqb4q6+G0sNvgm2L7w8Y/5at84FPguld
9WlXWjkk7Ffpr9k02lTHZHeA7BFsqrbQOreSj3WOrijwEjojB+YQW6VAxdYKzH11
1iV06xBN2Ph/6zVzcDb1ZJSVzL6wfJZmNMFC6K/l/uwbNdRSD+o4HsdTOz5pvi3M
dzdMudDydhZNcigN13awCYiKhMfmFzWubtcLf2iLB//lmzR8DVKFQ55SpRH8H6ny
ReY24kWPEi7nWMZOt3H2XlBEKOYfkYzsL7lEjSdiiQOpq/KYSqPFnSy020Oqq6u3
mkOQskXwjoit6vmrPgyeCE1Dlpr/24iP5jqwnvKb9iLWc0x2pFd0bVqL3E2lf9Yc
K2xMj6knCNwDmI+LqM18C8rwb/uREK5dRadguvPliSPuTnw8UB7C9fyKI7It+mUi
+AlSfHBYkNFfSR50SXrqTDF1AuPOjv1rw/gP+RZcs95nMtwuOQZmWQRlUNlNF4wP
sjK7xQNxjpijQBrTtu1AWPuZfW3K/G4wecyUOgOqzxUw5pbewvwB2+jkmEbOGzj4
TkUHPmF69vXw18GSPUnXCNil3KH3Y8OYdFgvGC88KOHt31+PrJVhZ10PofGxlbPK
Bf8LJMtSY9hSxYUguPd56+RHu3v8aZ1QIYmED6tIFBkNhSORsN4XiXihWebLNrKe
1AkI8iHgBr01uWmWYL8Svbaia8pecLJ8gUWVD4SIj5nwXpY2bQCHZvVMFdHRmKSc
uycfBcRDJj6RCnw2eYVbk1rzqu9RI7UPo88AxcO660BNu3NQgHqD38dNACmMnFKH
kugH7Tlk5ZlJ7yQi71VSoDcJ2rptXMhT7oVknGXHqHtHB/ySBjgsBFGsmcluqLbq
Aw0BondoMa1HdHQehotrWxgY5eMJvmVD8FHcW1spTufqMxksR6Vyb3rI5NEnyol+
T8smzekM7MFB4yyUzsu8IfAozzs8VHuDVJyhcU4wrnC6uIG6q9p4uzmpRp+Max/j
FYCTNdQcCfZDVabmgdOQJojALaBNFnLnEo7WR/en6vOGuB4yuFh+tODkNsel9e73
ugIhbnd9ttfg/CGrRVtzPkEU38egjSm9N2CH6gFZkjFB7yLQxGGr8RznrAXrp8mF
VF5woDFet+r/TNQsrx60TS88zeJyeb6c6JVaoiNol+kRNVzfwT88Ln7cmAhwB7nH
DXIJaesukbzzTI7EVH0qjNOEypE9tlhSGLzhfngR5x4u1CcqqVq0ksMHGmW/Uzbl
pIBySeTyiB7aWVAmycpyLx2PP+cB3MklANhGI+JkkeQukb4wtu9QjoQGT6OOg/4R
Dv9/+1an5GNtT6mUnQosbFMt1WxsAI7DqEspznkUlQUESgP84qhVWSfjwTjeLjOc
FoTJyOhhqB/rZtqqMRNihpFnjpvqR9FkeoZOY7a9A58bkvUdzWxB8vcqp+PCBghw
jHDNBROVnNpMhkT8f3r4KE2ECaZe22F8sg5ecykdhH749is+FHgiSKkSfJ5nyVNW
omQeVaCcPsL35IBSVKyTBf8ywY1gc2S7FjRq7tKUQAk1AxXLZzAZkOV+MdCbvR3Q
aUQBn4fy62VHegl21ZE70CBtFh5nc1Ni/1PEjEB7laR5b/qJRHeiaav9gAPgaxeQ
PD9gurQKiRlyPc6wsdA10edyD6cMBr4lkPBj1w4gGsOBOPLk4n7y6HbNk1vamAMU
PzKIaFjOhR4DdZTzIhqhezaJAghHMuyCSrcssLc8kxtVkaMFtRowIjc+8GHQryL8
gOCmrh2Dvi/Rx82ybBT+gIcV9fmFABGdD4hO8+npqTpHm7vs1kYskPGLiMzy07lo
lzRHy5wr54ZMkKrqriHjapCCTqSf0Xr+zc1nGfr9bw1Jy7zMKx305dFCcY2NIMwM
Sb7euQb/0qxcwBGhKcLqjAGzYIWGl8wpmse29h1nixdSIgXfLwdgbYD/84L8j2+d
JQ6fSZa+0Sy11c6wnmpfXLZIUDpM20uJ09JJceCzNdZ7rEvJnAzw5oJ/2selx3AN
sgfdsIbn6cCkq1M8Hc60aPonknkZoMWYjm6AKupjrtxc2McguSYYjGcO3HPeL6Jn
ZNzOhOfMF9anvQqQSkCe/6h88cPKNEsX+MYlTPBauERWCuVDAUph9d+iBAxjkG6C
f2CxafR5qQqf2Rj0xFqvPw+vcpwZA/YRR7O0hL3oEKZhYULOitGgPpMIAOpH9YbR
mkBgvq5hPZhz2cdQnqAPEgyQNG7IlYnJMCUub3TmzvCGWhGdw0xiTE6fzS7ltbPB
+rCOg8lTDc4e7ceZbQIL3Ube7WoSzkDLx/tOOLsCwOWj9kAXW7CRM3fbRBjPWNrm
QMSs6DUIJYwQJ1TSPaCwwek1DHQtef/1IYzSJESshMXiZuDWyaSFRH/4BIaz9cRh
Gv8G2ZDkpwROOHyW7+aOtCdHHCbqO6wgUIdx82o5wPwx2Znyrz2756nHhfCc8kFA
s747VukiKGqujabBDCxxYHMzwUdDIkCGejzqgMT/bGlegA8N5qq/OAeLLFxCnqJh
bMvtt8342BI/9Lu3925V/7nVtd9wqBXdwfDVGSJo4chC50HW1frDNbDPmiwhEBly
u8kFIHrTxpCz9s1CNwU18Eqqg5rQWz1nqzZEO8l9Avf9fcZaYIvOZE3y6+GYnU4u
oEiimac+z9cWPZNOkZpeEnyi1MS47CxjJj1F1UD9XHHTaP9yFJD54rBTfKVhfMjS
7X5ujE1azp7hp3r6dRCo84TJw321GxxjsPX+AVvrTisx5qhuvnk8T4vMi3Syz33b
DFVctck+39enZo55wXOuYtPVW/8Keo3FuSuACMCvxor3rXJoYXpkTCXDE7/q+ITC
PT2eXm+c4WwvO9d1t8y3k36a1kRbvwMo+0XQXJ4EoaRFRqky7XFT0LzC4RzYAyNW
LTJHM4CPB+loNem6Cy0NfQetbTrSyfhUwh+uKfDKpew+HxRy7D6BWMajmrPEDmAi
m6j0hIcohEx4j1+HMSpGNbsa9gy2j70JbJujm/gHit9MH8pnhDOnM5vVCivGlhAI
ceTNsZ85cdmw7+fj5P/3uyRnm28NhSx/LY22Zb5yE4+MWu2zLPZDO6rGjr7trsqN
8qb9dYu36rF9O/ggKTgGsCIdQZyoMdBnheSCbGppdxABLLvqxKLNyvOtlXOxXhd9
CX0JnZFDlepbBcv9XIzRn028/zodB8wXoLVqxAviph4Qc8vib/0DUxhPisvuAQqv
7oytWFBh/qYacJv9k76YscOy58EeuZ7QSQcG/E+OokeUgheRCDdcimFY9GgzQ9iB
PAQaRRfWGVmYbJWtW5LE6yS8m3aENV12BuRuQuWfhwldj2DWC47unDR92Sl+GiME
5zUSKNxaFfmnk7sRL6HJqfrbvlxkJEnj0JuDBbjBB8nqLCDGSTITHC2qIQNct+x7
iAB5BJ8p+6qO+5lok/I7UME7y7JEbMDva7RFpYKv5LdI4Hq4oGoAJf/gmADSRpkK
tH8eVeOxhuvRGTq+wRpzmaKNQ1t/7pQoElxtydh7sQC4MDxJVSHCGizsqBI2Ndq1
e5VG1Tn2gb0bEH88ACmpr7tg8dFqnPg0rJckjzd6ZzOhagouzkJblYdQ9jpHL8Ec
6Qtd2q95SguBGzk606Guvv5/n/U8irEyGJ1dDDoRQYQNrr9wzevhoPN+83bjXplX
1cc/bGwe/wgkeGqKfG1X7GAN1NTcpOLpLNN3TXTV3Vom6tg+woyE8jVX49TF8Kqj
mmMA/M9XjPDQ1MAHZxhvtDzO8pxgtsZ2yx8CIcmYWmyypxujVm7vUPXcrAHvc6VR
aGd2iBPZERu/kSHxbN9a568+thOpC3Ptiz8qGXKwWXy9W7D7EjxSnPAVT+XpmND/
HD6ibpvW1jDUbZmUvJtkjyDz4swaBTMsvtzjSjcv88YyzyJMeCBsY/FqNOjgbd7+
YaqGfp28pfFixY7qiPxgWadR74WUbA4BIcgxwy04C4PxBAfNG0f2F0JS/zjPZjte
9ENdR9+bdHVJBIIH0ivHYyF83MpJWUQZn+uPTp9bhWbmXDIPC5DMEEHUBBdZwuEk
0eivTdBM/pd6k/I4/EGcm0Ie5Rlb/M3JnSLliYEHfwBQFZBSqQtgQEJ87qA1QXXI
P2cYwM/2kWatZqdGaENkbzLckK1ge5jOjdcvxnpjwogYA/bbsGGR12UlUHYgq/Xs
mtHE/nUzz+fvoqf+/38/8Tmxb1QrU51CJ/YJ2WTs3Qxl0ETN05D4WOqy1f3qz03w
CWmJht0P+BloxwiLElzluveFgV1KEfPqFQFMmikLrQQky1/dt3bMlh0hd2yI5nbx
lGrzdAITnOKzHUNRq6RQE6vLk7cAgzRyH/YxWTNhZ7dT5LdZKPofc2PrL9F8/U+b
ligrv5qqeXO2mWDAWqe4kUluoQIojx/epBptjH7zRL3XMFsROHouPNjvwkCc2rDH
j4eHGYTANZ09LAFuxwT3dJrOnGZSGlcBxsijLKy9FvjbP+Vn/UtsuwGXGBCb3mMT
qtn+mXUomWLVGWP0KJuPplEq+n1u46gfqJpTqX77NqMuiY1utojibrpdIfqwGS4v
mwpRjryLfL+ihPK4FEvOO+Vb0qa8gLuJUBhbGZRndaAP31bnEr6N64y+CJPzNYUg
5Cx0dgQS94arSmb/7SDIxx2CvIQ3CjdoqLHLowi85QA0ncAJl56X+fK08kjLHuR+
D27o8j4le3ibrKbG5OS6tbuL5VHyckAVMQAjgnMFfBZP3WAHGWP7RTJyFQR3SbYD
2OCm3MdZMe3C1nUfVPvqg/lmCjMA1wRkgMeYKwKvPIwjBbnQAOSNXJ7ycD+tJ5tT
lNFrOumiz+9uWlxQaVJNnhCB74BN3Nlw9M31HuXahCT/7yVkEsouDtnpeE2tvdm3
sQmrOGGx6SZBSorVYD1AaQZ1oPyr6LuX9I9CkVq08iuqIiRuIrko0ZWKc/IdlZAH
ZFoNftag9QcgT2Yrfe9JCo1i9Xem10b1QBBifcl8GaiZvCZOfbiIt9rcwrbIDwNs
SSZ0y5dZ2U+oaaSsc06nXsSNAPGpYvmC6CtdYFnBYiM9l6ct2Hp/mF3bsHpYO/fK
fdbqOsEFjUye0nkRz7fYn3wEYsbgXEDi5woG60v+XmuoBBUpDjyNQE0DvKC7eWSD
KKWIaZd9+yWFpI0+Z2yvKNQXRZ58OAIShDJDDbcdVk26LaN/QgTyg8oiUtmaBjDz
Dbuvc0+4kQ8EAf6KASddgKmva4Xn0c+di2pVR9MWP0hM6/BXA8ADcnqkF2R2htYC
sFYp7/lkVIW9ydTTvjRHjDxJhYi11j8yOGT9oKQB7UOn9vK/cUY2bdlw7Otn6QKZ
YSQ4ygMDsaHIyZ4q1yFQ1ME1qLjZWHqseCIfQ+JsT6GEvUskPBQvFUHGdav7zvqo
/MWM7bH1g6JqQu4Pynp7CLS4Qep2C9D82RKQ1i0+ExGnW4i1kIaf54E521HC+L+I
7CyLAVO4/kNJ+2suVQvkn/sY+AcLjHaaHXcI6iZQVvnyZhX13tn3eItz3pZtaHyf
zGhLTKkHx4SpRXRt7vfi6UiCA1E3NFLlqDV9zEbQKKjhqvGTE7b6M/3haQeDWPi7
sJdlUnSCGOUDCFjDaZX3UJRgkE8nsgQdXfil+Myc6w1EGYMbjIs4eE+km86Jf/1w
HWBsYGpv+NE7jXa6quugiAteRaMK9G6WQcW/shJvLbM1aAA8/UMup4Sh9HBrdoJa
q0IfE5K6Zqa8Ym5XjnuAaDX2daQ5p7dMdre5BW6Bu4XQrlPDbcjhOmojCt1ii24a
k+0+WxI3FXP1pq05RhEb5YXAJgpQwUIpFPxwueVvUK3jQk/qFSMmw7IxSo08PsKK
ddc7NUjoYAccotnm+BEBbFUV8lOENLNX+ztPXlIWSx+igB9oV15hsCmMLKZUb3Rg
/5qOlzoTbH5J6cGqqg1+b142La+GHAKvjWHqlyDkGskmyiHue7kn2/8hGQyRfp2u
VzLlFPQ+y/kqn0se71k+WU6WnzbkCENqKqwxh5rkrT5uWhJsajr6tAWmVfT/67aB
mMvqxEi6Rcp69YQx6aUxPzZtZWFBeVLtoo3N0F5kBmcEhjuRn5xntXDZqYQNmXF6
bCKajaZfdPTp8JNway9I3nSlblFWaBwWJkqQZHG5dDTDNz5oqqvMr+yz/qjvqYG6
di6zR1UdrMOOsbdDigEO+32zpoHMEcb7NkqBPOj0yLgh1temoW14MBFEUAqb9ONt
UNTG0hLqENjTz08BmIJnurBIhHDp1GjNkrNPGhj2p4afWIlPtRCnx5Jk96czo/vn
0LDwPk8SSY+tBd9W5rKItG8d9ovsEGKuFE3RD2AcizxguhGABb9LTU0iOrLgWiAG
kC80AbP13NNSrPZU7rFFHJ0+87C5aJn55AZnn7Wkk1Crds+aWczIBuyOjeiqzSDz
hzz02dfcskKb797ksr2t/FMSmmQQNo0jQZMcfeQEuY+jNHt84OfsYmtPHZfVU8+E
hbdMEpOtiZVbf+lfXBtfszJetzK0WjHzoToaKP+7aHBg5lrEWgDrXCGkCYI0SLiy
xAIG3EerJYuO1hSRGYH7FHtQRlzgJyrQzekQWFphn9zIwzbzxbfViQQOb1EbVMrx
O+oOAWeswRvzXgIMGuQnbJcsTlkvqX/vX+y3UoTcvumWj/zo+Zq9o1xd2/NJy5X+
FAlQ50+m8R/ITOH2v9TI3YswZAakwnVYrY1/ayyh8pMx2BAB8g1V3nc0xVxdHd3y
f66vkRqq8OgRr9sTpl8uH4BH7sFSIf4QqgVPYYDERs+G1/fGI9Gl8XPz5axYyl4d
3RqxyOLqip5i+BdUAooQKhe934dVRPddTO/gk/WerWgW+yJcU9FoL0mfD9GX24gz
WQS08Ox6ZRXwpl6NbaNuFWgnCxEvWU4WXdYV+sGsaTVCzN8qW/a8mAhhbTTdb1f1
PKVZ5hNLO4JXeyJ9+FpOHwgdQ6D25KvCmzgKQRDVQzA/WaMSlPyxiilKKsJehM8J
tHywLRxaZXoX/Bf7CSBj4JTroFrdwsL0JDno88TmJLay7g56r15cPpzKcfqctYtT
8svuiKv3QOfkEM/HI+K0tEvmuQBolvdKgv+OjVTT6iwW/24McfCcFYWSZjEBd/0D
124R5X5u5Z8QgF0aCMHX75s5RSPssBhs0iC+XVd4DWRjCd+ZEpsKnqefOzy+CxwY
lMLvLqS4ejFEouQ1pGk091wS2u5wPXrt0+P5/gfRBvo8OKyAsETb834PYnuDCdw0
2SoiEttll6LQiBNrR7Hl67KiVtsy/DfysPvp1cPMjZvsnZY63ZNtGFKjTTUoxXOP
IekgdRLvbOQODyTsEbg5FgydjlzgVkJ1/GM2PAutz+XwBGHxw/HY3PfZsOxKcoLJ
EJikEkJR7y0UnAxc3QA6SFriveLBPyxPzZaRVcZSQ4mnyujygzXCsebCgMlDUq4f
SSp/O7oBvyWH2LX1Wzql9QNNCSVGpmqKJivtoN1mjjRoz9YuOYrgoIVwm1XDqX9F
1uQh54Hdw3ft7BdM4Fsc1n6scHz9AsHmL7jYDNqO+i0LjOp/43ue0lIPExTY0ela
KYQKWg0O80aslp1R2fR0SgCvCd5E01R92KNpEmqEWGUF9BZJqni0dRHxAl1lhnvd
UsbRkxFvhmAwMooG5lithX/FMoQyrBMbt8ycOLbfClPAJY0lHME+kJ4MvOwmOBQc
PvfKDcKeWJ1NjOVTa69YNEsWAsHC6xjq2SX1uCeyko0owsDNiEVN+IUZ72Oz1FIf
IbR4prg6HnBrmHaJoReI4/IKQ2pr8jsEecrY4J1erIwkefBGcXfth+f27tOIMto2
wFGp1Kl1gHsbS4wx1xrdm/XkcTXEvR//Zt8q8zrTpSq9ihpdrOCMVn2AGwOYd5ml
sNrTZ0LH/cINumwVIBmpIsrti1WCOwUC+cMoVY12CcFJhLRIv/0WPTii9yZkiqvD
wpfzhGbbGn7M+Iek0dm7FW1Fdbv7n8NozrlBK1RYLmjzJhG7tIFp+aLotbUk9xoX
53p6W+RX/Su6dsH91J5i8PiJ3uWU45yx3Mjg5l28lxy8xIVdYCcrJvveVJoKGvAR
xhvza3ZyqbE36nWNVtIw5JzE/pCZxMzsvdtb04j6igB4MUQ+8oeB9edyeFzgWAOT
zSCjTB9t2Qmy/kDoryXVZFRDylu+vV1u61OIBQ2E3te8iWbEz/MDGsJ21jdXdExI
yHYrWZ4kaOYd9VWrigMY2TYNFX26YAHudYY4uIoqpKYlikFpnYz3H+nqfeH5HP5Q
nMPTRMZ76bR9GHBVqYAi5kyoDssomRq9YrKKL/MjOGxF1pS+zhEhd/UQBSFWrx39
r2Nicnq4bHA0GEr6DHVvaShxMi14pcad144eP3ShyxD+F1PIARPzXaXRH5Tsn1il
M2DkYdjyXRgA69h12yCPzPJklp9MMX7h0wtnedl6izGBgIh4McHvDUZQIOe9EIhz
s69ja3oW8qnWB/sCkPzJJWLPoB60qUO0Xy3LT94GCKBncHmQjsi6IdGhy55cpcYb
I0RaTVnWNeU9txnWLwkBJKb3anIWTLGGd1hc2fX2il5VNegl5QL93kKU59kzsIbd
9Z+KRbCT7hIV2q1+aTsianG+e5yyubSAUxvEbIwbXrKB9EiGu/0IpPzLbVoABvLF
T2oB+bUbXiEzUcCKZ4zaAScxw4P+1WY1OV+PILgRN3Ddb+OVwwxPU5eVWKP2s/fD
Ogtb7PYZ8C3pWwN+g85ryYrPRR6qyMou7ro2RzJRpYnhA+8kglAUZu+HgJX+K9rJ
4ukN9M3rELRoq8b91QxSXcpDY1VydyR0ywZRdEtHoFAvpHM1HPNOIpUnuCHOvCqM
6zW+r1sNKv7U/l+edFAEZfIfk/awPbp0S8mSFv2EHpQs8zI70+lcKb+KAeAwB/U7
cDiKgKYYQE96/8itf487WXqlbh+SSevNx33JvHBil7A8iqL8vOG4VIwd8F3GWSeb
gSxggu2Hoeo7DyzQJRaA2RLRy2pxNnCoAcZwDsmrOuQH3qXQDU0c6SH1KAPgLRbv
2sh1no5Dd9cQKdKotGyDUjz96Qapvqa2441lNAD7mjiCQgwk8FsdGTnor+AB5quL
UUizXb3OqxbOvkzsLyrwMC7sexApbqYPe7ykJU8tKsH0/ufsEkGmud8oOAWRukg+
DfUqtbo/4B4/OdYxXoqNxf7V1l3XEnmKGMeET4BoFWxh0jbgx+2v/3E/zNZbaKpP
v32V6esd5pHgnMlpWL1BPLoStY2sG26dtF9WJKL7gGYfWr+Byg0YoRmcc3BNy4OS
PHPnPgVt7pdyzoepGYv/yIHGTC4SMqF3seV+D3jq9CMfqkrzN1MX+eOgGk1I9rTk
a+++ohmWS6cgar50On0bUD8v67V4smjtHnpPt66PNoUtDQVoOOU7HTSQL7oArBkb
SkOlzi8HFWL+p5GUJ9SRunhjQWfUK8E+PEpc9YFFegOU7ieAFGTOnWSQXbhEC6Bd
/RmNhvDerz8tHXsbk/tdLPu//3f28BzAy61BNyTalrQBBqcpuYBrlqQWmOrENcZ1
0DKVSUpj1FHgIX43mv33DqZnOKD2QK86jYeVAwWJo5BW6t3YIGx8cYoRS6yVW2QP
Jo7I/t3XO4egWT2GXcpBvC+mzp3vT/9qmlxOnpc8bVu1guUtTCjYCDzfeeEqGD1h
uVIFRUFb4MEg/wZbu1d2YKoW3oMy7yjqMp7nxL+InNSDNcbMLjIII7i1zhEN/vTX
Eq8lRppCUAu8KVWh/27oRtIHj9otkNiX9FChwiV3GZLTLGmQqhHGqtP0p+DcxHxn
97adR4na+zjE+7fY128KoPCG/WXe87f3bCm/32d7E2jD/2OuZQ+l/k4zskSMCgPg
GSVbx2OYORE4eYTsk+LYJRaXqdR/J31rfRU4vX9h6DVghZj9ZyoV7NKnBselAnLP
lRTP4N2C5yJkamJEkPyq2BN7etQM321XBF+fefRTz+fk9iBvlFGctA1nVtktwqan
FwRkeCNqzbDHwMAfMWNqa6ahzVjtvmCJnXJwtWhF0lq05Q3J0As9yblIWHqXfgrd
6forXqci05md56dBJ1cZ8HEblhqZnKkkUDGcPweeCtjVfJa1kHhBK3d3hAtiiUv/
hTjVnK5SAxxbXHcw+gf8AkvpIvD/T1UnZdCTpBcpiiA2L/bpLaZjDJatLONVd7V8
vx2aT68p2/m9MeNFAPgoop3tFkZdh/maIOsMzppnnvHiHbPHDJLmrJXhNxaLwIDi
p2Wrdcdx8Q2pZfgpdm1YvSVMTCVPeRPk4Q/k90PrTt4XeCuzte2hEnaf8+AYcuCv
FEshQXzGbRpr/yRCx53GgOqva1SBjMhtWfQhd0OsivtOPQtb/HdPyV9PZzmZwEkg
sZooJehZ6VUPuSYTXojKqYbpFtksHZQQWw7+Q/SCn5dBfOT8cZ9jR3+bFZ7GqbdY
44n6nHExHpNueASJKOekMkk0Kspv3A8WqlZsfhFD/YshHU4VRfvCF4vgHuWpEdsg
XUPoi0cU9XHDxIvm0jCCjg==
`protect END_PROTECTED
