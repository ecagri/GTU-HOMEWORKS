`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+6ZJ1LiEsmhbxAANrFWIb/uWFSCpCRLo5Q9PKFEjKEHdte0zfYmWEerJvzd4ZkuK
fKtye2Bf4vp33fbQHRfimDlc4LbFZss59zGH9ECH8GG3ouEAWyN0ItQucwr6YLWT
vECHBEowvUOouytJ4qHIfGE/kH1o2EEdOdwGyG6e8OzUVg0lcdidIAJnwfiVAQay
ssM+4aqRwKdRyZgo0uFPVJA7u4LAIA43WcX4xM7XSyYI/R4pzuNZXhxGhu2M04Fw
pk5ivjCM7862rcB4zboqkuH3P3diXQ9uJTx59drkXvXFbHJ5ehSpf63/P0vKVcgy
sVQP+GqNtrYDvT8fDv7T1M++kIG0eItBqoic8vfNQ6C1IJY2Ln8lDq5nb0yi9g+Y
RvVrO9KhC4XjCiJUhwG2j5nou6aJRVmy2zd1hdZgZf4B098K3p0HSmnjn67GmRsJ
dv744kTbIeV1S8BYLcpIIyARExEQmpxRzU3i480vqLTvar5NprXsgLfjWJMQdJ3P
CS91E2DY5iWtL+aRa6+xou7YZgegbXJW+EWA9RN8JWu3/qKGHki6Oifds8Nd/2QX
5kHfXoqcYFxBG2RlAilhbDzP0taiDD2OETd8jrvFiNIVg/t629fM3DwuVAFuLSWf
aDCvkNzOegcbi5yrapngdiKCwwl9PfzC7Ib9LMTFs/KS38ZXZZUTMXrjQZl4RA+i
yr1zjYvqdDZluuz0MQFf6J+qIkPIGyRBMR5r1oamKiHWR27NPNZsxinPu2urV4rh
kBKgiRg1M4H557JGDPaDKTJWyhekBPIcwbpSwtw4ZCd3eNjk6s58W6VuQoL7y054
ZPebR5A86RclYmx9rlVm25nE7cl6jA0DOmKyXTnfLrTmzPrZlSwUYbV+hNGM+jkn
zh5D7hrNE2YiYocQPkNnsConsbKbm5XZh+8wEbP98npeIjAqk10PN+4GEI5Cm0Si
CVMBqHbfCMGOAtvzo66W5DwjTYb7jyUFV2dfETsi50Mb5fz74OKh+lttVSZ2hK3f
DAO5XOwXa7sGG+iR+b8FJ1FLjtZwNa5fZsW5m0qzvhFuGBlYvQa3Ql2RriMNiq5i
UYJ+wdMREOZqr9BlAVm2NNcAC0+D66UI4RbVspnkapTy7QqT/ZJbvb/Nbt4HXhIs
Lszfvx57mlylPWv0EnutzDVp/CHMw1m9l7fZ//WzTHnRjdXpCvcAqAmv4KRGIIFu
8hxO/OtVkdWGtnLwQjbA3r2JRNpW+QrZw9KVC+uPKEq6eCPG+Lgs6jq8EHgTz5Kb
wUg4mpJpjOhrFIz21n7Kho6Qk6JjY+uE3SvCIxiXEHcPYihBvVpwyCmo+F22ax/+
jygFE77pzo8QE+Dmbs88IsiKgnidrSvCmmECl+DEqU4l5Wnut3pmW6/HeJ5g/abK
W3fUarmOAdCwG4iEd0aFNCPUxAp2UCfDnzl6HzxriODLZ78Pll5ReQBOTwNjExZk
iDPJBVL4uOADErwetRHhTaLP/OkYwt/pBCZ4EsRgP24oBQ2+teSP9wp9RMJ7ZLmO
YrOIZH9yfxinFekqUu5IdhzUhQMgp1HU55vHDrQ0w/iVrMB2uaOuQ0zUrcDQtm+F
y9grJ8PnM0GXvOVHhRc0R0sbz0xqy1P3iPMlnf62iBc=
`protect END_PROTECTED
