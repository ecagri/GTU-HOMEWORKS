`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2PFq0rDeqRr8u/eP6T/YP3f0ISohJWRODuO7OK8GLTxo4RuO3gyOeNQqiTkJei9K
TbRSvty33WEOh3TWU3MS77mKCA0S3tx0/yUiFHrsB/1Pqex9vRzTO59bMBMH8eUp
iz8g5ugXN6opkFoYxqPYgaEW2cHSKl7+iuIeYVAM87s9F4mNLf+iapwGHFxK7w8Z
SGBXIpP1tj1ORn5faBTqzMeeM3mDY1ruFVfx0PoDV9q4iNIFEkqaJUDwdd1cPeW4
NgMm0UWprsU521pu4+2x7VHNrnZBUZFjoLV9kfowVlMJgpxOy0NRcXu9YUwCMxsm
7YkyCXvO939T4JRv8SA1/w0tYbTfb0XZ7Fty3Cv/jjUFw75oKqkTGyFjmgMkdvq5
QOaZ2fdkIdIzYG+cmEY7f1nK1cP6DYhKNwut2NnGwvX0ISOItVoTkhah7tEivcfC
VjKHNvyi89hVDnG9JLNtE+kbKK9Ze9nF6uDgbGeir9HTB6x+UlafGza+qfuIWYuL
0mxOhp/79z5K0eRqhjQOVjuppwtJz+WjqmOkRGGouby0dXGKEgzGg9pZT+2Livxg
y3EVAFPwkv+Ei9SKUh3yxZzf+OieFtRr1dcWtFvS7GCQXd0u92tvoOmpoVlv1TD6
wGAhWMy7bib3h2ygOIRpdzV/Ge7ImWEE8N6WUna0IwefLmIQycDUN8NdxCKBEULI
c+v7xWVsgmOV5OvE24Kt8K4CTxImFS2kY4RxQ5/EXnCk0RETAKeR2fKRyj2YrmkX
7D5qZFU21E40r1soZ9Qie6QNg7JxwpfGB02Xs9YC0v5bVRK9QfdIrbaQ50xZOCP5
V3uAtf70d4ORwI5yzqBfZEg6cuUgrXgap8/jaR8jeLZfJTB94rTXSiZdyUO1b0tx
bAYASMUcE4y9o6rkWOs+BhBDZC4NW4B/qJOJYz6JWoZl/uOEhvameEFZ2zaveSMu
u0HMSN8igeHKUzsQJcFuMvprGicZWCY5Lx9+pGyFihlIE6Y1QFYiL19caUn5jDLw
+wiYZNG0Fhp9bSkkVPB8y1CZAPb/S5U3WWB5OOVbWs1pLfuowWeD/VKjoST67A1l
nps3gVL8VuKYowq9bWOinijDY8IV9+qwoKeVpFzCNDswfuNjn8qlFoVwN/hAsRgr
gsR3BkOXPThZod9vq2bIA2NkHYhDd9/qXI8nHDoi4LwfhuFHhfDaGy3R3VGuO7eu
Ro+s3VMMVymutzTTh07uu5gGlPdt37hpEjCBhcFJNOx+6zOFvgeSnjmruo+KwmCL
OyIaUbjsNm9qPJ+yfYmnxTUd+vzaTGB6k8vG1RP29Me22+qNhZ5AuLA0cAn/IH/1
7h4VTFHxgh+lSvXni5VHpO15RNXxZ3884se+Og71vLRds8SvqzITjvCMx9TvvHXX
W9qn/NlOW6ZIRAm1bugvSjW2E+KRKEolLIW/K8GXzeDfs9thR8X+WDxpVJwAtDJI
CKUK6iUxTJdXIRY35vFmYQ==
`protect END_PROTECTED
