`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tjTfguMzEN3tkdH84h56BX1Q3anJ50uuLrCe5/w7Q8ng8ZGWGW2CK9IjgcZAQOTz
uGWAqwxW026iEenSAiD9HlMtsSqNKAB4JHE2cxZZL/TE7Ew+u9cpiq9Ma8owYU+a
6QstDswnhSLzYZG/vt3dV0so8FTjg91BqGn8ePk2AFNDfUAhYQJl86akwWhvJl2a
e0OdKWssbC+zl7GdTU0uHT+aCadOID91bOxWGmDJJAoSq3WTpSAZozgFoMaaDfyP
5KOMUXTOt25X/+Ytt63Ju6Ry7T/vvBvADS7OAHlydSZnmbvVGbvDunGsHNVsYB7e
cJ+rhnh1mzwnByG/xE1IFoIM1oQB0qH+Z+qhOHnVh1GJ2aYsQbSJlj1Zehu4aCt9
f2+xVxRi6p6cqdTmct721Q0YuPzx8wKXoTLecVeX2f49ssOUtv8IucEOTc4yObba
W2TQjgsABW/ZVa/3St2EAVaCOTNbQR7pYPMSeC9dELqZTSeGLIfvUaR2GLY2Bb0k
g9GWGbHLnGPmC6vwYJv+w3UO3God+xF/T0dIVTpbqzEDvpzA4LEM39V3DTZYtOIe
kny4vwsdx6GTwLkPEo/uaIWiYMjNHB9BhFQk4k97pBEwmNdd5NVmzi1gh0QYw7F0
6cNTKv4KAALD1C3Dl5Kx4P9MkNtAK+23n5MzaO2ecKvLOx5F42mxLc0k27Xlm8oL
OtRW21hlDTWzZU5/0FP+39C3YjB32665V5+tQN3v/h8Grbh9XlYiJ6HVJdal5bSx
kYYstWx7LWOlCLIFWnxWyQ==
`protect END_PROTECTED
