`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mp3fzrFOSaaE5/M0bnbaFvTwCvyIDENtpBuHm7pMeOlX7As+3zJtgnvy0G0db2XU
YAEkJtCgoo69b9gT1bKbUQDecLybj6u55bWEH+bo8qBd+Zk5HIQgHutXgpeaJ1uL
j1DtzB+TIZllAfPphQvdTQiQLTNuVImQ1uP5Sva+3MY0Neb0hzwkN8Fw/Ct6l7jv
4n0aq4bb7YNeVH0b2ibPhw+xgRBdNiBE6WXfI30hU08Zy8a42FxJ3iNanAwyq/w+
SYZOSs5EUVyUk/ADzMwEhcJA+BrejnOwmyjzE7xLiEL1OVYUfJtp8tLvLQ9KXnbs
HqyaWXyHFuEMRJ28s/WCXfVPfOEcange+9hidt2b/nU/PfRX4j5QSnmQhgpN71EY
1K+/4FpoAzsTwCA/y7M2Kiz+L5qzjl83PrQgBuO6llJ/eSCsrQjkCEfXWoTOaZJu
tfQNX25nX9+SKAcRoTTRdBAWh64cslxidmBaOnPZdCT52mcdg/mCNSRg5LhFCUqc
JwIRpS7xGm+GVqR86cilq2+Rplj+MOnTCcaf0aOegoKBhs0ojQExZmaKL/SMGWCt
G7u7G26V2Xt0T7eGVm8cNKoWyf8S3LZcGOaKNqiMDJay39TQ99xaYIcB/If4orrU
FlfVre6T/5C+z01TAOX3/XcfGehCuTbyw2+lFQ9zw0H/yu5Ec34CXoYGmC7s30Q9
6l+hj8fA7mXgojBNkJD88kQuO74OewQfGa5vsrvxL66QC8PB3xMWRJptKu8Btu0R
WjjOZ793l9RwJnojoK2S2LtRptw7dZ4k3QQMmXYyBIm88jEPCJ13UW08qlyDBDoM
`protect END_PROTECTED
