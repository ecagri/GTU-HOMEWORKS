`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5fd0Ln/D1sokALphlj97u99KGyPZO3jvtVRMNfmsaWGlW41nUvSEjvfguNZmRD1r
yjGmYYj+Hr5FzPItT0Jm6spbB04bx2CjDln63QVeJyXgHcvqmT/4wyl+BAtOjilv
YmTS0sqqFTlKxTtPMEFogUlGWbxfslcNlCkj6Fm439am+9tBd7u1JVqsXPfSj7V/
Xqy7bPiZWGmsZI1MHHARdk9WWRPnEqHJfGmXwLNNGEAYiK02rt0Zr/qHTnxz8X9H
gQYRCIKxVM1EbSTg/P/K8RvFfR/pXDGzWw2D9bs9pNJLq8Iv+boP4Y6qH37FEEUG
PSWq9OhFRufXlF2k3iiEoV7iCavum424gPDZ+fuBHsXYlVgMiErkYuadlUsnhXru
4vS+xAO2XTHqXxAxx21l01MOHs+FAZzH7yBQc+/JG9780KV1UcpfvztDnRbuuP4G
jjZtcxRZ9GdOjjhLwPt1DwyuGxNApoEtx5mDLwGh352I5ov76f1WaCPm4lyqqF3o
ixWdoRx5dOaeKggXhqJYYvgj2nJEns+nOxavSIa2HCp83pug6gYLsIpUjgSTHaEI
SXg6HyNtxD0p5VsYyiSwVMC8M2gFyhf964pEOSjCI+aV6CpGkOmyvqjiPJGuHqLv
aFxHrEZOYbfagxrhR8HFB1WhzeYYOfhyeZNml2ruqEkK/dcl7YmQmqe2vz64QKB/
A/ALJMAwaYDEqDTag78g1OEmg2FSVMsiOAQk8ChnxFFdzMcR9YEgWIiWKhqWHyKJ
VCoFZbdp3X0C23p4hRUsGtU/TkdZ+WnDCr7izaT+fGcdxH4ng3UBJnlbhsGWkzkK
9i0BMk0kaFD8OmhyyxbIPLK6Fv0DlkKCJa5LkXqWT+iYshZA+q3kfkC95/yu3HpR
Fcqg9chQrRR1wz+BidCy7685NWDkDtT9DNssxL3CdQPDOWBVOkp9p23oNCJxdxOn
B2PhqFXLv0inYocoEDbtYSWSe9APR9W1EYzEjUuQWlctvnuNhvpop24kEe16e09c
TtjzOjCQ7ezlUeZsDC1Fzx/PQ6btWzO3atMl4SDxqOIM0Y8huwS7oDUHCbJ3uxsh
T7/NGWA9D6b9ZLM1KeTA+iW+kT2Oet9YesuE8qhUnWDoZn5VvrkVaHlW1zMt5SSa
fDYR3RTaC9YxcWyS7StUQ2OcLO+ayntuFPYkARC1XUrPV4xTooJ2HnOlFuYkUd2d
bpREqr0xze+xKxUmI/hclw==
`protect END_PROTECTED
