`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5f3KzNI8ehOMu0iiH5DTMzDsXut/KBY7+sXnovT+oQd4nDO752ZyJaTWWiktuEBq
fGpUI7vcRaql1xB5/++dDlEHthTvo2t3FNw5sdiBL2X9j5HUJMf5OCnu+i/M6zAR
S+siRnArsfzgA/muTOuccxe9Q2VvUClFxZmRDE+yDCIFYA8B+lV+UMfJ7/R3LH+p
0HN4iI8xmrZnKGlMwQGJ8Exn1aeMh88Ze1ylQAjUObXp43+ODdtRv49p83tbA0JC
0QOFCO82JZJvz1XfHLL5qvFTXZTTBHfBorUvuXwmRZQsenemhvS5hWXxb2vDfKb+
qwTFuWnK6BVmSL2jLWTSAvyPF4NyLvsIrRUkoKJnvKOwm1IPNFnU3hiz+HK9P/w6
1utvNtBXZTSrbMq4o3uw0vEuZGcQjoRcAR7T3nzKL4fxdB2AYFBdKuT5w+lnCr+V
BhWbnSofDbF/avr1dJMbZJKbOcOpiA0Ae+/fsLAdE2ySpwVUfAiHbC1+tssSD/25
QwaSlzK0nTJa2Xf47Un0Jpzg/JrtsQ2TZp3JR7/CS7QIxg5b0Y2hz2mZpLmymJ03
QBTHMFjBPum04qfV4B00Xpxsd3gUnwpL3jtE7quEV8PU7xUGoSoX4CMxmFu/LKv8
hR6jQMxZ4yTaKSpJ4f9UO1WFZ5Fy8EFTyCxND8PMf2AhdxcGE4TIlOSxVnCvnr0o
fqe2ZciMNGuczz9OUsha3Rxeznj1XHKlYmxfaMP+b+EUOgmnD4KLzWJJoca+WtK/
++PxANi60aZ/3wbt1+hQx+NhJL/3mX6wtB/hAEwn3BAe2jVUoett0VIEw6d2Zaug
9VlD1MR/fCUgCLatK588eZ/ZCETdu5VdFTqSEy7RB9HQqodBkWHRRRNCtWIMhx2k
d/Xp0dbT6L+Z8aLs7zO57Isyb+KjrcihYgg08K998odAyFay7M9MgU00zKJh0Hk4
i6Fgd38+JHNkT4wKzu7qOBoUA1TNJkKwblVeK1O/1JTaKWIhdvJcZCeIugIaXJlT
HDK3/vd8hJ0Dy3MxCbw/by98aUYxZxi+HHHqrt2VEcdiCYLdkrlIYOivu6M/MW8n
KJHLibH6JEdx5WV5r77Nt/vsUiAhQHEPuotarK01Rhph/fYE6YP1LvrVoPCUXVlr
7QT/g130eWHrAlNv1Od+0QgeOsbf7n3Rz7aptphfyxTLua96IcCpGmblpbPt+mia
lFrKwkPBOO0FfuzltUUn58csgqa0vnKUnZSGN1wv0c3g+JnVf+JNVjCeiO+8lTS4
alGsNnV7ITHMouZwU1muJeKVcut3vfuR/rwX0CS+f5DgqWpc4edBsy4GTUldC/mh
2/3RmWW2G+t/benE9W5KGHcs4Z8mswOYxhYuwcUfDPoz10OEzGBXAcXft31wQ/jp
VEFF1OeIvUpCk8rMFqIxxAUHnwoVR0s1aNODirCh8/ToflqgpvlLxDAKhCBbkQtA
nAJOLRMWd7QvJ4MQQp4lHkjNY48iTNB4Q0V3vWMExl+1fYZP1jSKbKBKNBqBIxOZ
SxbmwkCvWpaCs8aQCltbirUdI9aX0BPZE0exz/Mc+XuALicWMue3tJnLJSMryYR3
o5KbIzSNxH/uRr3QFqMpCg==
`protect END_PROTECTED
