`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NxHyAB+1xLWiHBRDkmcurixhWRVuEqvHeOguMzw+4e4aOFBw/82UbUxPTRkb5iyg
yDkkMk2n+rlS0zKQseoh3EYB3tQYxb0enk/7q4qlDsNbytYvJlLCtDnGkO2SdkKX
VQWu7HScZtpp+B8MDHSqX3wjFUf4YJftUoay82cD+P5M93IzU01f7XW17AYkpF3u
oHcN5VHY3VC7Tao4n5YhvkXRc7kO170FM3BTb5NHUaTSdO1YwQJNFgcwaPIOuT6/
jOwTl8FV0SP2fqWs6/u7UtQviBIUnWZ/F38gmF6Ln7URC1n/lkB0gvLT1jqWAoE+
TB7VbxRRPcYeXeNAg+BmHXD3VuZeoldtfSwEehrKtuIabTUbcco5vFZe5NH9jFLM
s5PppgRSilP49ugvTdUzZuEm5vWfvCeYK1bvLaJ4MB+rWeMgmKRzugZnsoPXZDUr
4LOMqvG7vqy4aUR/8qxWSqfUDmDPdzkRQCY7Eq/jCxQwHa9SKEKd/65iXpGb4yfp
GAWz8R13QeqrBupgFCF/dAuJkfbbzl9WYPPi/Jz9BDW2jZPH72PiKzedSpOnJb1S
a0YgfTWzKPuiBw/m/JHpJJaf9gRENxhcKVQJun94LVjYwUFtrl4vSIsjhSUkxSgx
RtwR2NAFoiQxLfOnGc7VmVNI4LtkRMFxRJuqf2MiS2qsJNuv5cfEXQvMj1AHVTpG
tGtR43xd1WGrn0a9Ah55RWHh87iaLn3QWS15jrx5z4UYiSpyA1uCq8BOEXRUTBRC
KbjeBOfTwrWuG9SeEaPuJ3mR0j81dPOsSi7BIFLfadwE0BmkbfnHW9UnZ6iG6QAN
ukLYHPYEotRKj1js1UArLhdAsjXeAd7aE3hfVyGwq5gRGAn63/rFNRbD0hwkx43B
kc/Ls0weEJ2xKDg9E4eXD1dNLLUN3vWccgPquvXdK/+Lk8IIJxyZqt4bEqHlYDuj
OjIB1uM7vot1Yetev0AYTaeq7rRo9NAHa0eMXwDNupBnAMjdscQlu4ntksQ7eOMj
n/OHCB5SxUA0UFvM5xSDc1TgY+9j9rbDNGG1twNVIrHuigW+M/t0Wvkpr6IHbOyo
9tN+PL/CfkRSJmrHMASC2J1Ao6l+JXo/TLpWLdyFS6SYL3Dj5l8bHuIUCAW4vhQ2
zxXT7iOyfMOv3+pTx0wV/Maers+wq+dtFzM2Eh803Wfoq2s0jxHIuVjhuIYsRRjI
mVBgGWLAstDkIJmSPNG6xeKPJuHnL3SgU8SYtXMIryC0aIxR9OOt+4tu5C9ThfiG
wiLerj7gcJzEXownay38891Qw7kpVYiH/BCA8qCsDqoOwe9eAyrV9RK0wXVEcGMw
UKMqSnxG+EjNqFD4I9e7qyuyXoof9gxmwQGexeYlYNY7/J6WNC0Eewf41p51sSQg
6HW55Of33R0VcrbN0RLTTTYNW5ozcLiGAyP30s6MBN65uN4bDrqJJk+C7/YvxRaf
qa+NUuyw6iDJr4Vm6xDf19XEJx1uJ1XUs8hyD3jTXahW+WHDKApvypFnlXcQfVRt
Xrp2NIUzbic+bs0UowccRV5pOafRQtZ3vVasYTwTQCb82BvuGBNKCtMMK4R9wESO
CsrKaulFswgXpOySPrAAROfobmuZuOLF46308y6z/2JXxwlVME80NMDym/wYRFn6
LroBYtiWR8xeLYzxW4Oajr9NVIUvAcfCchetkHIX6UaNzX/3WdhzS+3gYtiDfETB
a+gIY+DdrRR3ofr/iDts+C/gE2rObb/1zU7umqImrAqox5ldop5HxktiEnElF1PT
qejLrRmdjQBo3jc4v/yZuTgeStIqc7Vi6PunqTD41x01hBOwtXAB1urCaoL2mWVW
azKozFTBr6BnfTZV2IvKpBKRD3moTnJxHW4Cd4LGAhH5G9zBU3uLXarIczpaaeM5
WZ3/4c+ttCt2CBMLtd50Ybqe7BGDlYt1y75G3kRQhlakgmFwfR4C7wxjHW6g2kvw
FbPDNZ+3iYD27Al8iraqvUwxWVkjNjqyG0BfWlP80zuHsfnFKddAId7ffBmkeejB
+feget46BJtWXzO5fgkqo95+bEZAkTE2BWEyEUPQCt9qlCSvHFGJFkGQDzRhv3Dc
RTw8ai41H8p1f3IK6bVbmpHY26ly7XjCoBzBFy0GXfgr2hqeQDD62+xzFyoW8DZ8
+41ba/BMvLcubn+mVanP4Yg2PypD9QyF1hvXo2PPFtl6EwliQWKJlrBLHkaD/rJ3
JjcyJ3W/OPgh0VF08qrCTAj4HtSeK53oQaFC+U1nud76Jy+8BQG8rxmoV9NXxWFe
kkHl3N7y2BiMlZ4RDgySfJc4VqdFyRWRmdmz5Js4UDr70igdTD3RUYZhtNiopKNs
fSPXLBeF1BsZ8+OfnYmfppv0mcz2S7FcICRWLf9uidS4S/OdoEoFZGQaZNWAdx5J
qDdwAP+cX4Gxzj6OUW2OQD8rwydJYf0D6gxy9pG8vnMGGs+gsiRzyNcHdDEhajRb
Htr8evYWwZ+nm6CaiPPIkg6qqvVwOMMRYZc6XJUfrwSclC8wVjQv9rxGgyKXJ1jM
/R6KhDtdeNhjTEQefk+95q5SsvqKZ778+vVOzehKjMn6HuhhU/Ftf5xlp/isNow6
CEq6tMBLymnsbi2USb2jlXCPAr4BkmfF1pS5uxWTwiuBRQOG90ldI2JdXnzZWylQ
VoKEEbyzQo0C+Y7eC6SQdVthQ56/e2LOcQQIIoKpOPvB0jXYotdj3rAk6Hg9uYB5
eaD9ab2VAPM54rccE6Nqygn6P9NsEoYYXa6UVK2tJ/SM5nc2e4Fr6FyCyXmTo80K
K57BAa497sV8i6g+N/xEEOkqll/mUg9VU7QkYb9j3FbXmey+WCTJt8qnT6bJa6OV
OH+KmT4qh7gICVcbbZj37OI5KNymh0b+IlHLJ7Q2P14ugVh1LWrwYa1Gz//BSJ/V
taqvmpds5zFbcaRO1aG0KkH9E9aRI/EyeFqsHJOZZBpiUJnRQspfM1U/t/CMfl+1
PkOk4pR6pprrNGJyTo4vDsXIMYykL/5F5+v0XB7frY4ihO0d0JDz5JlDxkHS7+G3
XEKTEFHLnM3fKktCJMPZ/z2HKYr7TYb+BRl16v/WgEt3WlBFgZau1qnKPNqmAa9Y
VcNejH7ewMsNW+ewq81Ga13HSpjC0We2IKaIs7emvkoVpQUU/xbl4HBtd+nMAVII
6D+4jyHK98X3qtB2SaZ6n2LbWHMjujlMaYR8RjnY3SgbEqXYc6eNw8R1HwhodX/i
WxIAPg8BQm5BIO/3GsAPQyB2RANE3UxXGW042PxltndF3oczT3OvqYKWJM163Q02
5BKbkGCvT8P+0HyQ/o56TzM5UEsCVavfJ5Hf/PFjuIk=
`protect END_PROTECTED
