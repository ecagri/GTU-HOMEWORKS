`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VXIQN5Tauyb1vBexG22P02QH6j3dN6KHDxU2tR3L5fK24ndg96Yo2228goTP3pD9
ZLRLJxe3bdYWo5o32PhUQqhDNnFBB/GxOMIaGFqyKfX2xQUj6hd8+xgMKS35wefG
QkBQ5wuRgHDbt5+ca0JeEpGTAuXqu7m/iZCBxjkcZgv5ctkYNddTmW1ihBZ6n4i+
oxwDA8YCFqo3xYeLPXKoC+8x1hP7uXscsePC0ECNagYtsxlGStOYWxz+ocAVwb6Q
vxmxmdTXiDA+Ps8ga9ZGbnAf5usAnCfZXbxp8XbjmJq8A50FUbgmI/r4sDpHkmL4
iuqNitYWt/fnBGB/IBLtj1mnHQclzh4zm73z3yW1hoBt2X0qcEEkacIYdqPyJE6K
yHpRAkbuKgFTzM7/weyEdu0wPziCCJ9uaj8G1NE48SNOCQkTaw+GwaZhbBiuZpwu
tVaUZW+wKnYc+Gpk1PcVy+Mhke02oxwUvLmJICPRvlFFxbPN9/Sp04H1t/4LNVND
46GuRYT8zqIHshx76JQ/HEV/k+CddlIWn2+8o3RRFPvW4RtVGjL8heFEOE9Otixr
myml7hQNKEgmC1cN2WDlGNOljXojSCwcHJIRKpuQYy6FhKCoHab6tNYGQF+XE/2s
KMl+L9aLo/FYQiFmWL8uyI+Ch/f5EgKOCGpmZDCrqpIxdKfSYq5THmFee5wblalK
yWw1CrQC/ww/dlgm92P0CkCa9APv8F0ZGgLKl+Ej0aksoNX51sm3ef3S0dZTASUP
OF0lWak0mcoXlXBxLijyDzMot+stG0avh22JO+Z5tVOpqUCxf3m0tiwr8D4wAQWY
YiXnybYScSyfjF/rPBwTwzwdxtX9rTS0F6Mkc0psG1tyoWXJQroGKiS/QiOJhq9T
tgsuiH0lFoTFy5IW1xhP1mhBnCEbwpmdrzVtXerzFpUbWBrYzJbbTnwrwIMn1Hrf
IkOTXU06pdhpB/kh1YtgzHo+GvOEMT9igYUaTlQwBleSW43T1L20xPj/yhYzrH0F
NlJlCsKa2nz8mLb2RU3olnqZpn4JN2SHNiMiw7AS9HerneSnX13kMFLJXBG3KCLL
Y5SLJxKgf1hIljvAy0k6NSJamP5c1ipLrMnoyt1fB3BNDVnVbgtDG2ui9nSH/1SI
3NceffD6U9Ob/IA+ygh8Cn8ocTVHxzDDq5bNCQ77xKIQKOVJSwwqx+VPDSF52YzL
ujDVWepUHph52cVi49MDwLFq0KFq2+X3VKcZZjEOyJ0IIMu83YpImuLtJquJh8cn
iZVN3vp2bnpjdmzD3vfVZ2UoHNlAHuz8Jz5TAUuw/sp5lY4zI9bIWWNCad6Uu++u
UyW/CboT/C+FuEPqDb+vQHwEfdQFXVyOmzf/jGYqyKcGjqqxJ/DYvJaDtLIqRGAq
ygVjgrgtB/qld5m52AVBuH9oxh4K+G6aClEZTT0+HAk/gRaZePpJhIbGk4Ex34AM
Esjov+m75LmFYQPWildMgImgiGiNOcFsS+gRhMjGhWZjx2jMpWP5pZ+UUlr2U4LJ
lt/dgia4pjSeieJFS0jxObAuq+fAY4auHPEJLdDcf3DpRyGi4hwXXIpI70LRgrgs
k5y9qn+y564qd/UEk1pyjY0HgZak4TljhebhtyG5tVXfFWMTiNl5FUUnCrZxr1nN
JrTvg5RzPaCgUOx/XaMRksI4Sx6kT52ibXZCXqu75t4cZ1ExxCyhLOxcLmftf+x6
cNEjMITgfhtFAmubLZxNsugKJoj/Q2UNYEf68Jrz40cadY6aQIm9DL7TMZkASAdM
130Q/xJbFuhGkxt7ERsaTFfTH05vzw4dz/vXYO+8wkT4gtY7TP3D2XwavSwl0mn/
AS86G+G7MwtFZ9QQ/N7g+0434/xHmAjHPoGXmKULZ3RN4dG2d5lPke2RIl2nsuZH
GWk4W5g/w5EW8ciXLCS8BI/Hs1hYn/X9HlJAPc2X7bfIRQkEhjf9uIZ9oZzu9xdw
uikZUk4qTQiBHDW+/IlCFShgM37CpQ+TLX6ZJaO5z3ZA84MG2W46Dgmfhgv/wT5U
wKsjPyC5lwdZHrolqiIq52MI7dYtIRTO2gdy69eCtj/regxP5fzprqR+2wQng2MT
YEZrZqp1h7hufYHiUaRjlWHkyvbeCrZvrF8MsiHKSEzUy0ls/0yWYYaNNVG2FaUD
2vwAcQ0khYH4AE94vVglud1jbOgDzI3UPojZd14rQIJFdE6gqu6hcthK7c23QhIj
qp5UG5xlDq6CW5U7gK0CS/o5Pl/U4cmGk1OHxMEjXbCfhiEBl+DgMBHM6+HuZFP0
UjQgrrUUqA49NRyurAu9FxYWneDgDwxv1v/Ljv1BIbFYQvyQjU1gEMgeJSdPJawS
xbWgbbJAGf3slwIp5Er+ec2sPU8pChVolGuDAz59DR56yIAsWAHv4jAqUBiPgoJf
VNr5qz3U6NZ4rgu5MUCoETeCR00OCinGYzXffOOCRzt+QWAbIH+8H6LXElLJ0JIt
H3LHs0PcJl3omxk+VJv1XDrOglrXbGY1h9Qo6L7NrvhYmixJrieSzo3ue7Pli8fW
QClEWMX1HCDwEYnJ7Nuf3QhljflxiMksa8XDYGOCcDF03wG8gqVE4v880PeBFmYu
IbUzbumS4P0XcktTuVjbCiMcSqricBUpS4EijgN8NybXNE8EC2LCj9z7HayZJUmd
amfZtpvVvkIjbwoMSZi1vAFsV8hwAwH7lwn5jZk6FNCRTPUnP3kP6DI9+mf6Hhc3
k9FzW+g0L+gkLUCOFYfPMrb5Ichq+xRuVKS+N2iwOdmhgXSnhxiZ5nxwMoHalUq+
/YN1ca/i6BHV7G1N6qBa5QZ1Z1d9t3Lumvs/II1aoEvtQlsw+ZcuIfXlyX6LPXWL
xMKmFYjp6TOvxDRlfBofCJRQjtCLNaOmJJ2IVSa/a0a3OVhDOVgXJDj7f4F+fVZU
aTCgg/Man3hp1iTLB+j69Y4ls5rPJsJ0juzmzFmR53vgt9WnDYd+KcraBH5oG5GP
c0RmA85N0WiprKu2UvZewdCXQbGM7LCG96zafDc1JgUX4CgoNFIbDGKDAz+W4UcH
kf1CuAytJbn9LVef3IhQiS2yGXsnYNpleFPn77fLNKMaxXnb26smTjtRlhwiRcKC
7ALj/50zl91XHF73Ta2hxhnGJbCjQX4V3MXQr2htNSwjh6XOxhHhTCHIe+Q9tvDX
hz5Vtv4nkStzPUzAu+NiX7DRMJkyreZ4CBtwm8Wbew4nuHe0cBk9YOV153PKsZhs
g79c7luBslqTtPc3AsNripwb9AUqm86MZ/86OssH2wBiRs6KtihvxuYCI55zhdrn
xKyAYCtpKZ8Y8gsZwYhfyVGgdX7/r4nDdoiSmeFwpRaX3Ut+ueKVevT33txQbSl/
A0OyZvgAU5hjMQ9pRg6xnBYbVoxj2CbO5dHI6VDwICzQxVGcmz5e5BkGEvI/V85R
/wYFz4etPf0sL9qIPa0R+yCFR2ZvSo0dN3d7lwj2f+C2MdSGJM0aVAofbWrqKoLF
2v6MaM87kJzLTfwm7aa9Jxuzy88k3Sp7MCGZX6ZG9FE84ocYcuMGITrkOnns+mTn
4k1BEgYEJOBWxe+gE1VP47QrQbLPUvecgVysJBRiK57D8wCz/clQcc9XtyI1Adef
gN4qCBywyzLro74rKrlA1B0i77nOPYdZIuefaokLVJZrY0bEPCoq1LTPxCcdbDBf
oHenAWy69kEOqcgJxi2jxr5CyyXf2Yiivk2CdXTqOtZa7uzLfw07pBHC3f/2bZMG
SyzkpSIRA6b+vXEUFuS0B57lvwrdIxxO6myWlAaJyrlMtRL+a9v+5A4Q/ADuAPxa
4+gayivD+uBNbuUJpzRAHg+QrAwRm5o9LtKvNf54kz0MD9fNyW3AGnhn9jOoKPC5
pFEbEgPQv6reBwKICs0w1PtbSkhmEi7ib46pMQLw6TDYbFyOZtI3XMRv7z6oNATj
RipFUhrDFSxrTupVPBJM05tn8l8wGMDmnLx/ze+lzeb5DGbNElsl0GyR2o97dzYY
bHBSBxdALqHix3aTAZwEk9+wSpz4Ylgb3JPT7qfcfqLmX4Xncfmm5bhAWO7MhLw9
zG8ayn1Ns6sstRVxoSj6e5YnQQtLIahmUppCt6lOsFyJTzTtWq/kMagK2RsnpE5s
Q7vbshaV1D/H3YcvhjX8XRHsgE7JVYjOCANFQMmgeWPE93OyJ/32ujdsQKMFqg78
f6Ho73YeClwl6dLoaJa8o79EO0xNOpfLhOBagNkjtJuIBJtRTTb0qdX9TR9qkA25
n2L9HqKLy7/KrgNkDE3MUDeinh1hMJDI0VPlkTTFzFDReGPdVH0TgkBP37s2Ktii
gefzw5LyBWqJBMugOcimvIC2DiyrmEdOy6ceAqiq4jRrDvU7ljwiHz3Ct6vxYCg5
P3m/kKnp6ZPUrn4LJ+TF5agun96dyGFTg5Xp86/XLAL1YMCI39W1F0+/JUcUtD4c
hAnJXVpkomgDTf0/pRFClY8syx2dCqjkoaUt5Y4oYOfXZTGeRFFm/sKF7WfL2ADJ
ECNp25QShEETJu+fEhDT9jqWUx1oD5QQ78AlA1NEEAiP2qklnSktJqzh4XE97thp
OnkD0tTcD6D88N4NogmfCeZGgQHwuJESny9JlhKBfS64tHEWq4DDqYT3kY3GKetN
hb106ZT8MxXz8Nc8oKXJP2BObkYqiqNBN8zvgqu+LT1sad/6eAWyBhl8hlycRF+r
7iPQwfv6S87YAdlaou27UxhP41RLqzcG6dt22QE422wxVri2ZaCv0Xbg20hRmsiq
iaqtMqwv+vLoofGzIeRnDXqk0swJR//gdTAtwDWe//EaCBvEEjCleEOcU1DMHgV3
r4wKGTCx8hI+KjI8kt2W+uddWZa8M3lPjY8odtcrijZm2oPR7SllWo7GC4pro/Q+
FjyyzR+AELt9SYAfZaMOzEfhymnikBvSJMJzo6C/1qNgLYGEnJfpu0xaVJv9nVXI
1AVOELGKuIp8z9WXtNiq96/+xfaViscZXSi8CJ4NB3ZXoi3mSI14YDboMU/ME+e3
I0ugn6jWRRkZj7QB3CE38eu7jVE4L7aFW5QAvEVWTKn8/rXvB80E8QruFquecv2M
ZX4+c1qkCTJ4L4Vb04HAOzZflysB1Ph6XhG/iSZs2Ha1hVsJtcZE09ZP1V/VEJ+h
PzNiyWLl0p8Dbutj07WhP1yfqVxcm6Oy8MQ5Hd0lmb5C0cGFJVLC8NCixcKg4Fgr
xoPU24rrZPDaMMv1kG2yuKaeJNgWrqwzn+FJGG5EEPgn3YTylOSvcYFL2em10h1q
bXcXh/zr4U29dBGh/Q32Bl1JgWmfk8Z6fapVYDq7jLFXstj+o3D2EVCrmDJss+1S
yawDXRNXZDCdjJV3Y6y5mFP/r2Ue7OPDgpsO17f5SrtpHUtciV1RG986J1mdHP3x
QBM525V9lp62/83qn7OqZGDv+vx9Fd4EeJPpL+0DbS+XUsG40xWzikPPI4tRm3oe
dPii4XVYA+97m5aV54I2qpUt50cnpe0JRc8U60nbP9J9r+Bz53XM3c5uAp8j0HU+
QddD129m6VFOPpwmye7N8Dv+iPxwW/3E/Cozln7bvk3F2PVl4lJiWCIyccvLOH2Y
yfMeKmAaGLvhUOZI5eGAour9rTY8nhReBml4MCBvFpxsTuXuBMtxIeNcc5y74jld
Ojq8R42u8OhJEasBfb+f6lMqzJuZ2QFkOxESreLQn99Tn7feQ784K9bgHXUvSGun
bix4xwMmdo4eJ1stmKI1wuRC4/js0sadtwCg2237RZU+dc295QB/1CMWzybU3LSd
1jD5BHIhdZtaGI5ADGwdX+ys4sftbXoYkhnsFcrHHuR7CMVCO3/g9zDIUuWjz4gb
dKYnbxn7S1o+xNidI/NGfPNGpZNzcIOXbjOrF1KTh1nAJo5/uU2DcQ9lPs74xGZJ
rJBPPinxq2lQQlfcKv8d69qfU6TLGchXQRyBBfa6hmU=
`protect END_PROTECTED
