`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hjisShj8h263WW9LbYxOOZUDob4QETQDg2Edb22jPP+UrFF3BbQiDONdIOGQwJFG
u5TBGlpPhr0x4Sy81HqEbY/s7/QRiWm+MXzZsgwQuF0m6Xg1iUkgVCjiBVMvHPzB
C/qk8AYwwmItxFdbUq3uWKyJAXZBtVuVBCq/v3NhO3sT4UVMoYtTU9iNuIYrRQaa
tMsOer9ZzGucRXTqs4k81abw/cxrRoBWZvjtJ/kfcHbgnEr/jqBlBk7A5B3A5nHs
ZUTLnrxMuB1/dOm3mDU7UxJGmRpVDk4vHuMqhgsa+V3ugtBr4kTN4XBgKs7RRAK4
LjcxlscC+N0dXIcNXPsClRaBTBwZR+t2IiXgU2c9jM+j5lHbAvRAq2ZxBr79MluV
P5d6LZIjLXpC/KTEiJug2Swszk3ZNJdfwthyP3Hl5hvngiInfNsOPODxI4m0X1+e
hlQ9oDKMMLejzpcKp4RcT8nwIe052jHa3/XI2Z1gAHIrQ/BV0+twMBFgU4l2Mv4h
LW4nQ14g2PVeeByvzqBfZm0JhvVDjQvPjIrpAAKO4xTtFzrhJf6siabsLw3Sb17Y
lGdp4mLiS0U/rOLj+U9tVAOl7E0nuRzkmlFP2Z/uhJBC6nVUTFOKNQQLWJAcIl5r
zjRjjITlQQPE3Ch7AtXyHY/uaoh3JA9KyETrWJLwt1o5XyGxE1tCbEL2wxTVBa/o
K4NGHMc9vNhX8E3CGUQVI+zQfZRN4RMoDshaUcXPo4t4THmFvavtJsKnE8yKwRs4
+WaEvvfWiBwgCPxxDlyqvAtrmPygsyCSeHRmi5w3BQCmHQll97ff2NJU5s5NThKw
lT6o39m0YY7UXr0fRyLuro9NOdGKZjj7etfzgOQLFuDPyxjd3OQ7j+1FLplV0dYa
pCvIoO++bjhwS0ngSbo20yi9g2iRISUSmATI/H5oAiWhtzLz//dNYv2oiC/SRZIj
I/+hx3Ce2ROhdR3iVLH+pLS6cxlMML9REw8j6XGACnpV5BD4pwVMM14YbrmrXNQG
8b2pbnIc5WBIgnmkF5/T4ob3SbyovwZdqtBmbIQETrr0OsSvcB6/d4A7Js0VlBSy
7Tajuxa1SSdJmDxs6dkvvrakBL+YzBDfgEioONgZxLqvsKLY3GBIvD7Rg7dkV6wb
z0iB7hZkeVoWDJLtiTxreBt2ZfoHnxNKEQ7NJDJhDidS9UHpCET6bWIpKJMUuNbz
tBYDqJyjrSF4xwLe9Ioehgfq1nNKwsBo3Qi2b2sDLAV09iciGQ2ota35RkIhC7s8
F6cMi0XUGy9ikAUAR8VjmGUOHjK628C7XiJ8AnOgplojgRl8jVySxUTZ7gvGqp+0
p+kNauQ9C0FOO35Pzej03NObWtEh3Awa1l4ZXk5539B/XNfd0FEukLj/1auyjp12
yyBqxo/PO0nBxwXK3LFWtbKQvLwdjhWawZZiiKm62pZyhPMfP/OZLdahuJneHrZI
iD3obLocRGerg6mRl8GghbZo9+Y1jumXROT1JzdDYyHXG/g9fRVoC4rvBE7jO5zn
oy5xN9WMhWDya2vJoDuE+2/ZmwlIhNmobyiZhnbjNQbfzcmLv11yl9Fr/oQHgM75
p85fSBNeEffgVB0PzXNzVGPtugCVHNW90SPOmcYkppcgdxkC0LxMX+GSxxZLxxyv
Mnj/81PHTInJeoSeO3enGNrHaDFMHNsVlEyFChibP4JsALblxoNoKaow8HndY4tF
1e5uC+HS5EZxwD/bWeDHA0ZFuK+VeOTSUL3gh9TMW3BOokP6v1xauhx+riBH2nkt
/pnBQ22ZLpjP5KsBJXaoAjh+6teZLp/O9Bi8Ydga2WpIqK2Zz8FgdXc29DikDftJ
3NMN22CS+HC3MFzgl8sS+i6wT3bIJEk3M4FOrDOzvqytH1IsJybBvGGpxkZvgkBp
4sYh/zpoUNS5fkr+iB21pbhaqU4ZnuOXsoHfEbsKeKrvNgxsJyHF3Xsbz4vdbkpT
9rpXAxPuNAQ98f5rwtotRWNIZXdi8ievQVz215rSAa5BtVLDoJETVAk5HLHdBVur
qsXbniGHsm8mo2qry1kGLXsWzs3W/FUgnH+b7f2yE5OLmoLGpHg7pfy/LcEAGaW/
qazwDwGCl638jcBeXsaE7BgeWEx8Ne/PjTUdLif0Io0qW7a7Sb5wzHUdnWsg81Y5
PVtmPgNlQK6TTck8xUXP0NjSDu2HbP8LhXRPtSQvwOOxEeJMIg4iqutFJj7KkBy5
BNu+bF/uZ+ATpUbAKWjI/5RBP+mj7w4Cv8ycgA+rSPIDouvS/sLy9hZqmqYmZGYw
VW5cY94ePaQLA441vC3d8LDaV78kSZSCTNs+Ez+bYMra473wsym4gEn/q3sgNF3M
H1/i9Jl+eBg9DM1ut5x3DBdO0G+Bui+zNFE35Xm3L0qMs5dRhzNwq70uFVCwQUgd
DyWsiSHCw0ChR43Fe0ZmN7t0iD9VTHtKidQk5rxtlsp9qY0q5veQvFg/0uNIpg8q
FM5Fl8wP+AHxGjKSOLYLB4BPS/iQnBu2vQq5/NEg3FCQ6rNoeY7AkIeMZkNZem7M
XEhR3A0+aUtAADZOO93C1TXecSJRzjg8etBzXxv1w6ZqTgH7ChqmdmDtBxr5Z291
fLlWGSelw5SzfJJgBPAJfKdEhTj6Quup52VqoWcrlQDHqaP8LiZ9EY7evNP+hH7w
wfPNmSPzkWpwHdAqzzUKFQ0JY7GtDXWiifu21GQr5BPHnRdQ1dCQg78OzXKHYxd6
/SzC7DBb86R0QdfpladhSu0a8hg9m0jlle1/DxBZUBZhhQun+YFnKPecN5/hoOm1
my2S1tSn4TRIK9EFAspmd/J+VtK8Mk8baD2wTylK7WP4YqIRtaiR0is8Zy3X/cKp
HABgk+sit28f7Gkv4G4+zIj04e8P5YsZJmPieG1Axke8Yx9TrTberhFP0QM453KQ
qC8qzAO8RT/CwtusqcKNK+1Tn5oNqrra7YhU+HZZujL1Uc20RvHa8gsOy+MR3Pek
1Oyk3CUHgXgrl0GrRn6xu/SJzIBW1zetW+J1LGulGZWqDZTiPkRraalCuGqHwqmp
dL+tZD+dKjcDGmWzTSffDBF5OtCuiLfmked3L6IaTSzYKJtbhXLQmRt+DpBGO1oJ
IFrFIV2l5XnRVfR3zdF0ZHrX/wv3jRaz8pD5LD0K8eNgZMOrvcvZc185oIEHn6vb
HKEh9dCwYaP4De3jdUp9QEcovX562ZdDIugnwqBIjzS/BWPnvjf0VA1A0q4wWaqi
dS1ITR/jQWInTnsrTYI8z/VgvfmeAmYq849F975g54R5BR6R++7ol0oA4T6fVubu
QQxBwX/heAnnqfB82cPvKsbVaZ/cesuPep/t8Vm6nL+W/S37GdljDbgxE+VgOeeF
ciRoRQWloqcyrEBC6UKA7J7S9uCejJV31buSA7WB8VCNsa4oKQ145EYSQmc4Sha9
R/DinnejDaCx1wDuM4G/n9dJT5QHVW/irt19vP4zgu0dMjyzTWypsgi8VpUXP3gn
uAkt2dZZtBgwgcxGcXhmhgqWxNYLkhq2IkT2b8SauBEinBaWXbfSTeGLv2S4SiRP
tXYzPTyCH+AlxdJMTztqJsI0LNVwKlCsMBjn0bleJopvs7ZbvjpmregrdIMYnxAx
f7ERMmSWzKSgQuEzn3az5zPL3ybwNBQoJExetajHu9Jex/SviXpdGI0vFM/dILCT
uEF9t4A6WEd8lFT8ZCYNPO2k70t5C2pOvpW0pf0uleXfPYofMtznrKnx6sJ8cJaw
VkRCJdCjRPkUurJJq9iK3uo3B1INP4mdo2dK9ySpB3co+5wNOL6Gut0G7vVdka+6
cj/CLukN6jgJZSfhYJMuecPVZ6QG9Pkkw2iyMhGrfRbzJko+Uhv/t/dMbXoCTpE4
csfc0Pe35e3gDy457TifVZ2qdtTUtstB4mO7kwtazQj5DZrntzq60Ua4GdlA3+XB
VQ1ui5OgIXEQRG4lRpo7nLQMMCQKRhRWwSDHiVKhTv3cC7ukdYA0BHLBL3iNGtGE
7ZjvDwyas8vY+PYKvyTC26M7/zOPg5nKq5/eK+kVJRJRfZ5M6FbLcLKZEIfNb9Pt
Bbx7imCfsQrSuK6zhGfx8//sEW4hFGQgAJ4/Oi6CqKtwa6+17ab5xAvV5h/euVtf
3sXa5jDL5+KcHHc6y+No5wlQn/InNmlhC4Id+RYbgH7AcKC1rAzr19GCC0qT0cIG
FZaqGSyyNM9+KO0KQgiq8TizM/tMMQR8IQvYCD8fxtU7ccjJ1PniWE4Hw6XC1kay
9GnAOe7iAdhkNxHY3Axt6cMlSNy5lMacR+MQKG2caBlU8oVCGf4FIMHVeG6IEr4i
qpFBvxPM1gWQmf248DEnNPzNH2OPpq0XuI0EdzZU3jxdWfiJeLng8o9VB36rggm3
UxuKf2+OmkuSHY7d3ZSCz4s2sWRfROVn1nVo1blXkQe0DSl81zCFfhh2yi2U5Rp/
HpcwXa1+l7c2KttcS9YKTsy8vEpE7YE644+Wr8R/K5jQQhfzLKQG7G9IBkErzyv3
qAN5PvKzyZnBRQbmWEcR88NYYTrcQFtcYToPpxMaSVJU2q2Ro9Wb4UGYVWRJnGdg
q/RTP4Mk8du0tn2wS9VGQtts8b2js3653byT/oi4eMybGIZoZAX+MPEfZe4EHT/P
SnWTjJyCkwifa2DqKK/1hlZDpCruj1Wc+z1wmOOD0A0r3DHxvqTCGif61UPsU5YC
/kxiHezCQvY2HVVczlEjN9eia2LPOgAcSYAkRwDjhbcII529Cc07pJqv0UE/Xo9n
UMKIuq2M7sbPIRmaAmNL683d6LTYmqvwGMWI4Y19HUb9TIwymY3I1aafDMY7awdi
zigDKMrisBy1ZKMCHOgXPS0SHgnAgA2Hdf2KG6UjJaDuRQsISkDRSW0cWcyQzNj8
sfd+O/LMe0RpQuamdxrlYhMyoknQabTl6E0m/bIB69dYImoHjQpCgtmM0y/1xqir
4P8awU5l0xNkNq/LCUwcEjhgSxxTKLDTAGMIq2kDwcRc2Xac9kMRv92GyAcFh3Bo
7Cu3LbGMDSyLehaAjMeZHUCdk+7eq/D6pNZl+FLwyT7Rin5wAKeglmkHkaXVGIb+
dI0PMPqtrcFtiNIbXgJMvUSzE5s9Yj27Qw+2dIaRMqrQua3WjvzYIyt2hKmjCd41
0A/mzrUcEQF4SZwN4ajbrBWto/HJPp4hlXAatak7DdEmYuIc4Pae8O4U7P7MZc2i
J1VY+raNVp7ZH/zztb17WPgcp5CTsvD8xlJZjpr27JBskpsIfICjbV/E734Nc71n
`protect END_PROTECTED
