`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C7Rrnb6GN7VFQH59wWUxqLg3BpBqYqLdhmrpngzCWH6VDu0QM3gPnC+9F9ErF/az
VgLxngxkxf7JbgUNX1K4dYlKzgKrhfnwX2xMBqZt9JIUoekCZMCZ5/U/WwE6mGpA
a5p2YQrHqNNe5c8aVaW2AfVHSIJ8fvL8Xl45poAbQPP8wq5XFc6sWhTCj6KJOvV2
7e0bzWD2f6cnvElgerEmY7JpBATHp0QQ+jVmDvvkCpLekuwOHSlzCNAgFI8yW63u
bK1+elsAffu+haUkBda52dsK11HqYucP42ob4Vmi4gfDQcwIY7Vi86AiB8tsVT4z
q0bFmv0FJR74kFXaaekIYn015tLuNhi3LMP6H6N599xM9RiZQFVUKxusozU9TCMx
oJwbpkA0xStY2iaPU2vTcEdC3k9TEWIHNhSeZD8GCESfD3EjLc22VlNOXXzdzp8S
kgYDGST+N0SbqsI/IAe/v4CuHyXsUAGprnirArOJi3zExXo75pAf8F3uZ+87gfv1
DDUIYmR0vADk75suQnnLxQom6e9yTllp5ijRK0fapTGOGgK7BFAPNtra51uxZ63D
JOSUwziY7hkP5FAStycj2W7sWgc1j8ZBbp/1lD6MV74mrDT512EtBazNpZCmgXNV
pEU3FAc5tlMF1ytoRdb50hLX0Xa1ny+makdPyIPc+kaEMqbj0qDq4Bxj2GR0926J
AYUG7SLxUxQ0eyKh74iyLTvirZ+e+Pn1y/m48MDQa9vdyxh2L0CiI74KX0O6cY9T
VKxW6OQA6nsl4G4ZnOHqmIVzn0qqYDdD3QxEVxLYKjjH0Az4YnVtCUT3t2CSf+MV
aCTnCrn1OaaQZWu2jiou1mU17zEgPnOsV2XzGUVM2HntPM/vHWu4JOZJAGABYkHB
YkwjwG+lyoptZuLXH+uRy5wJRRNH2HRRjDL+2ggr2M9DkrQycP65La3S2rOASGhM
WiSUmTPiNEY15LNp7feaONVKT0pxLlLadb9PN942V21f1uk08McNYYVcryTFe78q
sebtBqI5Lag2VVLt1mc0Ndce5aVgj+hmtUE82rsPctSVqdiNs2lD7iIdlr7dVOWq
HZVYKBWne7eLamSpTsCe0VEdo4ov/IipNgfsskpFQpYjMKUFQPYYV8DQheuRnQnx
mqvcvz/KLLBUG0dLD4icuS8tNTIKFiCdjPKU/YUHwuvOojl4VDK8oq9GHs9ruqgX
092RtI2Xp6vD3d6pCFQfvF+C2YYCAOESN15w/b2GLptWQQJyflDdZtP+b1VxXbg+
3Y4KtnhSshhXO3LcSsC89LmXbriIXXFA008o3NPpM6plk6KE0skGqzyMpWeVFmgg
N0XN8TDluQbPXuo0Ut5AU0HgcWMPPpR6m9NS7ejXe8R/6TPnRwoey5NxSRTPMg4f
xhHCgEi7CuZQYVvG2knpkJcXoieEEJ/51KsmENMOuO8+zvqgbAaRM/HBQlHWYTu+
mMp3/QCzflt+JNCzvkKMC4tdK7O0X/ai75AWGymQJr5EiXe4nR0TDThDc1n1zEId
c0tU1+RBwk49UnMYoxCWYVRxBv7GBkkANIm8LfCQl+OqUOBQcK3qURPKzofOsEpN
1Wv9/qgLGDBtS4Mzp1ek0vgs59HUNLVPKg3J1pwvP3zBXWz3X5UZ/vWm7gZDSqcQ
N7Z3ECiuJmpQ2sPzigKfC6DAIhVPNdmMid/IdgR5Y+wqgdqmnRogxw3VhFbW9ACI
o1Vp6RHiSVq3DfL3kh8BaQ29P4KGhRqfU0NSCRm9kkXq7HnjysYdZmkeRY0LwMsK
PbQngYH4hWeM79z4GQw1zhErriosJ4gC2SLyBuyiyx2mCmjHtEqPDTc8sIOChMHX
CcrQPTLlZwJK4Km2qaiCmkJe2Io9YmzROq82nkT/5a5psm0o/HvbKntSvZAXT2HD
IfglLXZiaxFe2qzq5mENTDMAEnVqsDIR7SPi4QaSJwcEc7coiXnlrtSsttX74x7K
UpRWgAlivSzm9UbWM3Zxy/wHVEOSaY2+PHIAQkR/vKE4ox9LIZb2UnzQsPv+u8eb
/ESKnEqGxFZ2htiBZJQkMAUKG+6R20YHQv0eEFcYcg07GcuHWtqxtNrS4JswbS5w
pTi3uZtGtUclgKQWRlsY4uc/5rwQ5Pk10cKVzQfqdNA5jETu6AF508bIWGuKaoso
RhBr7VW9lViY/7op3iFCq3jgmInLnUqLxli6E2nGVIm0gDX86TKIbW61DvHINzXX
zCoVSeCbkoOsqxcB9GGZPziiWGWMBjt89m5Z8TRDyf06V7jm12Oh9hYwlsu8DPXZ
5eDwLqWCI4sQB33z9umHLZA8Bs4Dn1PqTgNY9tfYzG5Aa1BVc99z3OMMwGSIXtWU
hAXphNeA9NSWIPS9dhf2D7ESY/cPfbmOih7kMh2h4A+5m1KXPlIMDtp/LUVAbVIU
5stMOI7MdfNumYG8BC9uGdniljMg4Lk4oycjHllp2AwtBE30KiAis7xPjBsh0x9v
3TqZOEUN4qchX/RH9fEnwT7tIG/NrGOUP3DalDwB1i106aLrCxDAeXwoRs+FBbGU
5uxa+3izoLAmOl8S4ei4SFhzYtXQfzyjrcfH3JQ3VQC3SU+eBD6uH6beSn1a6J4k
uJFCwlRgWQ5Z3LiFw/6FVWzEAy5Mo9/cDb4EuG3wzlgxmE3roWFhRt6YBhaOje8y
aAGXHcfOATMlgLrXOzxC0/m3+G/0oG2U3HachJhXmQlDgV56bdf9l6TGzMptM1wr
Hjx9HIC3ir3TXlYFntdDFc4orNMb7D21MRhX/7ezWvRAf62pOt+FeC1dBFIkwLMc
wAcVh8amZLZVTNgNIH4MO8b9kPnbQa9LAiCPRnrFp0f0GEyjqccmwscCVbLFp3xg
Q1q85f1P5+1ikZzhM1GyxSL9xryR63YTkmnYwxaOKBm5ccwYCt0PUOAh728WeedI
/Nr99qmPCdVozG3wgmKtIWl4JRFn4Hu6to5O/jy4HNtwduk3NxISrwVTPaO/sOZE
XfORULNeDN1oXGHTiE7iyYV8khoK6nS/5jWxhuBR2UPg9TGnrffIVAzksJCLCeZb
K8j6R1MJ0AvfhBaCvfr2wbhFw7PSOkFypvMwxBssBEdx1Z6e2uYHl9x00ro+nLIF
9yesPlsarKx5gAPATPETq0vgvlnvBJWuHARHS2rYGoUAtONnuRCDgz1QUtANeqHs
KSvXMI7nTLSFPLtvcfreXPNSxJGw0EMkphVkDciFs0YJMApp7VPxTbfYNE4SdLYB
suvqtdPD/7pqptfrUg44e7ka11l2kuotp9eCV+DXYIticsHyUgdL1H2JxJm0s+RO
tzte/suIVQ6S53urVQN6O11FFhzWS46Wm+CvtN147b5pzBUbVsVKKWtTGg+6GjCy
5EypLNcqwLDQBnhl4EyrMi1UoW+OnT/pAERS4L2dPK94LeMz2DsCFYoGKmcg54uP
w9+XOJU0XsPUQAeTEGwtKCkHJYJ2lDPTjwHSoiQ9UKDLNMKTisErYKHppZY6DXRC
e73Eobxm5L2UMPtE0124lt4z1mLqCknTQ2q8tqoZRejrXjlaGP6O51raGHHLBrqp
WB+3POUw6kkJ+kiGLlixr24fAd7Bbei35dch1K6/ryJxEO8KAiZyjLnSW4WsLRkG
qNsXhEkwSw+v59+x0XyW5evHpD7VvRT7mPJ9Vef1I5s0rIWgAZ28GQrlwsoX1HE8
iJxFc5rdo2RfrRjVt2Ea7t9nTtya3RLA4fpouZdaz5WNRlKgzVkfu8kVgJGI3YDt
dvpVqFX8+6RVS2VedCAkHUa0IJ1gTuubz3AKqS7Wga1XNlEBEB5o7WTGe6JYicJi
hHpG8UnEizl+BNYGoz+wKhp3tCJU06Dd2WaLOB/fol3xyLp8pfJileZtit7hVodS
GvEFrKWy+Xbr+Bluej2DB6AEiItFU1YrS7h34t1GFOkMf+euBIE/srpRplMDES/k
WKfVwYNdl7PanzHhX1RpKNCffKc5IQHavVrWXlVqVkOWNhsalCXDhZL9N3JYVeVo
aphd56glNeTR5Pf2jG2az6UisXBUVKC/eA4TDUlte4/iSREIAJofwBbFG4IquJ6z
15X/s/klgtZeZZeLubark3qHbwYC6bKIlXLzVXyOudFseeGo+rBytYnRnMRiptAU
o/wjtLKs1v9JnSFtqA0NBb5YDeYTEwgXDDCSkQ+tAKjdflKq+fctiboqY7kSWtqA
ZnWwMFMXBMyp3bWWNGMach/Ckl4LqYkd9t5XfbpFtf5IMLlrfWcL1S8aOqMqNBhy
Cmejwa3WAK7gJzQVhmoeoztlSftDdUwbOSyq4W4pRGwJ64sjj5kEUM870cpaP0eR
JTB4czGmG/wMufIM7t44Ufbvm+PjtVJNLoBit3sAV1pUOMzVMiNifEri6cKIW7Kf
kZNhCdZ24x+Mv66TTQD25C/0VfW1Ll/wUTYWKVuRK6y7IW0sFsPpIxfv4IvpkEs7
8CfKeM1rAV1HC1aSlHUOvzNX+MUz2wAPOiPtzCNxID1FU/j792Bc2+4jb6QmVz5M
3lRBSPMsgNf2uzt6iL2mWt4tSr4uZtWVBqv4vxLh93KK4oQB6c/4XF1X2CZyfS75
efCM6a4Fz/Ffqy+8HGYrkkaqngEoMXUOzT6dB+CTDMYe6hEEfaNhTPh310wBWMaB
Ac0Ul6H0u9gcsxG6mbseK+9LSZ45HXHRoSHc5bqpplIkDWF9wCy9otWa3wzrlBpr
7aQUaPc+PiMOhsmqBi2WgErfJ9c9OZHZu9kWPF8MK0YbM/UTroXrVWRtDv2R12/9
nqKwyuh590ATezl5IEUrimzu/th7EPpqq1J0ec34lryjXJhwCGJILMgGYL/QqIrz
gh1YPkfXiJDJxmATYW1HUEhhwxN6FDFHE1/7/LSxp4rcCOEqHgqDyty5KVTpHAHs
mpSBdYM2htDbsv+mOOzASgG5bPsGBAH0fEJ+b70nXsqMtM/7zI9o6JWGlL1ZiHvO
B9MdU54lmuK+Mf5m2EQcKFJNnLQpYzrUJYUBXswNWNrydDVREpnRq0SAJ1AdVjAR
FKy1RFA0An1C/Gc9SdGTZjfp2rQrfZspq6WU+cETY9JsI1mVg/YyE5dQ5Kbrv8po
AiuLEjhPZZRAcm9K0EDLhBPiNGTFMhy7DTMEmyYbQVZAxxJmtWDSJ64UlHdU5Q6h
UdaSQj0hANBTMxf3xGK2JHyz+MYSywZJ4wmVe9q0QfBjEMw4Vnp791Z6Ke0JsoCg
klVJRFhcijqN5sR70ADFs7qEu77s5qbyS/TFDCeuXCpWr237TaP+8i2H0+6oNFTO
4fFBjNq+u5+43K1pTyvKSg2snZHvhjK38w72BmsonQOugpmLMoTBH2CbXJzl5vVI
u4OsGlKfxezapIzhmsvQRUZ8j28n0AlwzKUGxHcQOL4GbQPQMeJpJrr5NRrMove2
U90md6WJGfkU2YVHARj7YJ9NZdugJR6h8yUCmKQ3K1QB5vHXj0ZHTeyKZ32uRf+G
akoZojx0iDB5V4O6OJEWFpxq34Vssp8UDTKzcRMt5sbL34sC93FZl0TQT3+8GA7y
uJxvP+kr0Xue7/oK8wpOFBzwz9AI6NMRYdyr3308F12erVHl9xwN9w6LcLTTOoiV
ZuNNsJY9SfU+qaZQgEeBRBUXhOKHtlIkYO1Fv4HaIrWpi89GxsHqwXMeeR/w511d
q0Xd0SvV12h3FNeaObsHzVsKQAFcLLaEElu/JT7uvQmQdGUZcI3r30H4cXKzhXZ/
imJR/ZpXQ1rl0KwrV9PVfTKRF+NyK5NzHwrCEF7Df4O3c715QBZ+dajih1EF5t3f
TYAQY1xSlUA8cUQ1eVWmtB/D1kOmi/dmhkHWp+n9Ez1LPDEQ3hSI5cwTAcJxzSDv
Okc/c7kDhm93Ycpklf3nPItRCMSOQ8JgE+dd/HqlILdJsqHYq0FYKBx4OHTqIScQ
MZ/2WiNx5jULlM3j/3pqR7WTZML1K7wdxlsmS2uRvynuw3kquh3IvENomja5I/u8
eDz3KNqw5EOHoNXk9hreDriAwVgJsGgeTHoKNzLxSQVsUvJF3VhRDIEYIWQU/mAH
dTdtRUiOINBVHnNOYYoSONgIwNjAsNfp5F8mYx15pHpEMl2Eg0LKb3KCt3F75K6U
bYeWJBKKwtL3OT/Pk6ercpI7PJUz2/RG9iW3v0iZTEna0ePZ2+efrX5lMgfehV2k
7XHkWL1ggLgOEhD5w5Ymi3HGkBQTZG+Bol8OCN0NnbXStSz0gfM+rlwR4r+RAYzp
oo5MyWVKFZtXQUs8/HSGfUhasCEI0g8BFEH5pGyY6FLNeslRyqR+tZ0wNhrwoUnM
rRWwSfhMKX1mL7+NYBQ9VJLEBMYMAQbXiCSbzFdXVoehVmlDT4rjO8V6/b58W6rV
3LswDJ8r27VWM7v/6NUdaWqE0x4FSh+Tje++ppB6j3mzJJ8Xnb5E3qiyLUiTc2No
89zIOtqqa2VlR/Qclmi0fqQRo6FfWAB/QL5EvKHyfgl61NFppjean3XeV+kSZ4Ba
J3Q9skIMyofEqp4DsnpKcP2Widkv3lS/OBfK7FPWuznDCecQTFIQiuhcH2ByuzyW
jtQFcwQ16mWsFUtaOkIAEbU7SQqP4/B9abiwaRC2/OOlwqyQtlAcKq+E+aOxES+m
tw3v8YqC++maYhb06k4PDIa7WR1yVaKR1Zfer7wM7BieCADoq8T0DHkhDY4TSD5y
PYk4iWDJp2zykE9cCmgcgdCAz7DzkqhJEgFOW7XUVC5h9QW2CD6RMeTUT8Ig6OTA
9DNoNox92qAm2VQN8Y826Vsbvn0k5tVc1NDlDJjj8T1q1E8QymLCg1QLFoaRQr5G
V3o8mwZH0zVp9hTASFd2wZ97UY/WXaJq6nwXfmogQZzRrhh8vXJOSx4O9TM8/JuD
JD0auDsmdfNLrFN5OS0au/EHkaa5lpQqxJiZza4rHOloMxNx8X7WojIYS1BEkSY6
kesHjxLYqRhe9gDtEWOPu717QvrnQekRA0VXSvmmo5ttWf3NlvaPPE1Oq4OHpJoa
50J1MtBTb1pm1xKfm7nU0nUMkkJvs1yTn8+i+T02ojgZa5f8vhCXYma4X0qGLRsG
W4X/yiEyKiijPEP2LqyxJvsowmS5oymDal9ZSqcbBllP5V4o+M/fyiolF23OM/x3
hfEL9sc+o79Iu1Ox12GvFTLTWjXI4koPF2QMUJOlGJl7lIAmGqDp3+ZC8cyrKauA
pE7n6SirpntKimH8bpCycSoTyAyK7ClziiPBkuPwHSBIv1iYSwpzNS2NJmCSBlI/
HtTQiD9d/oMnlTj78UZN48TYAD4gIKsriQ7qmHnaRnleCraxPfd3VYdde7cnCaYE
gNs04QsHshErhwxk8XEPNNO8x6XX8CUD34T2KOq88YDNSL4NsBqHIFILyk+i5g+b
pXfhd0/hYoPe24lj6FQOeYWpHJ1+VSe/48Qxo2l/u9GYGbGxYHPToRck2IQTYtRh
txXce3mqv0eUdw4f2Q9IeF9o13b1v+5J4P1ShhRuDytpqyqVD88HFto7IWl73w56
g23ySzuYQLoJDozCs9XA9vWdELKaucAnUa38n2VFzqxEmHw6Du3YK2FzxV6ih1x8
jVO0I4obnYVqo1rlVMuK/H7EzRIFPDUUY+OUaqM6vdeh9xj2JDpUtY9Jazp2xRhr
iA8ZfVTGO1PBQYc54NnlqJW7uqKOUgXQTnyCZ5vQvX9KFG3EC6DznH/B6wpIzQFn
jgkhB0DI8Fa3bFt2amVfASXULjBeq10omKRxtq6DGxM92ZLXeTkKg493Uf2FwLwE
JAxkvEH+dyr3dcCU3nZH0nLsILEgVfrbNMSNDpc2DlO6XnDUmEN8oR0BOOFLbpOE
Pm07Z0MANpC/Gvpn6WfXyd1GvBEU0CAEu5Y1jaCzhBSzzi5BWMv9rIX389HRk0xI
Wa9hH8xEvcP5+y0P/kSi6D4ZHId+A0zn3e80/nP4//85U+Hy8dX62lLrb2kAMFgt
8nsyJO6wExOXI7TlWH3p0qc0xkCOgfFDy5u87GBVg5kHyv41JslI1wIKuvifCnGx
aX0On7cjYhbBNJN44NW8Hur6V3Pg2tHL+55457duqzFOBb1uph8WgNQMzarvtTe+
/xwltcyt1tQudl6ik+pxExJ2FvWGprQUT7lAwgNDO4OToiqjwuTdHZB2cPmPoMnu
JRticBriaSzIgb1bvOXEMfOIiLJUmGtG8QJ+tBOB6+t5wYRcYOtxOW9yJdSl0aJa
TfQD2YHP4kiLGbOdYwCwBhYqnerYY1K8kIlRQi56Lb9C6A2QghTICf7BCbN2L/NU
qqehrqFen3jItoMy0ctXuXDlCKs329xNUPEA+wblR7q0dgkdQnZ0YB1ysWv2FWm/
VLODzar3OgVV4N/q/cobo/V+bXIN7sdxYiyqOk6jjrclltCGmTNEL3W5PB1jLwDx
IS3PYqq9zzkZzxIRy7rFTo1FFCR1PsNQGesVIkvHesf651nKMRR/dG8Fj9C5No3E
c80FDgc/ErdFvScUKfwnEipAM2ScxmaSJZErjgspkxJgJwrmxra5GANg2d7iz5jz
4V8QG9yTYKZlbnYE5H58G7pKb9kPdY9zEb1pWf4+OxC+poRx/dP12YdgEzTC7AP5
f9v1WEG5SpgEwBGybE+IauLq3Rndd4fWvuOPILypfVvGY2cKqxBN62m8BGU534Az
mV4enlni/9XCQk2DUliedGp3uLaXy1mEDh+07LbMuaLLR/sRI4UixNrReZxatacO
8PhhjZQZSD3UeRGE0NVgXh5hB7qkb11tzlzxoNgH9Rw4kaPOSB65hurbmbooJuNB
B/KmEfP3lRZHIzhakPDQoBMLKFQEeC2NlOB32qRhMo+cgCgGrkNJmtxX+wEn63U9
JQscq8GZuQauJe539RHvP6Wd5jOVPXU5RqYkHo2JFANAK3IIY+JzScd3CUbqaB+f
UiLvNNhcc9lnb8ZYrf9GOvRozlrAxGZ39MWJyPZOjf+BimZ59D0IwQv2PtEsDDlI
h+F4/E4SbDtFKaxZ3+j6NcEzOHfaAfN7CYexiVeCmsRu6o3SZp4lk8VpDJxg1FYp
Jma69DCNNEDiASDl0iOdKYzkNhFdCVdMJrKkg6m1MP3mv9k2r2YpQKEUrq3gmHCj
zmndg/lsC+QurOuLpX2p1WDpFKZfSJPQHtb0hKM75YJ2CL7+jTUNt6g966iB7V82
IcvEgo6SXWgPEj+JXCHwKJpX1w1wd0Job+61FHiQnr75FqfNAx1Wy58Dcnw+FPXH
R3idy8+UtSpZikK+pnBRWc9kwEpoiF4oiQamtIXKp6t/X9w9zwMzScvvShoZFAZ9
WA7GqpK1fvrgxDyGb7CpsFzzNixuDUnNqf4NELhb0J/Y/QA34Fwst/VBMXwg9Aim
6AAzI1mkvuVI4aGI/3pwtbIbu5iBn81itRWMk5gRdYupkJNHgaV6pwyiRSDMGAws
67xgKmwMabH15Hso1ePKvHCUpZ8uw51bD9uuA/ir0xLddBOYpP/Tr7z4U1cYOA6N
24htQRBVfZFnvGpmvPUnC8bmoCqpxcsNoMsf0wvnUppVL4rnp07Al/TM1arHl0zT
dYfyzZ3PZybRd/o9eLIXhG5J81Hazz7I6pKDqWy37Ov88QTlkXuRqhGAYAqFzLhB
lhz81nhV0xpcaeXzT86G/tc0Es5wLI5bcPSNj1ndMxoV9UvP+7ZWBKADXWmQoMhc
lF6so/6O35REpN/ggeiwxP8OyJw33npGg0Pln9x1kPfOCHVC7tPcWuDg009TKWiZ
Kp9dCpwmCgr3UP0SgCi/NMwuAcF6WojUZgBxy5oizNOWoWViAiRuTZUETkTQPwAL
OM38fR/mo79N6s9ggsAtfKDSyFlSCBWGgui+vXtVqEMUMhb5mayrS41ls3QbHWi0
g9pCwZ8iF2phOl68+zeYufaWkSwvB6wfbp/1ZOH+mKkESBYnC0RNnHW0IwnHQquA
EbQfP2ZZbhRh3knyHwLXgY06tuvS3xw9scg3GeH4YnP2uEObO0tk6yL8G8TrtO/F
3WuYxl4uJJ0TLQIH1W5XEF/0E16On8ZmKUzwwFsBw0Ri3Otf8HcHGEXpQzS0+dAr
2PgrVOUbDzF7TGrkchUDCOFopLp6LB9WI4g/ePnPO0+10dKMz4BvagdXhaHAG5gx
f0//oXu3P5tA3VBS/uGf6wsapOLrFkfkAxA3PaCTLfIfwyzcliJfUIu+jyYwFbEU
jK6iq571kBAfVkyh12NGSsH22H3GMyFJJzvrx6l4juRv9bV+fI4bGj5Rrl3xPxln
znJBwpzHHTl15tkE1FewZCvDoW4tKLi2HvqPeR63kFTbwuQL61U0+YcQOudSTvpt
zZHzJvRAld1hVK10div47ckC4dEUtuEcmBrLxTwzudCwozogbzBJ45UC6vMNWe5F
nJPSqc6bHBTXHX6XNgwPc3KitezB9kRWjqS9JeyWtFODeFVKyDUR/ocfyCvJgB7A
EynCGzGjSdTlS6BNtIYVbh1f6h+qISxx7sRs/wpC84YKCC36cbuRH8HtcsNq8BJb
jt+2cVcVkkHPkObV/eluBT+k5K8hlJLeId1AKfUVUzAsWT2J/CFDOTWs3MXBKwV8
hVHHptqDJQiVWwp8WkqKdACsakqy+ibkEsyXJ/X3lHcE66gKICZH/yPfqQZHDFLY
A2sVadUzAwyJIvKtNufdroCiiofTJY26i1WYtjJdtp4MC6fvpuQlD74KMEt7gcJe
ICc7rjtznN7ASD9QBREd6CVYUuYIdO6KbAH/SakqyU+QVgu7izOEjUz3P8C2Fibu
uKLmqRW4vp6J2ozkE3AMSdBBN2DpsCW/++EY1M4vNFqNs4LmaF/b0fNrM4xfO1Dy
FYebiDPIjiaOH8YB2vprsLqYqsO+lx6GvPytzN8M56A86LMtvB7QOYMA+NtteYEv
bRbwWwaiOL8MP0hU1MzeXMsbQAyoZwX9tPcaKishbL4xCwFjh9JBbexWzwTHT0md
OBtpk9+q2JW031Kxd/cXZulj2bVmVuyUmqJ5K+803uSMRXm5P5RfM8cXh//TmfZn
0xB7JRS/phFBBq3c6O6Jr4atfSmcjWW8kKC1LUG9SHtEU83IwqcoxsnPci3GE3XZ
i+mByD19iS6CBrdnyCSpA6TVcDpLzzffIMe313RpGZZKpgudx5/A+bJg3umXUNIJ
GJA/howE9nUveIcEBMxTkRy0UFZsuUmfsFipqx2Xff+BPLZoCR/6BpEkbR5btoQB
N4dA7oghP5mShwlmrJfeSeObIqmMKxwps3BGlADonMfjJMsbL5gSyqNVy6Dj8Kuj
OJk4QCuErbw6MQuDruraxYQ8+6ycUpEJFx0uuEchEZ1RABpvbaamL8U0IW+Pp5kh
srO/XMMx+SdzIDhm69yxyayx8L67W/puPCQbCdFtdipYc/yTWL5VSLN5+a0i7xwk
1oodFk3vewLRiNHgwAF3V9iwuMi+WqiYHUfY5peiq389SG/ntVzXYVoNyjtLA1m2
ZQ8g3NVsBZ01W+DqenS/vpSVAy+aas9oIVQuvANVDLM/yH+Bi/gEq+cX7BSEwHGU
D3lYakfeym92Kv8cvbxoZMMIawycnk1MZ6f1vstui+peewQIC0xcUg8uTeuzCwso
xrEt6UZ9b4ib7eUrOTMtpdRI2CjuoKtyoK7gGbIj5cHfLQWM7vgRNooPYysGksj4
pl0mAfBi+4RNN8W8BsBEM8ps8t4/ighKgvQEjyTudg1Oq/E3OB6zOWMYsR5AHdVg
oYP9zZacEEe+gFz9vSEky2USI/DhbQSDa9qK9DIkyewLbiJ/cKFJvOiE+JFVfuZi
nrBMadrZs/bZYlkl/j9TOl/MtPkQwMDn2K0VNiD2vViwJ1o6e1fejFaWzUABVwpT
hPJ42iEBRxnC7kZP4tiaCgMYvW0JzO/b0KJwbMKqfHf4ZYRZB6WIcVONQSA+z97f
bPSa79fMq3uSVr/33xXvGBV5B1ju/IUezF3uYmTLG5aD5LZ3up/Rzk4VNbkCuIKL
z4Rz0rj80MCgzTln+ehMyPmh3oe9gjPAXgyE6Le20RbPyCsQA/cLhVDIjeVWgRTF
T6qgSdOBUsQazna0kY7LLXrZLUG9Lxjj+rKiAnQcLezLFE9ncHr9sTpDla1ojcwQ
86V3rJ1pInqLfr+hN2UbURSe5xa6VtWtcmdsv4jx5TZCImHQN+Pg0wnylFvthxfs
AGK8EUgdHMOIix74NMwnb9kPAUa8TaCp3YYXLKtFhhwNoWlwjwjjzXXbSWwH76GF
MwfD7va+h7GJrNY82x0N1tm7Z1OKkHfk0hi3j0eRSeqAja4qM8T2ing/XqsH4RJk
iAKntWLQjvE9Dq6NWUalQ+vV0JNcUe23xJaxyFzVqfqKsdEXEDAbJzhLCC72o7L1
+pHfxGfOyNZkW+WK/hOEDOxtpGbd7B1bnNyNy4gTiwCKstKpHNU+bNDI3KmKflt3
UBQzv9XI9osXLLgDjzFEvFahz3Y2Hhz7BOk+uMbpPCnfBArAmdpgkT7+eAXuaMQ3
IGMf9ynynZQBZpn1Ez32H8xsITdqusGj+D9pyOi2WZeoPmshJatLgkFrBs43sCua
AiqcrjrLKkIBsrH0GGvHvM+Q098TrYWmrYkZAN9PEFhleZlrcBiCE4rD2RqOEM0V
IKl+hF4rHlMKyaSLDSKLBtxISDW/mxcBoGH+tSBo62rWWJ5hDy3f4eEUHC0k9UNu
TsJJsJFb30V0O6sDGCeOyuVIWuJv1pDgbPIxIjkOEo6mURVjMdIXVF0cuhNfYswS
lmnDiDNhCLnyrW0K9aOixeABMPifJMZ678rGaUkXg2oBVC7+qhkvXG8+mxRbRByy
6UCQi8HcoK+ddHfnHwAvud9ZR2bdGzIlRYwz9SFMXT0++cOfcHPfIYaa5Ei8tBUj
lw1QN+Cq4+EI8asOxJDjZIPlAMkv4Vna9VVaz1J8cnAoNQCp7XjE22PUD3VgfGkD
jwZHJwPuXyR7i9kUy1cKtX9SiTDQmDTZ2J7dFO9HX0QcOVZHo0f7V/wuduRmzuXp
dxxkpCkShVDlpz+zWWU4TXQxIRfz3Qvw7DcbH25iF/WwdhAQerqmeV3V45ZPTEdm
pmp+A5iNY3xzL6lume3oboVTxGDH814FPL1b0MOFm6YN4Hxi6pmph5i/fZYsZioy
4+lbvEnx70JEQthNQfwqtk6MG+WV+5yMEU3+NSox0o6ue6sdTC2ZATxBZjkTYLhE
RggVbID+dmlfFic7PotOakSkgtQAr/ce4QxA6jx2v+XmLdj5TL6I0J1UGB8CGxy0
ZY4HeyMGX03/cTxNiiAKBCeSgzkQ2TTeODOfXMJtlOJOax5t24hlfNlsHNYBrp2V
PSyJDgORlezUuucxh8lGN9cgICL9fKUCOEkOMrPBOh1JbmnrGTLmF2bVTUoCyB6/
2Y/bsD2QmBjS1VpVYYMEhjmSKAo3kqA4w0vG0ZLdk9V1du6TJ7fMxdjehA4v9swE
Lv+sbg40dW6tZB1jVivr0MjYQbah2Oe/ydRdOz3A5Nfy+4oj6PcakvvdxqlggywX
iTQpPYaG03KbUAkHiKEC00R/2OqGxoaJIWGXKDmkR28mbEG4EmU6jUZWtvTApQXa
whvb89fEgYaDZcCg+FbWaOoNX8oWk5npB28hPv2fEIrZau7z7uHzK9w2pS0yN+dr
m47Kpdn+rpeSvu8QEYO/7RhKEXUbf0nr+OiUot0OLNhqAGE0beNuCls5O813u4VF
iKjjunylvfEncINgX0W5SFVKppO36JPNbALgbChiBea3pqLBuKYcIrqC0zdec15p
66ZG9/lUAwydCLZe3uHeobPRMWwEKVTgy29xYEcv0zam31K+UMRsZ8dexqtatNL6
UV4+xRnSQD9fKAMzw/I+APp33sFRX+6CX1YfozV/4fErlN95SGNsXo6CT819Jt0o
s0tZmQoNNB6KaYTN8xKQ/3sN1e0+WZ4mDGt5l4qP0gQKYmGNAIISTOqCAwzcsLva
fvT+s7mvKehs5xCEL055QIDhPFnm5nh4q22GyGaAsYlzfUiN+yC+tEE3ea9TcNob
j1Az6QB9EKbISkUnMxK+rnvXOUX2HOhV+/DSLpxln1ZuJPlLKy9+Q1QXvooBgr/5
Ay2+alwAqlKOlJumCcrE1tfQ/J1LySEeCR7HA8++vuu3pqHSh9ErbhsIJmOS+tSe
DQlAAfynhzGKM6aPMPb3p96ZHRLpn69KylikD8jalNSC3JjZuPlwvyM2Pn2Vqifl
8MCarbTkcuH4J/F+miukyBF30cypw+c45r0gH1GZ1fDxd1luI5y5I0KAvtA02Afs
L+4SeaQnd+wdhJRc54bFL7BVzFoFU591gGpi9fg9iLIx7iPbeDwrFPF1PVC8tM9C
WlY+ZKhlpi3HJE/rBnNEgJ2piHKo2KFNjz5sXqXc6v2IKNGP5WX7DUDqOvq/XlTS
lsrFMQoKrZlqwVIOh0dqMT8fyyR2rx/XNjvBcOEvFziCLiUbqOyZ0UZ+5U9+BU7Z
lK07iEdTavZ0lDC8R4+CHHgJXuP8OJbewhjWi6WGt2F4gCi3iZuZdKYIF1WB3ttw
p4P0/4DB2wH0vN9YW86pzb/AysUbxOSE5xwlzjzmpSWLDg9HvovSWUBiPXtpvesA
oLo+/vhJaBjVWggpxlsyI22jFUlIyzFfBiuo5mOr9u2tcpsiKz6/ka8+4reRzI5Z
ML0ly3v/zbgyFCQPsZ7gHUTb+zWoSSMNSteEhvVlD+vRUCGYzrvBbHIgJYEWK+ub
YZXB3evPa8kF6RLoPd6xLDL3VkHzNlWeSqIEJ8rU9h6BE4N9hr5+QYTPtsQ+3992
K0yKzbomxUBZNWQHUtAaqqybF9/Zh1jdb6osWqCGf8pzts4/EfK5cRa85T9FHn6Q
1c7duJn5F1WcrsaPYqy7OqesfuPd9wKC+PQ45h33tRzK/MI1UvsUp+BPu6+jRDSM
a52oa0IpLkXUWR9PJwKPAxO5OiHaYEsT3BqBNTYwF/QNvbeWr0cSb/sjGFR00rqc
m/9XkWcPaJZ2+bAoSHocmpKSRpsaffSW/l1YL1fqqP9gMo4Ukt4ysOhEnDZdaegj
4UyPZeDGNC5JIM2FhEWA+iWyRHowHS4xe7Uu5TZSOa7HYgvQF4E1ghnnk6uZAYTR
qZPnZYCZwC+gqHcpo7O+wVZYflKtgnP6eWN6t0Wync6G6kj7iI8zxaUVD+Cgh83Z
VrY1bB7u5y0FkzuUeVl//eaSJX83FkpHVsn/igHSVBtZ33xAoCf5nyqUzu/4yCdl
SFe1xvRpuJlRD3SnH5YJStmwSxMxouuOsZ8mRpwB+9q2f2z1uyccv8cqNw9Ih7KB
qTFZW/l0YdCtzQ9ryV+62ITOkOI5sMVjttQM5GWYVOxVJbvzS4jSBc2IB43/Ws6V
1d1O7QVGDXbOzkC67p0bocV3QHMT2Mzc8Wy2CsqBFAFypcUQ9x16pRzlZ2StF+s2
XuA5DYHBkSeBg7bowo7jvc7RzDrkuaTORsNOMPVPWMoAaFhAhh8m7rm1LbAW/CqK
lSI7EaGuZnm5HXF6O4mQLYCPQTS7YVMxqQVPGPFVW2PFOhULO7hJPIWGWz7nlj+7
K4Z8PLXFcPqrIpL3/jzYfAPSFY0ajgUvetfHmQn58aLgbEIesf11vDPOB6zVUQQs
At1cQt6Ipg3sV/yCdDWKV1eCYvdWDsAIrxH030ef3/zlgFCRwuTXNPFz2Sl4GBTi
iAv6faQ4J/vf3IZng40+K7mBy18FVQAawZvlrpOWnKfwGE/RapxTmjYlolxucL1C
mjOl1L/SuGY+FuLOl6mYJH2Le8C55PzUNTNmX6n3JdlHYlTLMs61Il7jvNmw4bwm
NtSjzHi/PT0c0nIhFtnJU0WH215uCFhwnwZ9R5GAquGIwMb0n7sAiieYjVy5+TGl
s4ett+E8knI0rblrFkauCd3VxfltRMvwjWKUuvH3viIwB/L+HfSaOz2ujjkXJDFE
TxxM2BCg0n1eTrt7p4ibpsiz00jniG3+GjkcOKjO838IjzHrPJSNKus3ixl+KCmG
tCcRPmnfrhY71m5mCqy1/VgkBPvdcsAtH/JNYUg1z9ncI8vMq9H2aYOWeGFo+Zej
mXpdxhjtktsyBor6BKO9BAgiyFS3cbWaaMBbShNWR3Q480yun6DxGBLSFhcwY8MM
OSre1CHRDHX/3v4mEL6fFTm1H5xLJ+JtXe3uhqb617VS+lmPW28i6sm2XMzfSWuA
i0trIXm9A7gv6mc/eurVKudn23yvYk+AE/i++J1CfGCUX4Zr1DgAe/daRG/V1+zl
bUai36BXo7Z0ZNvjOEjJt/eBnyhszh2fOOr25J0CDMyLjbcPa99z/sJqIQC9wP1x
5CFwgTj1PkpUtiB75+UY+aI6Bim6VwtV0Sis0clPCR6igHlfsphVKqHulYBnajD3
PlbkEgpEdUWogNsydJbzRIrnkXHLC3lVrU7Ojqf21SHQK0PONGkB9NUtaHJ2xPSF
jQginAsiNVY/PAfFhHXc/9+bOUXSGOk38CNvks+dYUelBjrmA43FOAh0TVO0GpC8
4vtXeqW/4RkGqcWhJIbDb9qSFDdYrC2eIwdRvLbaKmD7/n2ZuKlQHcsTuUGFo2r9
NrjL4v3PvsWCGDEiQOvcqv9UMItat9LkoSwJsCstu1Dnh14jpV3/BCh4B8uDM62R
JU/XZR0Noyz+lfKmGiXNNqe0OVTW7iHjKANczbrLnxvVGcFU16PgvHhFr9F1pTEB
dQ82NUDLkKNGJ0FSkNpkFETdkTXd4yJrhUwfg0wDVmmBQwCsmNcJq9XFlxK8mc67
ZuTsLGLpDGOKAvN4rckbWN4JcJS+KJ2MnE9db68IwQzzxHikDoKbEQ/TgS+iwcHt
VI1r8AQSXC3OjEDQnRk++KF+dGA40hzICNtp3hGgMXXdLelrUqXFukrOz8GpUIAY
Pts7+12KIFkmAygHSly21InNx9+NCh4amOHQkz9PitruoaZ+TZBGoly1e47kRulm
u8CWJNbsQK1XguqGtx9snXYOkAeb2LpXI9UckDVGq438ioock3zFTWTXNpZ0Td8q
TNyOJWb8mY5vhVKwd4QOlI04tiiUXKv5BPWLtlptGxdnkA6Ti2vTQF1fEo1tA0Hu
6pI1LSXsASiNldc30xe0jHybOaEZGERI1B/JWbajnqgRYTG2HtkUjyB51egys7Mv
u1tkHsQ0dCARVCiyjG7BmPzUkG/c4TyzRdgrT2mHjfb1Tfknd367Wqoq8+Qd5hGm
oiokY4Z2u9IJynNBn6lV/xKmpMGRPmPp+N3Rw18PT6iqIW9mbB1gOHMFhX7k4Dd6
3MMeZ9Dm56AnYolx4cJPab5dHeKjzjYScLpOFWVHgut5+bZNnHORiEYgX95yomdT
UEcwRuGY5p/rSIoBvMqsQC6Hg2jKceHRNPdol/b/IvSYHRxfW2mReXT6m0ufUrN/
8s+Re7r8kkVV5JU8o7IPqeNHECyEtJFRBK9pgwj6uFqxKuMxLzofgx7wRQ9oTxmP
IWKwZo695XYH2H3hTGzn4pQ2EnCmGbKme/LIyuPoLcyjhpPsQPxBYdiDqVdrSESL
q1ooRTQdMo3bfoqKVZE5UFP3XbsgfYC2bWdlIzBqk+LpJ4EGlwwKER2DKGgIrcOF
LG761hBSUltXatwpZtkht292A5FQ1fsP7hQ9G7DmCBoTLffUIg0x7sCfBe4WRNU5
kIyt/KTh4Pny1QaiPCFuVl3IjPKO/S52cB81z3TmzYbRJ1/e5haA4roSKHVE9sRr
w8MG6B7qiKOuyCnHH1LfAhKJOzyScaFgIrx6SJTpvKtgqCzEKSM3bmD2lNW2Lld9
tV5Jm2TlvuNfzhbQdOrx5iUNR5HgZ7lt+ELP3dY8gVML4pJXe4Xg5I3NsOcYpGoK
wBg/y7PzmWYFLOa9rmFJHcyxkrSP8xjaYUSHR8wzDPM5Lp9pNWjuImsNxlGY766V
ez00DoddUy26K/KsVXRayeRcLfw+BnavegRVpXk+IiX3cuWmVLB0MQsX4HNiNDHg
uCfRWTGcfLDIo9ndjWPBehIme0SP/DFpVCtqGuwjWf7Hx6cgWBZVZmtb4zhaMAcF
/VbhuqsZ7WxbBWwIUV4Sji6XOPQZjs/t7W+l5KNgx2kv9t5W5HboWB8F8p2EXdjJ
MJn/2JLMq/yHwp+3qDA9olg3pXAUFw5g2nGyD8Evl9l+k+9lf0ebaUnXiOvfDYEk
FxdBSa8SPLntz+vMiuQr+rDpb+jgWUFo47sHAaXa+fzFVPcMrPF7VuBTYN8zV+o1
SmA+k+t0BNmb0nVYBbwELLBMOMjr3fl5e8+7ONuSmL1I3AnIdPsiHPpq5GFw95mE
kKVMW8Ahpq6ZWxLQR7y2c/r456wAgL5mWpx3+TkFshu9+bUtY4iUE7XbjQEtbk9w
RqBmcrD9pVRyQFA/CrwZL/MhJuT3RpD5zySbu8hzrhdIYMMP7gYpdHp8BR4yoEhP
s02b8SRic0gpSH5iG16/p/tHi19Uo2+fA/j5EmOJFYPS5C/awtYRqJvk8PhY7Vm0
z1xXa3RrUtRkwX86FVFcZgk1FPr/v+EaV9s33sQqwVPJtfS6//tsGY7MZeMvW7a0
JBYBzBQ+B1vOK5vj2tA8ZQmrTY5HjjjlP9WNqkNaN2GXYiJH1UvCXjPgmpAZdAfd
99Nmbb7BippzQMsk4HanrMhFyBqMrk2FOZVTs9xBx0eGJYIs/YRZ0ob5QvbfeFBl
9MWChscIgGVYJZerpF2f+qo2kiiNSwYRvUPA+pCmwg+iBtRZeJfqTyh1tD+cVshE
h+Zi47l64BIQ/aSYlVILQmq4zNZYXwOeR7p07FomHsUc/gCLFU8aY5Gy5RblaiAP
LaUDiP3Y6g/wNVji7BQimPhzDnsG6yHZ8wTiuJrURsx+M89adJS3y6AYYVRzD7ZC
MkTEJ05NCXvS41i1kWheRfcco7GTYHJOB5oRJLpdBnXaWJcWrPTBcUX6yn1+4Oab
prCMMxQtSROYrqfUf7CsEzM3xdOqcPfZn0zlJAVYoBJXqg2wdEOAF4WZgOJK2lWh
VfHmGXNI5bjhNixR9BMktqxX07gHd1ItUFcmWqhnn5SBllpTWY0KH7Vxy2W8Z25s
N1ODu4RaCeZ5TJeq3fxpaqs6cn5JA4+Z3e47DMCDHCaarp5lw5DzvvdMhvZxBjAl
BZgve15PfMsWzdwQzaK9tBV7O34ntfZhc/reZJHuSk4UBeswzXnd8eLiFGcVrFKA
1OE1S5TnW1URv2cCV1d7S+DOSzhWl1Ptrr/CAiCnUA+nQpZ4fGl0tElJiE+C/stQ
f+FAtzLOsr1FfQiYy3Pbo8EhfLl40kjlv1Sb8GeXOZ+rlk/mFZB6oegCx4hlRIqC
v5Gpt4ujf76xq0ScoNdcB9HzrBG4d8RpXrrJtg9bipAV9NjIh1ViHXabNhAP31of
kL2LDjZEaxbz4YelTG03sFDOqF3q5X+Hi3MUwjLnO/uoRBciwTirK/Qw5tiJ4t66
Nrodj4zX/S59TE00rGm/I3FWmyPCbO9gGRengIz//5ViGuY8wJfmiyfTCwfxKgzG
G6IJ+h92vM0SbyfJR5L7yXFAYriLZiu4NZZaGkFEwY0vsaVfZh6WgHAibr0cVQj/
Wo01gcD8HXYQbxEX9iXumbwtaAAHUjsJjt8bjXQUh6OL9RvpRb5YaCdDFqrBiPEx
sTwZ9ajp+T2SDU2epyEdjN3KQcSTRddb3Yz8YEab0+xPVzvJG1NqbnLaDUNIoVwJ
P579AWFNwHydtf+IzH9B3IvLmAslxoQsuWo6zW91lCCi8MnN9ffJziE/XcFrGb++
K4udyyUvESY8Me3zPmzm0IV+nyyNXPSCH6bE0CaRLBvt5kMUed3/p+kWgg8BhoUt
1gQyc0WHPSYA7Nh1znxgtfOgTGQm948n269SdnuCIVMN/VFIrFaZdIRGqnvEVKLm
4SmHHp5mqGXyJCsYnljIvEA53Rq5AIjP+7pyh65cjjhhrKIllK5ypBP1LHQGOdnJ
Zvbgm05dum5qmf1VrN3PAtIlWTmcpuybmG8ml4MfZWS5kXpKdDTAPZMJIpqdT0re
Ix8+k4YBU9LXXCDu9r2RtgVRlJlGd5qMb/lm8DF0CHO5f125+mSWWJ8XAnVLY3X7
+U9VmCd3Q2WCxmS5sQfHZersDgiSgkMcYJ7d8O+lvvgwoAwm9nDC+gScRDPe+jdT
vU4lQJuKdab1zYabs2+9+ZZOvOOa8e6VF6uCfc3QXvx2uL466eGo9l2NM2CaeUlR
W1dlJR8Uzd3ZcN+q8p3zGbjnNttYSjR8LGLWYEE3UkhnXcXibeWtUQQIfb6FS7UJ
KiEbWeHZJbL/+QcOGNAYBYKmOz4AEtAkgM4Bj9wldMaMLWOalwmCM8jYrrGALR8p
b81wsoeBN51/uicavvjH3MZUS2UDKhyxu1gdL3cby8DwvNyYqXKLSfOB/B8U2vYB
eiEkGPjnAbki4/+eO26+zkJ9YQgipWGLUmUS+E7LeWiE/eFgYzrAnXJSfN+Z2T2z
AIQFBL6RwjURPQj8PIQO8HNOIoFtSAnyo4sUpoDyCnQqAuzrsSNlDY4kU1N0vlqR
kPLwzjiTnWz07YD3aK0VRe+hSHIj+IdqIebDyh6TBrZ/ChMxiy64MabskN/IFKqW
P2frFblZkBl+j3w1wyXiLfHUnFfLC4lQzGsaZtH2Q7aKO8LlGEd/KF2hZS0If2r0
bJibhNnCcq9+f4iRyK3sjNXD6YwCmFL4ueLTY2L5qSdM+4eU2KdIiSYLeGbJ/gbf
DkZOFFDMzlC5H12MtqeQ/Lse0ZIfSQ0Sx84UNMBcMiQF5/yise5Wl1qm+S/BRbHg
BqkbmQEYhZBc3KHf8X9vZU5v9vWM9DdR0i6XNo7W3BeydHuWAODrIuq8MN4AuPxF
IK/f/1BlNAmQYzpRf+qfVSK9oIqDVO3q4exYjaw7AuBc9iRHveVB2r2rT4A48EYn
fJBprsFx2fIBdamoWObzaIvWOAb2NPG3157oCq7fYqvGFzfkX4cY5wTptfnF+/56
1QoyDOCzaeP5cJIHdv8iselsNbwJrAMzKsixnlkTC7B6H14GnaiMk7Q4M7fnBjWp
86XBkzIU4t5u5FBF5Btso0Wk3kZ49QlqOTBBCfuJG1yTXFGgFafKN+WgZurUsvU5
pCE2ytAyrzqI0y+Y6NkZbRDWKJ2B5oVSKs47/TWpxBFfSIAwnmLNbt4QS5zPs/U5
Mxfg813mmMdJ+yl539pEZPIo5oyk2FGGc3vDt1pUsJPM+GgdLNfTEXTjXUKWrg5l
aZfBxg8IuRlVSHpLWnLAQevGatUS+FMy7ZJeNSmVNmdxMTrAH3Qj0jUJ5aCXX5WI
tlsm4KL2+kbzItwsDSmiQalMZUxxSvHgaSZ6M4f9EOyfXAKejUUlOMfrQrIlrNCv
0G8vz+CR0kdKQTwp4AmIpo646eODPX7XMoBYZll/YOipHb9KpF3dTQL+sCywNGl+
jQcyGmBKBcKtG1mmexaWeDumRQ1fyyHQ0a50i+zrOtT+tTKObOXdcgq0UQ9FCq+L
HsOL3YhtSgz6nNowE9MqHLo+0jSKoypWHTxT0Afv+yWO3dsF5DvMNaOd45+4Sc3W
a4NROE0YdertW4InC7+OeBR/bvyXK0sNW9f6/vP+DF4Dt6Atyu3MNWPmep8As9wP
b7l8HIq6ZV+M6/8/g6CtNYI28c9LESPtRonFiaCw3/t0owHuhayGU9XHR7sdwmL5
kywUiKEKyxbWmnMVlsfxCd582irLy6vVYMrA5lC+VshmUI59ewkStS+289VDFUAd
7EwHDUOBSaW+aHFCCC2q43Vsl+YGnn5mMeQPFGy5Y6amLPLiag0EqRDwWlTHjoQg
sddBt9HCaZmwCDz0uFBg4kxbKkXJ4c470tfIsnbXbuMiJ2+y3LwLqdypZ+Ay0lwq
zm/31p+giNddj48yWR9Su+qHMeaQi3SLGX+GAVje5o0vUgkarhSoz7hNw+xACX8s
EEp+ZacUdzOABy8eQYow1+ZKIdakrNFz+KUnv7fuPddQRIaMar4zYCTZikP7Tek1
UCBLKd7QiKTpvif6NnjEmODtINubU9CJHSuKVCQK96kbGo5Xi5luP4SMroayZ4R8
eitXsFR6JvTCje7vMjKY+JLm+ScRlvrP2yU8Lv4vxVCyp65xlxWlR6jhaI43X2s3
dkVv6e8hESjAhYkICJxvk/w9vwys4Fa0si9iuibULlFKx2KAEAa6gNRuIhdCu4Zv
uvE83u1v6G2zYr1SUSKsJfFyMkuVmYPs4hUCmZN85/A+SeD768n1RQ4wnG7GepNa
Y/fEnEziodFAKdwxrrd5Tzufu0gKiZwjmxPJbmQVkNPiA75340ugASV5y9TSk/xo
ZEwf1Y2u9CGSop8xIgb6kcdMRpYHe82Ul8fIIRjdeI47++wJ4+Y+xGxppC00JvYB
MJVyEJ9nb9VpzHg6x1hd1D1fOVhcmpsrzqAo40q42yXODmOG+0BKuIwahFDPmv5I
Pe1kjmNVYzNDA1lAjffOrBmB4nvgVMmqDt/jJ/aj14gqpp7ef6KXX22DIrzmAY8A
UkACOoDfllORkgDNIPdEYMC9DpeuOTt+BzVfEqtYqpAQeZwYhsQsjo2w3VqGTRqH
NTXr/quKDNOprXWhd+mnLjr0SPkwd6o335nX5oOCjbb6y9vRoea39V9DFAsN+xYp
q2QpgC251IMmxEpa06RNpBhJ6zHx5BYbEqqYyBH3GFUXP13pNaauuncW5kUVOycB
BCF2Flb3OG5mtOu6SIE7GRR4Ot3f9PdS725G5e9U2LmlwxnuooFomKliYfPDo83O
6MOzektL3CKwhHerRjPl90q+zNCTY6z0XmSsmjUbBwnNJqZqa9LFc2Vd1MarAqHD
pqNthmj6Wp/8bK8M6p514/XBuKea76RswnyyIOyncjUmvXD9Jtr+FzBj+iAFZjM4
UOhiSDu8Q/ZyLGARgaHddX5S4tQfS7YUWcGcQVpL5maahkiq2jyYf105M0MDZzme
XAntBAUXY+nml9cmo3/bAn7qwPGTOvIuR3HtOS455JCUZi4hJBXUiJ9AfQF4lWJc
zujpAWkbbZrTzfjiDYFqnUw4jV0+J10v34+Z16epOyqDTn5bU148ANsvo6ciD7xW
qE3Ri82yPvMAwh53nWS6GI2TmxgsvtRS3hq37pTXHJ7TL5ztWS9Zrjr20TJZFWJU
BpCdjALzA+DiRyBhUGgah1ts+C8Ls2+lgISDWMRZZ5NhHa2rvWlNyiHUqe0O59nm
HkTEqTMlr8T97OCAI4WL7lT89VxA5OV1FhamaqK0L2tXcOIxodZ2g2FvQQ56NfBY
wW2ULAY0yxheBpo9RFosmiM0rAIkMBHNghsm2/fcy1m1zrECP0STLdC5SluwD1ic
P5TJYcKJbUFL073Ow2o+Urd7fKcAdEifDZiv0nnZVA0Hg8FRnptipVcqX1BdQg0w
OhQNcwzgoNX4Kdkyf2tpJ1Nh2UBiUuvu9FovzZnZDCvLk06WAuomh3+N5I1LFELQ
c0rPSdmxVG0hSu5jEthG+0g9WtBCEo8bi3ScaAKHvsd86A3F+TBpGIqkiP7m11Ou
vp8PFBpWkfrtfPKZ5YQgT8qudwHPw12rQsZmTFKM8BitVm7iwogWbi/jIKtE9fbv
JGswIOQZvd9hPIwUGqSPLjltT4Vxeyy1WaHXj91eExNrJrcirXmNQUJC9SRFlRG0
kDQGDtwCsA6WuuzWVo8xOPdophy/da5lKsgC9DRJW2AWffQf5HIWoYv95rAaOjsl
OGgtolSr16I9krydmjHM53oNaWyfwjfm58X8k+fXCs5Yg5ocXL8fW6hi9UZX4uE8
6RReEhRyH2NtFsKe60U5eSLF6Q9PTXvo3rHVln3fRuQq2K2LP42PAkjPI37y564q
liFjZjnhCtGCsk+8az5fmLhG2YU9N9t1Q1djP+9+2XrkQkbV44JyJ2pNLExYuiW4
j052yMq8DEYST2MikQRiybZT0+mdZx5ZGDF/q5ojtZNGcYZc9FjjiiMWcFnMMj/a
f0TiRdU+nMOYSee022I6OX4h9WntoKjSUkuH15Vg/DSo896G9P26YGc+jk0D8NdR
UGJYYg7FGIcGWWCPflDjh7NEsLjRUUwXJHkG6ESTYoKOdncjXVOOkzafNUAQS6eX
9gtv3ZWbuwjGnwXFyom0cKwVYdaiCieyWKuBgAZBl95bntx7TaDcmTFGejDpMeqf
YXD+rQnsAoya7PQuHqgTqOS3uP1LLyUXacbWpRTH5QtrrHxEnBPHv9PFJvY9uDus
UOnJJBgdyDm8G2J9ASm2Vzw2T3DYi4b/zLgrsO7YwacQYs4l3Auh127ynK9iAT06
odBfBz6UFDDZQDte5F9cNhdg7YRTgQ2EfzQGErp+tEj1iWseys8PfuC37O8U9yHQ
VZOLBNi6bicGaLWMEAg64hDDtpdtgIC3+lySe86OozN/h3HDrbBG2o60d1sYULbd
N5S5VNH0D8qLQFnnQQDJlKSCgMIhGpZocD4y0swgmcribhKFpn0WmEqACgNWdAVQ
UETWh/jvIvP1bu+HesdmEBba+QemwWnbgZ8JP2Nk9vrDIj1v0jwWqT5r9SWBIijU
UTK4ohu0y9gMrMtuPXOGRT1ROUKlbH16J28wSxFCF84PjaPCSqmh1ANvXnlz/zkR
NYZZ7NLZfzebX+v5OQcbt5ZYCT0EpOOL2ksT9/Jzt3FiOFKm4IOa3wHfdvLWX7GX
kdrIzxu0UoBP6wvy1Nt3EUU0QsOodxgxuDftDibqssJT0DgldNzA+MPhL3X3JdXh
Qv9PuMzUIS1bVkdl9edN6EWTI0huNThkD5ycRVf39YL8/22q43kyUHRorywGfFrn
R9l9XIFeZlif00kQyNka8PHJgTk69Mn1t6nYGJH/OtptBdL1ZDTDi1LyZjPZ2gMB
Gj+z2m4W1qICjc0UkidRKF7VqkApVqmjQhqcr32RsbwFCwvVoFmKlody0/5M/ahE
xm++6YgSz4+oke+vhxuGDqwAsR47OPkLuXNK/HKB+T087zjUcjfeyKboN3H9j+W5
tMvgBXTe5DOnOBKGhAxaj+vNoPRW0tgAzhkLyWp1WIirU010Cy5+Up623DTNSg5X
5rvpCKBcgEW/dYhsiLRpfS6UEmx2XCWuQ2MVCGWqUJ+BTn6gERLjytTAYXwO35D9
2xwvL9aFq0GmG88+QuI+Q8+aGo2S6ti5f8ESemKgIJTk9OSR5KYPBYS6qJBxT0Co
WsWk+1P92ytQ1eX2sFdVbtTEKLt00vCzH35cTxrFGXUzOR568q46YPPz3/AJmy34
IqZJNOwD1GUXONLHHKKdH+oXRF6jTOhbPTdX7Wsv2kB9lfqP/ubQJHs+9Y3m+FYs
SaXASNK1oRGtJXKlHOTAgqvQYeSwItaR6ciNsrSguDeppFipSmiBLpb9wqV044q+
E3mYC9X/Psj3T3pwtGMgyzC0BgHub3NZ5MIXNnpvopY9AEeTjCfMnvby4YglCNfY
+4ZNYI5drjaYga3IGVcdaE9soKvmattEqMIy0qdhEXxO8NSiishwT4O/xFby2wJ3
AKiMMHM+A/F6XQIpIQ5UZrm6UP4JvdblogZ7+ioSMFoBz7F6A2E5VBQ6kzCq601l
fqq73/clEDrW+pbmU4u9t+pNigWVlAE7Dw/7Y5rR6P2x4o8eaIj28NtEf4bVONoO
CTn+/5zfklNtvojYc79g4YIr/maHy4RhLP6ucOzxKvZZi89Z2yNS5XMXyJHwPbLM
KhNqsxPD4gzKIlJLScjRAz8S7/4q+vnBkaAGhlIEXZaL9vuqbW6kwSwa3hxcnFqs
ge5Ey2+1SoXxPqOoVCG/Yo9A1QRkNvP0I7rLAvDKpdha6g7D6nJ9EqY8wDA4NWe1
4J0yMwmlHcW7vVfOHWs7qbITesvTORXVn4zLXz1xqA7W9NFZS63eKO9NVwopeL3k
UKtvrsHSB/WpKyKFNxrZ26g9LaseYhug5TuL9PkKhiubGf/XjgzDfj4QiCQRboQ8
kR4CWCBRh8Rmv024uG3atgdHL8Yyfb447ZJxdFA9DV9Q9TcK22WremoblzsEj9UB
CcZEs8YB2dsnuzuF5XxOzrSztNvl2wmr6IUYxkgvN4lmNuIP/RTZoCpEDpsxVzaq
m/JdR0fNwTYi/i4R4Wmvi2ljbCyoGOs+uL+QN5xjj/5pny+tkRmm2K/52EWhzmW+
jOAyCgJhuTIK2Rd8WvPbtu5MxngR9E4Hw7U2WxNzIp/LtRBmASBeuobhtdeyWFc7
GICMmt7aPKf+sgOFY4zlntpFYQQLOw3dJYIPgCoYpo91CIEWx0YDAOldw6XjwYz0
1hTueuzwpNBtS3NbAk1zPOH1nIWEYkKZEv4A62QBLxcU9ZAVtEHwjaEHfkCRlyp4
RjIfZp5fPk9mPdP+YwIzh8FqX3wJk3uL7xw119bejhmgId08llJwInIkWVnOGyRa
gEP+a5FjLIsOLLTt+Iz81SootpTezUvtewVo84WfsffxPhuFXgvq/0lR2grn6kkG
fdQE39MXSEc1Kx+x4idzGNIJTsRsjzny9a+UZoF4kzVEsJb+80EPWFFXWMALRPKb
ouCSudy8OHqo5gfHU2+NDXorlvxs2pIelqMoZzdsrE+7hEB5vcRIPe3Cp/NhVP2E
iPz8PaUM3LKkd5LgSc2x3NbSIwq4mYDCURFGVf9C2JNwzU2lU87ncvJtX2yXvXKw
nhY2XsY2IzI2yqBLpyxjKMEZXXmaZXNJjwqLM/HMqkqhHfHKYu4F+wyKN1RnmSnj
+dzsX4qggcen6jjGv6F+w10xzAxlC+dc6pDt65APch1IjyqxG5/TdsKVBeBskOWy
py9X8sNpvXGcKBdoe0Lh0TuL/KV2NjwPT5GHpLDZdEwjNDRk2BmStirxqwQemDn4
u30pNkaYtv749mCkZtH/Rt5g4A1V1NHWQge8QXHYwLmAHtpxaRSxestZvoY+pcQi
m8/O4rnlKnUoaByid4zMzUpTxQLjo/sP2rfC+GE/tshTQBMXW3q322u+AKQwsXJV
T++GsVlmdxYjuPZsMXXvjK3XjjwJyxwVwjCLYIU9hXgFNKeteMozPnCPMRfscm65
MnaUB+S+HO6G0i5F4x+1UPnKFMY2dOb2/GIPmIOmmG2SunPnRxcA6PBSRLUAiOUS
DrLM3muYqb6gwLRlHWn+8cnfDPQnZp7R0OxJP5NRCtgcRXJKpD0rY/noTXIrpoxV
9Pbhc8yjtUhOagK6r19c3YvvIkrjXNRCIfdAdTDXCgiZ7G8bv1lcr0ydMmGXzZMm
2sLQ0oZUFUbPjlTEQXPYIXZcPfL8iHQv+oXw38r+NPkeq4SPfp0szXYe9GTOGAw2
YJLLKL+4d8wDdv77WweypLMpfHZtILnARbnrlCxD5lEjZOCFotskos3DkMi8ozp2
WYQ7TYHs5UyntZUGKpG8XeqsFosyHQAJO6ZPyaoNDhDIaNPfiAWa/SajMzy0hvcI
WTBEkh5OKMM9ulawqzk/FNkWLitqcYx0y0hOScoYrEseN4/8Kb+uY27OAj8xjCDJ
cMa8F+y0yuBXI7u7mFnjhwQ2G5HbM+be+ReCFNjdZclvBm8jP2f8HSeAWbCEI6uK
cq7hknzIoRchD0wM3o0lSsOBsgLcJEvOqiMHmalcgMQWlOnOPBbOmfKpGnLO4kO2
S5v003OZTP44krd930jPszvw4zQTxKzY3k+9n4wrDbiR9/AVgMm0WflW8OoSQ0c8
aA00O0yTpetSrFmFZ6PvDjCBb876DmrCUkB8jm0hkEvo0ANflucztdQwx8nmdjzT
wOd9uAJeLoPu4CKG6lIPecyRZWYx9GTupMJNpibfvfYSeowTALuizehXikQhv6zQ
MTf1ZuOuP5QBkO5qEYT3Xu9XR2d0vvfPokF6BBTcS2lvc1/1IudxStnasB5unVx9
0RicpHRUlAEWfimVFuCjDATojAnqbjza7QgRrSRIAZ18QWj1KKnpvLZbHas/JRTz
e7L+PfBFKdTmqAQC8nAZefLfSLtgCkEJOOCcreFK++dIzZeVO37JDHyVxJVd4PwO
2d/zkstAX2VkJRiD6rPXCYkUuLfXR5zP2S8e3m+b4DwH8x2Nj9jPIo484pl4h6YW
JMTdU60OZHVqIyG6M2rKv7LuWB1ce7dBvnPgs51lokCA/fYlrRYthV5U8+I3e3MU
ukDuzZ07YrLmlPnT0rs+90w9ZRjgGctxoLlxR+8RxsSV9UeIo3Y4QpHPgye2nIKa
HOliL1GJzNIpjY5f6brSbtzONG4XtMDos+FOvF35TXEMsqbcqb2iI8gIVeVc3Id8
spW/Ue+zS1rsknlepzFdV9BtxzA2I50bhQmhA5HA5H6cVueSSn5D7U2r6JLe7K/w
IhchUA1gjMKeUSD2uOUGazGxGLzWsgYgx2fsGns+3+Dn+M+d5C6kcKoSYm8V0X9K
Awq6my++D01ORifk/DPDDb1DQkMlCvrB9OH6jTwM+h9HhpdCZvQb1AvYKrRWcx3h
iY2eUJNJXznw+Dok4eYQ3ka1BU3dYDX6+a1ivSsVOxJYijtE0ZQuYkDZX+asPJ/z
AcsCE4OGdLJNTcbvEX3xVpdYu4KiF5uV3ecGXkm3Q2Aj4PLawIsDDTm9r0j2ca4C
Ls7ECxQzAdYbq1MJ1X5eUmHEn+7f4AMiOmnYYl3cLQwgpKGYkbvdaXX9gu6no2fV
8pp1UITUS9F5GdOsSNGs+Tdy7zaxqKbENqNbHVJuLI135wXp4c7NDWOA0KxvoL4R
uN07VggSsUyc9ko9hqRpku9JzgJUc4L19bU+rGBljbeYiVVqstB9DbN+c4f6FAXp
RgtlMXNVpXi1x44pqECEYceRoQcNlYUnOmO/J5iPp88V2ZxJimH5JIYiWdH3kuvR
rezbZrlIi8MZpGkyd6XPyTEMP0JP8y604fqC7spYHdZyhCVLa13Wd8zq+/RplU6x
54lhK/ne8APxJiQiSqYXZczmFz/kuctOsJqvFF3ueFSae3nDDaM7+HIXcLAXchDI
TKBTRmJ1kPUaIt/xjfiTNJ4N0B4iF1SyfV1mvjybU4JkMJC+7/jdjKeHHeIFhkGO
mf829GyH2udxG7BDSHwFsKs6QWXT4vRKy8VgWp3egwt1Sttw0S6p62E1gvL0cnX0
+RQLE24G23buf+4ckFl1Y7rDvuSC8jbp+8Z3p9ztJd897WrZkZKpjrDi7HdwaUER
PdwuelzS3vy0c4MRPn+Hg4ZuPaD4acII6ug1QZeDUF3QtutoiW+1KEOrQceslnjo
ABMLtb16f9qhl4DwKrCv2VFWhZgNLSCfJHU52NLDw+24TPEJwI0SYj0kQex6bupT
MgxAtVLt73p2eCOMm3DPagnM/ZWFcluVXaE7i0GGGNrfUVKMRYAE4+yhBNSlfF6O
DpHU64kO/SXiWB+MaSxtqJ1vMLmmXDjwpgrwZL7sier+lbFi0jKkXGegoy/1V2ht
9FzYJ12hEb5iVZR++YPaFCKEj3xrQV9K0NvRszyD6Fp4t8NcIo5QNQtkygrgFTzb
EVzNSsghzlTAoQTz2NoQ5wnKdrJ3xe9b5o1P6felolBiP7+V4qrHaCR5umCsE8z0
vvOWnxTXsy1c0fTPGrVvXmdapGPXSF/9jymMVFcGL+edXm6cRrpeLjXk/64CGEJc
yvYjoulKY15lkAbHoCDQbZMl5Ul5GQVlznoaxHjVRDVaHYUf90c8GZLLxzCCBDMK
Ud+s6UnA2+c+IgEpchn8JCrkXvlzl1Rm42NqQyEWo9UaF0x5RI0VTUEhhYj3REc1
sKi4mkxWvl0+G+DK8Z6C7IFLr+jl55cEv4ziNMVPcevlZW6rod6Hdzf1Wb3gojSx
aCfSUzH5AzsZGtil3EGI6/GYm7MW+6mo4Za6KU+/+lXnpg2p5/8EVmwW4zphGt++
bdbD5usUKAa+C0yTiUYTZZlbROU3Uc6WVuIylR/PZPXfpbt+KHgiEs98yJsx9fYj
5EugG1cuAcNs3dlwoskrEWdcINR5UwyRZi/LLiDaqVnHkQIGhdgo9fNhxWlFc9kE
9fL4I9h6AGhRvRATLGJJ+sLiyhXzjNHVKlPGypZ4z6MreLt9nQbv7lEtbIsmdRnD
ucBBgzU5zgrY8t3FAXMPMC2i57Bk/tY8JegOxtMKeDD9LjqgxZi9e7LV5NfeLzJT
WEemyToRXQFn0czAqaDHebxHiDQWsBFGa4FPgAQiu6ljzDobq3AbfSUjZH+ziRSt
KKiTpzbH8FUWrTOWicL3jE2eSPFb3UYv+qHRWv5/+4wx9AKheeuq+K+PZ+TWG9xk
r6tmQxPyf8K4TdlXjnK6nsMTVIkt12WIBDvzMDsDOAkR3vIv3PNQE5O1JRGQCxi+
u+Zo0L9UupaDjVOLIePBdEa4+RrAyZeJCSRGZLHKeciYx/V7fgGwOc1KL6tMFaU5
CFwsXJ1a+7rf2Wp405PW+4wVyAS1Kkt3L5DZWeEXuu5oyNTRuBCaWxT/U4iXegAX
6lnbvJ3zyqByHqPG0WBaK3DSEOdAWmgiP67VnHqIS6hI+pFUijY5M91oKFIR6p5E
ChHZpesoKTroXvHHHpdV5d164A3LtiU6HfS/Ms076dSir+ltn823ufbK5bKDbhFV
Sw9XP3Ce7DVnfhskyh6BU7iObjmzxj49s/zYce+JZBhPs9HsLMiy0sMMkGgb5Z4g
HRQ30sOG9CW/YMl/QxgMDxDVvUigZddPbVAj+eMNfewGoSrN656jVb3936BQGkob
MLP210WHkMgiBSRHGUhaUgDAFkZCwOrnDBXE3hVGpOAoqcGHqZaHyz+pIlqyyMrf
gI85yXwhCTxt686x7c6rltB2gQl0dmKb3NVmNx6aHLj17PfujZxlY8sDksrNREEk
I99WQ6uxanaH9MKTrfo1jnjuIcDHxsfv66lc9w/jQHUGMXJ0mV/k653pl4S755JI
zVs7ztVF9eFnxbs1PesJtde43ne0e4Jwx32KDzBGKv5M/RglfkxwPMqV9kldi/yH
NzGw57j/SfL2g3Ko9hXYp5R2XO7qMLt/ul1hHmchNRPhiQfyQ4IQMnMSMuR6yHQP
1exmAtn9uUkw6MGpGCAJ0I0O2Up4XUB6Vv42MEIIbWZSlnPx5oUzz9ehHPJLylIr
F3QizC+FrWGQwgE2jZEIC6nHffUTFu/SP/lfojiPc+DNrP6zFo3X/SJMs8z/R5jh
5+LxN7VJn5WRuPaNnC+yFhctzpzMpt2Jge6/0e/52upi8mfshO0G271RKAew5JPv
hscYhDvEXbFzXKpU5k6clqhkC1prkQIhey+sa+MdN7QP/MGH+3ZNJCVBm9zQNiL+
qe2D9ObGdr2PB3VerZaocf4lAOTLeKFbSTZfifxXPLV/84CozWBdC6/C0261dD7P
NqepcwSReLJs5v+Hn3qFHKp13urwutcj+FdG1+MXHb/ZOB3JqXc2s3Ii0lXGpMOH
rzeBQqvmX+wKGIuw53KaYWfDiELNHBuuyc9vYN6imhjnnr76cn/Jn6ODiQ0KRSjc
2SLCAOJ9fiAXb05bmCPtF3ATi7rEZF/crR4JG+t6SfguyfdQAAIzlQlcMIQGnclN
NBn69UhbvR91hSTkBnAevdgWF5U1FOWS/fqvZ1hQ9EdK1sj2+c3Jq5oGBTS1foNy
EpuoY/eKbMlFprZygqUHOM/GBy1gnRfY4JieeIxN5f6UX1GsLdeeVGeXlwhT55V4
UWKoK0KHhbBteMdhJ4gyqMm5flzCGBquUt/vrUDaR+IwNTIot6nSuqjiphOV7O4N
zELmZSjU5hnrsEAZlkznmdVBO2n57RHSWh+aze78yWpVZ4Nh1ZL3E/7GoFeZisMW
nPT94Fd1W/nqOKyJwOoL00yrbpfSYo0wbMqwRa3L3bHKrhDA4Qq6R7Nh5nLt3FrE
+rtf9DGJQKqAIsurKGhj9sRAgUfjg0d4kqAY3tWWpL5DB5HXCnkxAw9CtK4v4FqO
RFmEJ0pJaX28XGs9JGt5zHUaZwYC73J5+tU/64VS4oqemmTkv9WnxUjugbteq8/s
7dvzgtzdWbJQI2nzEMrZSI9drGOarLdzBKL7cFFSSiNq7UEPYxnISi4EcKWvZdSF
rxhwrEFe8ywYKhcBOU2jMDLc+nLvsgP6TQPH8JnA1gda0NBxBIw4HhEP1x7YBsjK
mhiQrACujEQcBG67bjbT3bnGPwMB7LL6TC9mabbE3W4bf1447CfxtF8BVFrOjK7Q
2vvqCi2wlDVn7SNZzUw770efM+SX7BvgRcL25z05Z/Qa7ZGfmZMquNkDazJOCyzL
m1+x54rzq29NAQlGc1fHXIzvtFSbnSaAQLRQ69CwBHzZXN9BQPZco79X/F6hx23u
tnbUVOfd9t9kQABEKDfb0dPV2PaXcoj5Fj+1CpE2LAXWXfnfBgHa9kbwc7kevf5P
cpksky/na3dv0EuFZkLXgj7dicfLntjNlG88wLvF2KOemVUOlFxSSdbBMraQvW7f
6zIKeJgMfFn7bb8KxFoScxlx2bwoZY0vTMGF2Hv7++UgMxlzsBVIBTIiraQKCGCq
14j/ibFNmgd2oKA8gba6UscTjW3Fb9RvPpVr1dNaXPdmfrVhhbtB2dPQfZvlkdTi
oyf/3gGdLiF+CP1FQQ6ORmjh6gkd/Go+jcCKoY65wN83rbulrfPxC5PN62Bee+Ae
P2X2T5x/c5XlVEwU4M9WPhuEj8TFiLwFnDNRf+jspEs946C/N1StIRel4Z0Jy+N4
8qjhtvAMUGST72FtJLZ7yohF+UHhgyE+aY24/jAkV1nFRzs2/O2l79KpAIAe+6/F
qJeHAPkrQZHDyL336TplfWVJZTYPsqFu5xazCEjEhvKS3uF4oMRtJnS8QUzYCKtL
OJ+FAnlCVvy6zm375DUARapg4sw5vKCDUwx59g8k+48Y/GaNwpqwKjvwlLpJeUfT
7iGB/PBWMiXspQp4I9tVg0Hcy2JJJHdjmuQ1fAyBXTsqLl7CpCLsW7Pc/+XJB1zC
lxUFhI8wAn6mop23NC44pIP9qN95Ixwaj/VXdm/KI0w4/SjSZL3QQ0LWYCXFxpRg
c4XcQGskVS8pD1aQ2XOLvr0YPRbX0R3UGdoE3nTObzXUKHh7tEQSvBLjmaVWfoKx
Vhm7ibDfwZQc9Ipy+k1f5ae2iHUFzOT52MfJB0wnIo1mwxhZgBFDG7vRUm47CV9v
J8aqT5zXgVJ71PTePDrugiPPGuVFih9JYrw2SvhS9w7eBXmqQzhed5xp1WSydxc9
wWehT3RznSi9s87z4jjsy1XM+mvglxtH3+QE711TJLAKJjF7j9f+BoNYkNt4q5N7
anv651EfFbrrAPecvCZcnZh3LYujaiDD229BpsfzlyWRuw7LBV64nfAx/W572RZj
HaQrnQ6e+TqtRIUMOcvSDwsNZWX8YJ3yyCx/m33/C2JBnM+/c8dZN0VmuS22mN8q
0vwGj8z+ha5kW/+YTvJKB8grUbwSkSlPcgvvIf2QJ7e1piP025TpgBro1XBfUSPz
gnNOGCBWbA5l4qkOykiRewUCajsi9ZeejVxt7Gl00fDMrFSuhqf7Ji59HMzbw36t
l2eILrTVBtBY7MvZ6aU9lPd+WpjNp//9gksvmpkLuQ8EDO+ziGmCjQ80bdBhK/iQ
uym6+E6+MzYDfvjXU5l6JWr+LjoxfsVFME3/psrSQTfVusXxR94DYc2idaZGWHfe
V0tiHoU1Czc8GCuLVho/x9bVVPAWu0SkylHG1e8+j34mq93vJp+FHQX914FpvZ0i
8ELpDqbkpvlim2UIlwzsmWJ86BzDpZMJ5SS1O/BOzT4hNYlGI/IcwBG1bwLQEBBc
SWKNutyPRPEvSCEnhrvLSA02vnOmUst4n3lQ7DBbdWFb+nznDM9ZxIka+UMLFEQo
72F+JdIm7EKD2agMTiYuGSNfBut9G2aQcQqqkjnFiqaiSBM9Ju44qD6KJhmmC4b1
kxt5CEANzJ6QMqG721fdFmb58rAW3/S/eupISFzfbocfrBwThDjwjf59Ldw2iy0W
ljqOkl7sT9PQYe/Ljy5dawtkwWqahKRkoLNkM4ocx5NQELBF4kvcC6F3UI5eZSTt
yB2C8hOhVPyR6jBWIPKZYzqPA/KVcalGYQUI2ooqM1bmobmrCc4G2uqp5hrjCuEi
ljhB5/IbqnXZKB+8FZ8kHlilEIahS+4UFLo0HcgEROS0KdaCiuBXeyGFdCrRZYGR
LRDNSrov1ZFz91tU4otTn4q8X4HWd9XenT0g8KAW5+IObALIPW3cv21ZCn+/Q9UD
cNIj8F3XIKWw+XyNFhbf5fijF/5tVuNmv2PZU2/U+gxzwuNMLvBsylx3AlhagTx9
140j0dqbJ/6Yvqv63n9ZajoearG1VY6gYQzN3kFdPjtYFGcD+ym6K9PDrZVd8PbR
1/Q++Yb2tQnjPWV01KoyDakqtl0ZJUHZbnYrCB6nv/8nLS6Fa71k2pqTjN/C2cv4
808CgqArn+7uyWd2hoGyF6oGc3LJwRJEZ4A7jM29J8rn9PhSMGyJ36tC0huRNMmF
cVrXq24nmIqVk+Yt8TUeaMIFHDCvHDlABT93g2rZlGDyrC9ZGRbYJxITJxzbO1ec
piN/7cXQ9dSlhC0MkcUsN77muPOpKcuekRLJ4Oz4QaKgyjyaoFo07uJJXd0QaSI2
HzmFCgRmbb5R2KnMu+XgNT9DidB5r6eAGUsIUONBZbt48N0Gbv827/mr3WhvMga7
7EdtXVfcCdS1jhJdy/UNYm/tdF5e+tYL2JSHgcchvOPETZE+u+NL17FVAsp5A0y9
cK2v+WCUmzugJ9PgLGEjQw7vAOACsrPhzhjYblwVd0hRG/0qZ6sXrCRlx5Q4UYG3
GoDSFYKXNpiNrUjMN45rmJVzJN5ViUs4fqKGGA8Uw8dqFJZxawdGT6tECMvCx6Te
dE1Gbxs9lKslCsyDq6gae1JVYfQ7Oq8t775iETNt8Z691d45UYBSGt4/BKM+QMlR
f9UqJyKib2fuqaqSiK8M//MNNHLE6R3LzHBbwA3v/phGNUb/9Jid7IrUDyWrCPc1
qj3p1GbBryfUGYoqxc8G5Vzh4SBYdUzfi9fzXUWON555KiMJFfGSMNhIoNYerWHO
AyUFgs3t/1sZzOx2RBOTVGS5JPqfUNvu4Gx/JQDF72xQ4dWfKAo4e9iTrj/mLRoh
nQ6T6DBq6TWaZQ+N3y0Azh1MsCqZX5mVIQeorY5H/wxKV3qx2MFRbBzRlrT4MAoi
IO5vAro4AgLA08/64X8n9WWs4jgc2+jDuGgOrJxTCF9hxPrLQTbNVKLUgkLoHDVa
WgH4n0nu+hC+Zw/asMdBy7bTjnPUB6wZp3qkp/LGYNRlmN2OsM4s0DXe96el1gwJ
CrvmUJTbbE4hldyTLdNjPDoemyxwJpJQ0AXp4DvLk4kKyZxW06iISujisUb5Jw6/
ij8kxlwyarbHOMwnHWvvexMG1C0DqF4fn9oXL1rJM+j3+6cYXsTrXqwjhz46Hk8n
ut5FaDqv5MChb5iRyeCL3DmI3AxuF5bkpdRE/Ej1gUC2/gM112lMn0FOVm7guVx0
cobnzriXc7oi9YOcvv1gB8124jw6NBmyH68jikATNZKV0mS7h2iV83I3/L7IpEJx
HMAKuJtTsqrqterXfvDfWO3beq4644vl5XlSGJcFRsVtks44sf7pMn3aDifrJjQm
7JxKnE0Lk2CrOBJxVESjrQW4n8367My1ezJcDL3A9G+Dl6EfcTqLNoIN0Njiqyby
QiatB9uRtkHbyz/P9ZZ0lSBvPAxEktW0uH5UpAgNCeV/gIL0XMaDymFTj03a+DI4
e4O6WkQBJ+ZTuigHdFZGs2lh5DSTeVFMRNFaWwzAgOwN2I+tVckZ5E0vV7SwL4ds
WLYfq9Ed8TS3nducSCokNdt5rTs+AVYTWSEINZLJQVl7GIESgXi9SP8M3YkGMjNR
BePx4qpl/MR4U7BYMbIYaWbUmKYzqDx1Lpl/97FrsK0tUtPVtNmW3hEOG59fjjdM
mrVCVMTSgPanSMb/S+XpMhUeELbiLKT/ijI2UdFturPAH4htfL7tCPI8s+eDnWFp
ZrDd1qTk8P9VQji1EcSOhBgn+YS9OSfzqu51vyF0GrU/d+Qe/d1kh6mTLM22blb3
0rzO78+0VjB+bamP16btlJJAby3byZtw5aMXRZgAsrhq/Q7QIxD8W5V9PRgdjGDa
dpcSzb0p1cuhX6ktCHDKUKeXrazGWAhhmlIqIoqXqqxLztxFCTm/GG7pPiCM4Rgp
392h4QRUh3W88xaixOaBFJFw1eXJmSG6MsH81Klx35m46tlZbwwcFLSwo532lTMG
EhNjJfy/v178LJgOrn3TPOjPomsvBpQAKv+me0eSWmg7qNnvsTl7SZCwaMkpo8ZI
SPmvoUuIFEzp6XTeFS9/RBr7Dj3Bx3+33PfDl59RmzhgmTH9A1c28IfTUe1MpHbz
UvLGUPgTIr+OAFVPisaKLVoRUUHkV/8DaS7HdLg/yXsIBPvfBep8A0bl7DOOPqhQ
2149Qw/s+yDc8v/V97FNeSWm/2APpET7mAocXp7vmI0m7Y1s3GYmQYxDraD1+RUm
Zo8HPnDeLjaUS2uUWZ2Out33yaeRV3G2ioFFmv4QIe1Als66uQX+6zvVwNU3lBRX
OIYXW3pqjGD/m9KMXv8fS0/1vfH4deFqxFPsmLuEjxHJLRRsM/UWeFfGwOS40YBe
GcrJQoDYP1dE2gAndgyyji9iRiDSnhC1983Dbc7vzUTXyr+r8mtwVBopFEEWbBbq
myZQhwENLXJl0O8q6ReaFW2zYkZWAGrviBBQpoiCxCNDr5Ve7he7Hf2bJoo21g3K
3EIbovR5cG/mJEju/5FNO2+8lkCY/0ExqdmVT+m+diCx10wceM3WANYW9/lJcASD
KvCbht1Ppi6lGWCda+Ab0m3iQAneh7E5/Ijk++0aL6+Fm7qPK1OpCrQjx6S6KYqC
IvUDTvbYvuBVzcr9VMlicCGkfkLLxCHdgrrQR1Bhajgl3TP56pdYp3/Wb/2LrfNF
ooeOO0Nr1O8e0s4eU/acPr9U+ERGvntJ56rGJBvtEns9ji5G45jN8gFcw4xUPS/e
tmlSeS3IUXsIrsWxbh95wUCqhQ68MGrleyS7FGQjHExVj3N3xdK0X9kruVD8b2vu
69GQ283pntK5JJryB6VCuS5KmIE+ZZGHWjXOo5nirpFagY8nkIZ1WC1UveaUyNsD
naaKtbhPZaEjyETDFNeM9T3dih6Ugi8eN9Ze6YcthChLCubUlumsMMYTJiNi9bhc
c7xZq58XDEDXTOZmRdKoVD0sfXm9tMExZNlWU735EeFrQ8PeYRLM1b38B7ATry1v
rmnNmq6r5/CL4TvKr8G3JfddQdRAy74w4ONSTUZhzMAurQrwLDdVchpIMVkqbryn
JqLLMijk0UGyQxqldI8xULG1+mdoCxAEo5OyWhKX8aJ0ofNz6sSQ9/e+nsSmehhO
AavYFHCBc21scwpVYKTLRa+u0IPhftmUPgdMG0aNmYH5U86LMgDktnzsJ95YfWc/
UHpi/i3RxTgyVQdXFKBUnbycNEdrPJY02XKQMcSRug1AE76zUJc6cA/OY+WSoae7
Qffcdi8oK8Hi4EdOImK1tTmYK9E5OxFZ+GZb2+K1HiR2shVNsi+KmFJRXesHrmx/
TaInUC7lig6Jp9NNB0HMkercXPw8fPs72pAbk2MWxLB/4VBEP2VaNn5QOJqz1FYw
ZkDlxXzZI94uUd7HbQIM1vcdR7xnmpzXeapo7foxg0gnW5/AaslT8wqkKc5Ikc82
a+oXaUL4xdV5L7u49j641mu90ha8HQruFedEdRCvvgoBKjI+zungT31pmo3zG0/w
jDGdRWbqRL/v6Y4NfM6xGsvwnFviRjuo4zrnE+1tZ/v3RpuhvA9dbr47fH3E4DPI
Ml6N/23c3vdEwgUWWJwiCD9nWHtuOsRwKxnhm50CeVi9rlmxsvj75LzyadugSGwU
URXWxL78rPIjvHg8XqR/F3JxWxcGwI4yQTXBmyo8F55mcYA5ZjDrAQeXb0hfmPdp
7rIbpiWGC+s/peRJD8SNcnhHz1aKglRFcz27Iz/lCwpYhiBurAm9ZNlf577YpthI
rDl9jTIFXPYdWEhDB6x3lLmllATeIU7GH+GrJ9POwx0rJAbYFE+7QYXjn5PuZDOY
6HhlEoa8hKviKcHbtiqO1wUTxQbMiDd4Cy2HkbGi2btreUHa1gnob5fRWUCy6uPC
AKJdSfIl8ec6zYhl0HCerwQmgHGmNqnKWxTAPXNU0I0Yr7BwEyBNrpYDaApErxQ9
+7LA18lIdRr3ZxiL1/+HVZL5CNtA02oCRT+Dpbk3/TJuXweGVuzJzP2jIBQBnIDG
r938lp4GN1YhQTpUy1Fj3OFb8CvcN9jBcQc0Q9l//RAowAxJzv9jm3Hqhu+ATmEm
AcowdK0g5n4FW7qqaDNI1GoUnfAwfijMUIXu5EMzIw7TlGe36Wz/0Jt93ju1zgDI
zPeG3p4DtPEzcBmEcY0Nm6J69dsioDkPIz3j4Z63d3riP8DB9zF75xtTFIyQu+5h
8/1NY3VDhr2R42mpTzEM5h3o304D93c4aOO1Y2sbJcCAE0iDNS5RfOZQNCbA/S8A
nJxdxSgMJ40hjfVytyzdhyUIIzVfXaIE8Zz9AbOTyn5H2Mjw+Uj7gX3s3ZDtRu+P
P/zHR8f7OxKwu1O423R2Zv9ZsSlRpWqdXvDDLTZzeIFT2WcuzmBigTtHoYHZFXtJ
JMSziArHGDyXoIoPbi/Rgl+jVfrRAGzvlolAxSxudXqrOauOqPzx2MmnT5iWJyyJ
Dg9JWC+FY1U4XYb4kU9uP4Hg/cUSs8tCUhlhl+TDSa5eSkNfe/FJMItENJ1Ak3x/
HZjvDwSK1PoGhBjPmWG63XgyOZNIiDrBlqSkG9sH8TyDALDx1pmhfNL0CuTK4YwG
Iy+S86xYEUsYA0sldCbhQuENkfdArKqn2OgRy+FIfg8RxSuG4beY9HlnPyIJq8/g
I7xJA0n2xdgybje69EorjEItOIk8LaA2vDXBpIzyJGKQ0+AU3DjwZU6dGuhlogQX
aef3PvArl6cxaxUQ6TicC0cEKbyzWTCrWGw08CaRwXB7sUAfok6Sd24sdNUSPtnT
LD6mKhQ8JYF48cXbShnl+FNn3RdrWnlGeqG5h1YcCCvlLmogzCLnmzrQK3tp4g0M
p2Tp2XMpg8+aL87g/DSxLBuEL3QQo6POY83eAJSoSh/bwe7CQzuT52A4U5Z/bcbG
bnp5NOP9xHtwDvfJcB6Aj2dFNPZ0u+DuMM5ZHEqlICnjy8IAuIBmDAhtJGX8SYeb
8qgUUuqiwjL/bkQcq36fRceym3W34raw6NBFAmLVT+adUj2M9RkO2qosdwap1ymv
AyKdgLThksDNMgsTLHbgnMiLCy2G5xy43+3Q6nnyG14AEFCOwwOZxR0PcUuwGnGk
nW+brtC5v1V28pH7iphpmMGPMSyaql83qnHzc/SLM6C2m+uNK0U+W3nmAou5kHLQ
70QyQgu5i6/VtLYF7g2G0ppfrpxYRj4GIWuvbyHBm3JDVOuD17+yITriK+i/7Kt5
PvTMJ7Z4NmclJWInb30RCT3oMCB6Ara52xworU8uTYRhQ31g6z615VJTFgqtIKx0
WjwMwRls0S5YJR6d/wpF1J/cCtrJ1BpDll0F4WhtzvxhfVaV9rMTu4ITzQ3WZtO/
0+ilceDBRs7EzlFMxt2G8IGN8ULrInByvr8ZR6ZJUI1I2orf1lIlIIjjxGLZFxhE
Yu6RvgLWNNVOBKqftFUy2Cd/1D9NScIV6rkKZmVU9XQbbFv/Vd5ONtQ+PWdfrAOT
30oYwJYv9+J9v8OIvQoYw1o6VFaVcyaNYbCEBlUIF7C4nFA8P3XponIr5wDjeZW8
G1akWWKebnm6+eEhmw0P9f7IBW5lbmOAMR5SHrrad1o1sJqMQlOcGnWIOszegllA
aWyFjjuV/BhyWzqcs266Gy+pWhn7l0oHNLQAId8uH+nkghbRR6P3Y5U2tYoIZ5XZ
gA3+YcuBGQ33bc+oYeHvFEZXPi1+fCOO2D+FmNc0/g4Tn/cQKH7UgspnjOPQDtiK
83gbkm+YqWWtVuNJbevpaQzjLhqpRZ7C5l2udPiPdAVdBlXYzGEVHQ1IN7/fQA0b
mEdUcatO9rIfOjyfCO5LiRaFpsg0vrrPzJtjMsyJ9Jmn5hh56GQ48bYYQM30zcgm
DBCp2KlF2biBp9m63RIvDwlzXpTW2LnYQqEYjXJo43/uifuSL/skCVjZ8fWUBimA
eTukaCspN2fRCxyTqJPlgtdG3lFNoylSUxbPVNi/i694ItK0K8zlbhguCrPZFCve
IWEfiWGYSR3ryw8H7VL3wL4dDuW8G4uN4aq98RdPvwxHrusK9fN6ZUxwTPvyywr+
gIe5zTGUgmw6FD746lzkoS8HsusTUxk5NIrULZp8oW+4ieKyVY3AsKIlospPmI4w
JNCtZR+KJkB3Q7iqPMoVKS8eNUQd1mbeqp28/vvPTl+ZxvkHScxfxpPQRo+ZQrhq
WcHYh8Fl66JvwfKVWJKhUrQD1F41mPsaJsGxLWKlPqeftQp278deUNLvt1C9qAn3
XYqZeaXkO1ZuoAL+VPip6d9UpNv2ffYBsesTTFwTPbr5z0L0KgNKOTagkhWBv+rw
iiKWLwJLC/Ai5W7zONPStSa4GOHIIpLim+0Y05u2jeTs9oHpr4NTTe1hJNUnnzn4
BgE1SJ8tTErch1EPwZj10BnrP1C8atKFu9F+FW4ph86FbYgenF+xmLh1DoDCKzX7
AhSef0Io5hmXsEMp/tUcv6FS3qXRWJsSVOmgc+kHDbjDRN4ed7L4RdeihGME8H89
tjsKJeLCuld4x+KPkjq/tz0n0eN5TT3qIIPYbrLQkHa9HvZq37vDxlDY/5EPiIqn
QGNN3Uv1XZOU+IgEEmh0KMunTJB7dLWdbfhQZL6x3g9eMsGO4qZs1TRPbWnFSIMt
NiRFq1CjEtR58LMqdLY5eoGTQygQagU2pmvzg4bOVYXf96cZhM2hj5H/2mCjaJ2t
auTOYSZG70ZG+x/psndGwUt++/UVk7hZfHL3sthbbtLF+2DvgIM8Jf6xFeuJ7XWz
i79fZm6+R108mw2ISMaLs+iPCqOLN3mNJLlrCyZ8VeXyBt4M9Gs/ND+oLSXZWCTY
pp5lJvdJv3Uq+CqboNBlpqRHAm51WyVrOb5ogVmtSgd8EcrDKPVD+pExb91TQMUZ
bMBv9PKfOKZ0rmtvMriaJAg0p1W+2c5kF0+9myJZ0PJJ11CHYSX9u1YSJ9QW0cOZ
PK+/2evVb7aXbpyo0twd/0YKbazeD351UPW5fzNjBUvaKb3wDqU46A8xnBQtNmj6
9d7fqp5LplKuR+qF4UlJvCPxqtVZFT5NsRtCEebq+B7Rp1W1ueMDnAqzZPZCLCzu
v8f23SKy9GBQkLVkvUhkKIHl5v5c5pHPI3RzcVQyICt2Ge4ZVu+b/fKPWWvtEppS
GQVddLlQcg+iK19LvpXH9fs8unL8vUDXwQWHphRQhqC7YZvqPkjdeaGwVjE/rbcp
l1jXpyjzVj+Qifku1dAZNsCtrl1CPiOYLvdYw71WUXViVRcM9h5XeU4BMqDpYjHF
r0GbEfR551DGTk5ogPqt22sVgre0m9De2aKqH28RSoLlWQBYIbKBMye7VbhKs6WG
kTj/i5SEcuMQawsMAVg+t0ItOc7YW4qFlHLOTMBwPPHulPF3BNj13wMI6PE3UkM/
5cADnAvkpT35jIvPk7jQFW5vM5F9cY4IlS8yvYVsVe5cXI5/DjK3drPLsk8ROEWg
nwWhCHHU860vx2X644bSVKb+sGtlrBlVXL6Z9CJs1t8nms3mWkRat7ZyxZafFnEh
tCkdbmn7HOBeFsOQ6C7IOAM9vtSCFiZBQWYt5wOBFs7h8rbByFXL7CLinpYAUcIH
gTVkUWukcJyZG2FSalW57L59Ze1wSF812HMUuCXB4i1lJQJk32wTwamkAF7C5A8f
6c6WbrYWzXofN0AYRwLPguehcJEbo6OH9qY3GypGDmlogzX6F6v0HTkR9ubIzHO2
2GTClHEanrLwB7ONh/TtGsL2UPH9TV7omNfo6eO8ysaOcYU2VWuNCo4Orcz3W2h7
BKsNR8o8L0UXuyM8bhq9vf5cA9V27bJKK3eKJUQF2uEYJFzyLMhLiYcTFC+fn47t
lpBbXSuY4HVWULM0FyYzbgfqO0VdNlCuMWEb2dVjEndGne6qp5JX1QbHbPlrWRBj
+3SZ7x8fBk1uJcEnYLN6JaYr94u8ZP86Ku26t+MdY4XeWD4yJorNJH5Qw6SdHx3Q
1lIebBlrd/V5+f3UdZ69+Ia+dDkhTb1xcIzAbEguLyxRwcOlbF6mF4y4uG+kLrQj
HQ/Ex/q75zoaHfjTgmy34bT9sMpxbQKgGcUydoEduMGes/lc/yyxk2lyzH6w7nqh
qG8TE5u6ITacK6/aaRRv0F5A2pNBE0SAkwVDsL+OZrVeAZ6TNMEYJOhg52HU78dB
aWk0wDiWN9qGmNFaUNa4lT3ctSTU4X7SkuzJx32epEvjj2XkbNkfRgGjdC6yeGAq
zTfSdsrzV6RSxlPxe97rGespA9GY1Jg1cU8gY526OZD88l/bbTQa/5uH282dJu+l
q4zDSeX1slyLkSy//0Ru2gQTmwk984mBc3R//Xw8MPAt9ilevejTdJqMiKzNi34Z
d0uZyT2q+4hWtBoyZGetqr8pg+b0E762/OcxuOi8W2N7jAdQIW5cLmR31DYrqvvQ
cVCNZHdK+VGPGMHkEQB2t0ofDr4aRMOsAFIDrKgqYxTG9rCGCeuhxXgro0zNdBuW
jzf/BLilYdCpdWkETbWISEiWyfEotLiFpfBnrSFGvwHt5K9PH9E5dTG+sDcM+U7p
oiWnbe6NbCogruJjs4/d4CQFhFyxoHGADmnluTI5VeLxDL4OsznVhCchlbh0ukd+
TGHQBfRqW8lXk4WaPUyvEznwNegPfPhDGKYgOcNFZ35ldPgRyNYutqnEDLHE4Oln
ySe8zo6O4Z66AKfExdNT3Z0H4UVmDiPceRDM5NRtVuzUMAjR36sqzoTCj+6TJ0s+
bpXjhcHeii1xA0gq6GPQWYA0sqFiSl8RYbmIfh5I0z/X0Qy8GEPitF+m3z4jR8/c
7aR2bTkWNy0in7DhJiJGfqhKWxU9L/dZAsjhezFn233SqqR6CIb/QyZOuHKb97tT
4ycwczmFZfi3d99n2lQbPxnar6GoV9zOYPogCygUD6zpeiUrbJ78lGHVFLQPHjOk
V1BtxDY+oGbY8vQLCnqyVkrzTYhDNENJ3ryObmr/pAu5J3K2Nq9+49clv9gEPRT9
kvCclhsoj/Y7eD/akTdma2hWHmBie8+KaVAKiKHaqIRZDIafg1MNeS1LsChgcbum
ej5vgJeCHIs5W7wz3uGYAmzVlU43vigIpfucOHAi4yoRcipvFnzym67cGIyW7WZ/
hcddnY2qmtRTDUaORMI1UVcvS3hx3qpMvx3/W8AsDDEnZyi1Ik/XRDcBs3LHGouo
jErKj/0TIiXvNtsKq3o1qBLMN0nBjfv8hdZBOvSX6zPow6M2JNAXX08XLNlp9GTm
mhbEZxRagLpYlzzaeToJICKAFZfr9+dOcF/c+KbcZy5TQ+J3zP/O7gcPuV2px9dY
P4kCca0cuQp1icxFYQprRZW5oni3rc+95l/uQkXpV7eGqL8DHMGxizmoQTsIzAME
KCEw5rN04EB74p52pY5D9/zEGQRCNu5iGrGghlZHGrAx+DzzEEnB5TzArCiC7WIp
G4jFXmC4T5T3wO/P40tdpVLB7ZpBkGOcrrBlt11IhLXe74FIDn5t9ajtxN4SwXem
INBdpH+KKluElp9BTu7a94XbgyG7wp/VtUSQhojQOTYc3s7yXOoasC4vwzdtnNx5
XYObhfDUnZKMafDk8L8lmwlFaJH7ePlgwUO2xBPUCo0FH38aVvM8jg0yKpS+gs4b
22ElFdTnNSJY25bCC4bxoaeVtosQhJzS66ZuH6XK3l9OMekF4KSAg0xXPxEHVc7f
QclJk/K9UkkpHeGpcbUL93Be2t9T6YVkxFdl20kEBdWVIyfCMDdHKc7gbtj/qiMs
BHojyRn6ikkywOZKv8z2Wj8qzJX1ajSKYHi8mv2lDsMbIb18Oho1+FPTwaCK2WTu
5kmpRJiSZVrFXDoL/Wioohd1DdRog9v/Y9cT9QufFR7wH2JvnHtjv1jZovoUOHU0
ptJWrQliYHe3C2Q9bX96O8Su+ReNpJJkSt3uoE+PpxOP6OVmNWGpz1VZ8Tcu1iES
1vfU+8H2xi3q0V5BOFDO74sgORWrKHM6AF8/ef4oAIcq1rpJVJAugSIvSvrcZ06s
om1hr0vSTctP33yujqWqfb8kpATgyFgM2EbE3iwVZRekxRQfx+Hc2gi34Pt4+Rez
ALmt3NbqpEcuCRIldeCkACInpIXFLWdKC1/Mrg6MClPxFyAeF4BoiGBwEAmBrwXB
DZoXenk4omAkIQPsEG0BC/KKpEqQyVQwhgG9pfRe9CynuOoJVY0neD5cJ6ZWQFHR
Q3HYSpSXqtv/qoGVNNFPWzOEhRkwsQwlPRpfJv1PVcqEIxOmULi+f4P4bR1CQlHT
hefHFI5MZeaeP9AMr9cKkXQYNIMHInQcKG1K8choJbyDIgR+IgqTDnDL9jn96k/l
qmg/c7oZEPwZ1ouxbcabsBm6UI2oV4WDGWMdWEauOibO3fp9FKf8F9eDFwl0moek
RVyQ9Zf0ryOgqldtqYm1pXn5nN2PNJh+2Uuo9vtRquRJU5TsKjyHEyKUIIiAJJdB
Mgla1Bi8tksGkrVqc2nxPNdSuvnhuBxFI1ux4eq1E++OqE69DnfWv9Xf59JdHKiU
v9KA1jxZfpcjuvfsz0r8V7kuqf1/us9076mKSPti07wEfIq1ZE6BvBTTqR2StO5d
6hTCyNF/gi72Rrct9Ak/8J0UPfuAvcH9OD3lsEGWojuwvjk/L3ECONN2BdbB045X
6k/cWNiG9IoDilOWiJDRrfg5/wUC18RihAgA7RLfDIRgrt3Zyc76q0OOIaevi2Mv
UydLOLE1Ya2RxKHp8ibwUdjYjWJJ8yu/pQM9YUKrTCP8ipocHG+ASobU/UjaHQ+Z
EW3j1vEIyxq5p2RZKcfHyHgfEWBtTcE1xAjKK5NBKkIXeZS4pnvX7Xd3AKjMQ0Gn
24F0khrJbk4UUZDFiW7AetXa1qwAQGNRHpwGPJe0Mwz4ACHo/iG0bYaChT4VPoum
qxuqgTTmsDVl7D+X8rcLJi+t6Vp74zQ1hDqmjc7nc3z7LIgcHvQk0b04i3QifGOS
+IcaV0ZLYAgbm6oFoyL05jAga0700TOhQuLSFZ6956o538jd6/AmT7vZUGmkfwK8
OAUcRBuX+7iSVtLfsftfFVYl8K4ZeFZU3Pzw6y1lRsimJbBoxAUKHLYRFUImNg37
fl31EZm7krLUxGa4kg71h8c/YAHKyzjb29n1KV/YtW/SDgdQQz0J1+EfdpqORtxS
RRAocqpAtSiOEwgfmmcnKAHG+M4R5fpvxK06IPYxmnTYuF7LCBg6AmkZwR0+xF3h
wN88Epp10X+fmdSVjn4oQ6HgmzoyoQp9txzhilAVOvGbw9EYWyXw0kyjugnDO3BC
iWDQV1Q4W1O/F5qqPwYiARaAuwTfF5IKoVtsnyZBZ64mbDVY00pfLgqkRWl9gVij
D51/Kz2oi2G+0CvYInIEEOtRfEf90CzDmbD7x8Ly2aPz4Z+lnjonTHo6K0P1JfGh
BqA200EqG+7KodKKYa1DWGFO8ucgqUwgWmK41UV/uoYAyXNyTC8YPlXj1TEtN5u4
/X/A8Sf5sGC/oDqJFovS/5whQ2RVsSA+xRA2gA0j0khcIb9shhMBxcR4aA4xCgfj
HufZARgb6m8lPAvtqNlfreWJtMpS66KAzSw6k7b6yd4YQg5Isj/M2TK6uj0K6VGE
F1bret78yPfNDCI8z3Zh/65io8ugacMd3jdG9Buy8HbVF39LqCzDKhuPpsLjFfPr
hEwhzuM+uLWim23ipsdMqmnDnP8mEN/MVm/niuPhp4Khh19N7p9dtaXVhMdgYld4
+8S+0YXtYobUU/nqGxKKD07Pdv2fZpeMwkICzX0x7t17KL/Muv5CLNrd+pvNq0Zj
tCXU/pyBLqClfjOjOJAdCLztf/PM3RdHsQpENrAwnfCVsSU8U3s++bXUQ+J8Trr9
DksitgZTlIF5PX3juObXRcxrVzMGnwZtQHgQ8pwJb7itsv8ezQVUjwreoeePlqxO
ILygaNZxVCmuEpFD3hKG9rBq6VR0vmYQJH4G9JDVqeRYWKnFsl49Ek71Tzqe1jl2
jHB96oAuWOtK4dl5wJLemPWgust4CmQ3pzbnNSuJXMtO9VfDr17nKtPduG7ftuez
M//Ec9uMIVrPvI2EY1WoJ8Hb+wk1fSAI8vgUdBRgNi5O7vGP4aXEGOqAgZCfVqpa
S3v55qqbpn9Ee4zQnDpK4oib+BuJQltV+hGs131zUxSKHEaM9rcAghwB7329+GZd
f9x53aogsyqyPVJm7T4o2Aop5Zp/1p6OLaBqJMOsNBi5aLMB/OcL2V+XtHqOERsO
U5LpJqh0Sc/viYdj2GEfYZ/i/n+BfXPtn7EK6FwxEEyrkGTOpvpmEFe292WvkObP
2/qxSvxWKO//KnBHh+uN0t8VOo7nbHyM72C5GqyuK8rhlGix6WzlhixaFPvmBE0+
dFxs8GsBK0rVs//5z+MG7klpUGihp3chnlMMARkvuFYQT9iQYI/FFaXoOwOS5EiC
UYRlht0EGYPi35ZwIbrRW1dppnszv41hZcAcncTHdmLrpGgIaODdgs0LwIf0lKl/
zSWz2qOdaK50XDfXNcQ03CcVlopjS9ogt77ZX9v9qEelq+NjY9k6M2XCfFJEQCb4
jISgdXMXQuazKfuIXBB9ARTYhjvtTEJKsCjFacFc/o2pr494/I3FCq7yIrbCtlsR
Jy5YFdedQomYHAL5MQ7h7o1osvpwT4acoCPzycN5m+jDiPeP67btSXz72NsXe8R3
UIX7sBssTuV25sJ0+nDISA+80R5T41bbzkor9QEzRlS3o6Q/Qwr4tjxk8j+m7Iux
7IWgw1aVoYWTm31MoQUvw2mjic25jKCVhpt6hGG08dIic3C3l2Ch6L+ML37UvqAM
ZeeNQAWkOC3XhQVw75pE0/k787vyyafzuI8YYKrMNUNKeG3WX0NkNJaOG0Xo0ME8
kZtNx4fdAwbcvKdgrYWlOTgxQdHurJxLZz+r613OZUYo7gvW8yx3UEbEmDTsMBvl
a0N7scz+PADMCjKzfXXGdcvzi1DqaDQF4olEr9wwYs084q6rm7PwfLZqnSKUfL/m
kjtEPMZUY0kHkA8WuTxpU/oehgHhrqvhA2nMDaTbCXBzAH2RaqJnLSUndV0gUJ6R
Ld/cK7NZ+rnG4ce0+SGjlvTSfJdIr5v3M/BFlLQbecvVWnx5Gu/lDzV0IBaTKjM+
Os9Ild+QiKtJ2YlzpMUdqFR1dp0iEobb6Cnmi/LEicaISQXm5PVdhrapG/yB8ibc
hTHBempdo3frn0F90kbav/PmfTOQo7r6DzAjwWn1ehKrlRt729wk6A5jO4bm4OVJ
nqZybOuy81sKpjfvqqB/RsohplElX2M5jjfY8r27ccgLjhDIAX/lSUi3OCNQU8uU
KRGI81Cf81Jb9sgKNxDhZ4F4ffyGj6/oJlmkqp6HZJk3S3B8s4PclURy6Y0jAtaD
PfzCIdeYmNCByZtLMFwL7szqyMLj23kPAemR0R1a5AEF3TcMmSZazpCJbXBTg4Gn
Gfn2Ds7GU4xb4B/QeFuWcVTBdHDsaYqh1ZOWAa8X/pagVW5fNjfocYxhBs9Bq1yo
G5IrVxzJnzO8bbVm4IX5K/5HvrwTvXCi+DGg97Lp8b/rc+GpWzjKwrBDp6wVWfOX
uqeN4A0fjaKauHV8gJ3NpRcwwuvo6S8XzB4mQoomP1xQ2nHOPToQk8HafAY2FG8n
f9xGjjoRiykfhD4qDBhAA5fSNlKwIiVhRURQTbLhtXID+NQVgIXE1kElPDFjD26E
YoDYeOIG1HdQB2jgH6Z36pJMhL9gMW1y6jJ7VnpgdeM57rqPSPpiE4+9C3QqT3Vu
p4Kqf7QmFw+eml7U7V8wRacejj+Du1PJi4jto6n9AaZ1xbjDm3ie0rPBdYutyYof
9KaQTe7I7DAYdO1lkW8fWDkRLvMvGz6lx8Kfy44knpxdWy6lXUP1MPMBErykW0rU
6x6iL2Z8g/BEMDMYWDP8gbIMTIWXmLU3/XqyyPTWopYujpfTPflSDxewGAIPCDVh
zH1gi2TRm7g45v2+nPMr9wirO6Js0540WzC8EL7rNaIZ1DhGEQAsJHQFUeLuWxGJ
bYygmrVG39Xs//jLWIBiZqn4r5951Ovf/r1+9PXbMK/p+1m4ymWW1nUrt5UTtRv6
oOm4DxtPzrAVk2v2IqnxC/3k4eplDD9khkNbEPZRDAoaWLPEzGFpbAovYuKsBvAx
u3eFtl0Rn6lZdXqdFA5nleACC6+c/G60SfDDf+By6NmBT9biZyGegKxDWSISDGNI
99L34LaJ1lqIXdpFtwNR81VCCk5BYd4zFfiO15Zk9kx+D0DA7Yi+quMjPYNd+sA8
ZsaoDdXmnCGHfDaCaS+D3ijncK8caUbegyKL6i0EADHE3dLHKxb7LB+gODQmx4z0
tVcQDCS2ozotXL14tQxKp+lQUhmmu6eesOkdX2e/p12CSWfhf+SNfmCN1Yj6Bzyp
HrPxHIlji9zwJvHlxHQasMZMigC1mcmv1HAHlPekR4ACKdVoTtNgWRyGZM8ZeLb/
PpMc8M+dhaH7o0zlssZmDZwkrirOctv1XNM1c7FX/YX12wnDgIyhe2jVrtkhQ9la
7vIMggVrLbMVwmx3osluU9Gtpbwzh3F4WyzRLOt/lRSqoKy3wDrns+CK8iayHRvq
3tFkQkhdU5jWk8HipnoJgNwwYv9UyIxA82eseuTsqknLekpgggMCB7PZMx93S8nk
2DChiQHlU25OAVLzSKfqs+W4VtQLwMi5HWRYI9Y/yuASg+m/rS658sxJ9qTF5Xay
tSZTMXqQ40JqCSshaMVjWKaRaG2qSFGqS5qveZy0ezDbZKHYEOAND0qBY2EtySb9
QylaCRl/VPME6q36KgbR9WQrFpO9iCwWEehGHRxKjr2cZHJxyuqHlLg318dL2TP/
cAc+XzBCh+A6ODs5f1/T3zuXygjGlAHhv0535lWtCl1UeZlQ0fQFy6tiHho8UygJ
mCyGmXvmGSod9arrQlsZTqFY3fC3LxBdKtO81jJirLJCC/kWg22qYwUQibnaSOY4
RnwF0mSGEr2UHlboJteOynridVerTRnb95OC5UI7OhvriBBrhfnSc0J0Ra9zrjBJ
FIdoqbpvueBev+uFsA+Jdmw8syvANyWYPOPZ2hmWkWMHFQq8CK/KA38imHiTepXk
4DjOp5NSsEfiWkssQL15n8iu+4pZN6JkxkUYoUxOftQiQTSFvmA5+yBFKjwY5815
xcJJRuxh1V9T9JQjdfMKcYbfh5qC2J+C0g3DemvEnhDlEkvuO87jWiYQw+DEjYST
Mtcr8ygOZme/Mv0TKmdn7Jn9d89kj5zRkmJ2134Qy7Qkh/42atUDHKtJiU3nD1l8
IaZOYP8mmlOph58vTdwOk44gwtVhiFcsu6d4GjbuitEc29Bu+1T2a/NY+5NQaCiF
Yn5gnNcQblOewyaJvCnxdkePvcHOiZqb0S2XqkMYFDhIyHhK3N0pwqnTUOM0TmHO
eGaAArNY2CWOzX/GmKZyCiJXgdjmc6GYW/qJ1cMJsrzATcRCiMd9oDOvsXpJmmr9
uQRabtQWd4e2sQjXiqr0UdJfeb7aGFUvq4XpkZ2UcTZuYamqwrxYsGtN2RKF0Zet
kDCE8/KlxrK/JfLJXM/D7AwwT3EF2LUWYttioy4C8ui2+rX3fij3dQl0xBP9tqnU
4wZ4gBJOf8/rc0G93cjldH07L1nHSz6m5MjkjUcN2uWXfa94TmDP9SjdpkTzAGxt
HGYyIvU039D27xvtpqsiKP8h5poM9HBldC4oP/bHFXgulQHL7ePqcBVYWyNkjwRN
MTdp+ciQHxsfw+xYgviq3L9uacrhrnhd/DhsfFyC37f4AKhcacN3Ja/zN2SXk6xm
LPnfYbxisbLEpKGLo7YPVsAhRR/85Cw3R81+mQpLUHwlgZP2WdQshduHykZVke+7
1i9LaB3d1Rrof4m6MbnTg9SxYTasQYYzkagX3pM7ybUq2qACAsQHgbb3nqmgybnn
Nh+Kgk+PXUXhBKaE/N/BZWWYZxFeYduff9PmApYlSI5g5eynPDUUQRuXDHJNQqTP
G0jl+Lo6PTkHmwL9mYksjmv5pyyfbgEwFgqd5cx2qCRr287tF+XBNxP+BGpXFxHe
Sj1NWNVLmGWNdkhK7AQzVRlZn0SFACiBQnAx7JI9FrZaMfgUB3OkeNB24m0v1BGt
P5bQSCUw/tVrVdukl9XuKVUR7pvz5QQSbOyojADzdWuV1vVrpixVev5fnUoGs7bM
N9HU4Bf8vR4oAeKcInUWzdRCcsl4fnOeDX2z5IAOBQwYmlaYDjLvurEhwPve9wiM
XhSQmXjKh4BuB0HVnS48DgnFvt0oEQKq+WaOlMYh8j9rDPzgqHc5ajiOfmMLpbjA
rcGmoWmUNMI1czck64c2F8NeIfNhR4Aq7O5Jctr+I6RKRCYJKAaCvC9FXmgqQP4I
C9yrAdImLEvoL/7y+TxFYQHM2E2CxKi89216QO61osiHU5KKVOikVCRnMOQoesIV
16bXK+tj6NzRC6HnU41k3g8DMM5kYGPD+TXPCRq31fkPO33HI64CaVVBKMgIwEZw
NXF5h1mnfSdlR5iyBPYBuNr9GEg+3ijHy9VV+Z5YEtO9dgrV+km0RRzFQQPRMLTZ
znQ5f3ZsahpGwDcPIkQUVw/XNPngTmntSffsuk2mszz61rQmR3uqGHybbIq9AlbZ
6OZ4jh4jCkpINXbcx6hf4gl2OtlgUyeUrb1caIaZHlFh23RQrsQ9HNwEmxlpCmkW
Pxoa1MIEm3HHiZf8jjgKZgiN3fxBXymoAde2cSMh1dFJ8bghsMgGMUK547JQ6cB8
RN5c24Ixa0Yz5CntcmntpXlyOcVP0YzEt24ppKuv1Y2kT5y6nc0WfuiZVmpod+LQ
H+VqadV1nLx88vOnsWUR9Drq+HJd0keH85P1A6pZ6zDY5tnpDxmUoVS93DHecMbK
Or8HbEPnQkVraWIUzK56atnv4ssM/B+oNdAuU6Uz8DqgzImZZvlKqYu8hZycS1ta
XxOxePO5RxSa64i96H15sRpY4QF5e9nOe/05RR26RCZ6p171om4mSKeqgi5TPSRC
FONf1K/8sXkY450ysiOQT5YC3kP+dA9iU4TYoy7NATz9QXhOxsKLEv3LVU0KSVL9
OW9/Dr+ziZT6aIx3fpD9bTmj7II+DQODcsq1V6qH2awykJ8PBV9fT761wN3iyqfc
cvoeJIJ37UKk9c383kaup7aR2O5auoIyS8Oj0Y1Kk+1pbjeC2204i3xzp8qHN9km
X7TETNAeRP7OZWgFX8ApQt0vndE1HlXSjMF6TR0JKjX9jNvG6zBHQ2W+RC8QQ8bE
4uUKO2Jbi5hSdZ/dd2mYcur01Yd3vyrk2ckA+Zh6gfzN3OeZju3gy/o+4JM/fMF6
ScM3mMASBz7HGK5GHVgSplrJiUh0nSVOJuRuLILUQWibUYNCNbITfuHRo7MCe+2t
tm+Uqr7+eUSIN/6LDoLaPT5idrmxMGywD8uMEYbQ/fjh9WwUTcsZxP+6lBIqCPco
794M/ZLyi92qdSYKcQ5U+bjDMSJr4yXVz/+tRz3gTOsRtwAmObuzzu0SLIYG2ONI
QwBNNUv/PH+jvMWMOPQOPFJ48mmGnsG25NQcalcwLh0w/ebtBQFyQ7AgOgYNNhqT
rgzHsxOsKP7tBfBs4gZ9ZWStnFml13/4t9W6CSdds9cCm62R+8h5uHpiApyxU8hs
rhAmHO9X+P/8jblTpwDOQB2xrUWuX78n/Zfvg56/1jIZbvjuhscbCFAx855jdW98
/D+SjJUL5Iws5TgkABhvSrxDiKhxYy6mQ/1quBG0oGy1Q6KdXUu1Z4A2IZiwRiOo
s7uqAQqiKkQSyaALDejryBZcLQSBSwrjLnNDTbfT0CQ0/EWBQlioJg2x+lKkslI8
S4bkosgX7cnfyS+4kG7/oAVWVJEQiZstfSX35O0zzCSsnIWwdAisNRWUxroB192Y
+MseCntD3mkQcFxn9AWLfgd8Lrx8p6qsJeOa0hjJ50+GsSNrkfm3tk6BdMuGcwzK
o6i7BjCbdbhBFZ4iOWKnI2D0p7dpVM0mTrvh9iazFdwsmbQGTNgoWKZcnL5SpcUo
aZvpsaViE82TQ9J1d4X2iNJNmOMn2JdyotWSjFfg8Tt/oa+xfOlYxMDZ2/mYbGmL
ggCFDor1PlCIIxnJgVsOqOSx1PaqFZI79hCGNGOX0egD0aWC2RZBJGhHtGztUSAZ
xRpg3w6GbljZHaNqf9sN6OVSx5q2f+ZcPshEwAxKOvjgoPEbExB40xgETvHBTsOW
xutmnxCCkZKo9eG2A4GvskswiTFU0ySRr359Qb4DKhWZvCMuc1V+N+LI3w+hEonp
bz2kYgtJ+mjHtN4BJmEgmEdimQApFy4xcZLWp6TQb6pI3Ng3PKiI3uFr8wpHTxgy
4YQ6cJR+Wmckh8S+kirJRmsXhaOMTj5qC6qTLMnp8zQ6b0rQ17WjNnlHzByZ6ePJ
D8V958VzfVNQml8cQoQ2G1eWhJtduz3WNLe8uxUv2Fu9RJ2RVeZ+TDaxX0EWkDEI
jjObBwPexo7CpH7G/zM5SwTs8ZnCAC6/rwFu8PoKQLUaxwxNiHfS7stfGdp/TOPT
Ve9JZrULWtdWgyphLFGMfvLMnJ2vWkGnM68jc3c31yZQiMf4EA3h5khDf81lRYTk
pk0t1L/xkwQ/IWNjUOxh2x2loR7QCZxh/6FExhn7EeAE0YlnrpagJxKKwRvI2RGM
2C1NIOKKm5q9rY2ZXIOuk8cjZKqvEYLaJOHE32xcCsEFqbmA7XuL/Ahq8ZIhKfGy
lsv2889MB9FAijBfrI/RFY1ZKdpbSjus83fO06eiy/VJ8ENYokJQlm6epTHUQLg9
ANX8tQQFMNO8nC41ZdUsamLsRE4bMKukSJ50kwasTF39+wQPM+vubNwgshP5FATn
l2ZXluBm970m67ZeH0aS7i+Ue2DgQhknGz8DmZMNZQu7/4RTO5frQGRJXaOlA+rB
OOo5ufeLi7r2OSOJM///+raSQ5SLDfczrJJecfGBc/T2IwX3sp85x2QjjX1lAwMd
gI7DkSp6j+UME39+F3OxycQOKM4oRLUKIahOFcqMnys+8TLecjj4v72/DsU+s3Nc
eKylJH6dv1FKjoQnYw93C8Sy3sXt8d/h2PpTUGkeJHZfmCwHaDl0TQyWP5hum5aN
kiD7wjL2KdRP6XK3KbRlZNVC7Td1+qT0qlux6KPAiz6Nd2Oi2KTWW68FXMt/1aDp
cj4sX3xJUg5KpBs+chDPz2Rmy/nKW0wb/qrMwhFi/ztr5uM+cdnXb1C/xOfQ9q5G
PL6CMqSPcB33sH3WvT4aPFt01OQ4pVhs/oO+ghh41VOCiamsBy0Kibuk6m2Gd0zG
2kCxIIIC1seJj/V9zh6SgeXSm/CPh7fT/5ZROjERr2+QUow5R3U3wdr8yj9M/rtS
PZCM07A+eX1573WdP48WAziAVgBgpctRkgAxXSai1jNN62jnjMofcxlbgtabdRGu
ewzhb4SrpKqTsk30QC4bSk5VREMN+JSwUfJX8a7Ke21Ab5kg85/eU5dMtSDrboR1
BX4i7+y0SsDA2a1PAeWn5qmQZxI4uFFfkSYreZ65Qw0NFYDVLrWLmjskpaN6PBmR
JFB5wChUPRCOIoWqEGOvC6cMKCBSWbbAkzJW/+DhU2/pHN3Sv3kjj7mlL2PAUgpU
hrAsaq5tAsLQvyq7keUnfvilKyxxvOyVIx2ZXWQUAX0dMPlnDd7BbL2QThtGqoFL
xK30hrjQdNmikereFdaEqtf2t+GHx3IzvnqKro7d1U9hUiQwy8a+2IRqkj0eBLFo
Rk30827GJi3XX1yOSg7GmgiVc7cURPrsp2lpg8hI666Zl6FzLrzJdJ7osjTaNyAn
IwKLZYA8uEgiEMcxziubxYz9ouF1e9FO5vXXgnmwLCwI8Wg2mlfJ48oMaucUeHE7
`protect END_PROTECTED
