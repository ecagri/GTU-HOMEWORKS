`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YMMW+c+wehkCiX2t7TcJ16D+5meErbgZHwhZw05dZEivSFA3/W85+Rgf7Ztg9Xim
m+MD+/tQmpaWfNhE+ckp1qjP9weBYAItqQ6vv5mvBGtxmGl48ker3k1knakFoCJ2
339Y3Mese5HkB4yUEJoVgnqHgzF01ws0JefpNnj5bMK1JSMbpAkdyKi7kmt+mfan
vyrFntwvIGjTQjdl69t04UBEx6kN+dmtqNrWCuaNh7PWvM7K3kwJBT388DGUFD5+
KPtAlOxIZDJCvR1+4a9R03dqL3Sjch/G/Qc9Cuq3YI0chCzjf/2B1qakjKB+5UcO
uuoRz8xJKqR3v0V1OLhKj6YmAG8uiuxj8zbIc2ON5Q+qvgptkTURR4XSx3qTJXVJ
`protect END_PROTECTED
