`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tCLiZNMQyuojmmq6NkIl/9hkfFKQIet7HjoC8BkGaNXrDuqxnWiXUDEg+j9RyICK
+uG2uLHYvcRKpMLccORhbjZlW3ALh10xokfFQhp3Wg/UGXsyjeDcX9uFBHWYCSjb
9/6m6jp3yJaY0HBr6gur/sGSQDqr79i3CeC/qwyrOjU/PhQrsHJXqS1RfQiZ6ZW7
C4FOJp+CZJ8+ir/sv2mAluja2iw11oeZOR/cT6JXX2b2YpVSBviRwdlRUrtjOmsW
VRYolNKjUXYNt+ngS8KfcPsMBPYTU4lGmS1w0qbHStHuCSAKvMaB0nbOx+XgXHwG
296d8IJzmxPNjdhzbAd8LqgR2Kv3nn9k5rYY0+FlPZ2F/xPcRoQaGi8p+jfm3kW9
KN4GgomfZmkGmfFJTdR2OGzNTfQcgiThR4RKIHRHOxGrBgSU6ge/vVqMFHT0b6f7
WN+xqkHG0A0c4Q0d1c3RgDwfiM9SidqJfqriuoVN8TyH8uEDrPzmRnRCH09v/fAt
wqqt4GTiVk0mQPXXOOlMKIUJIx6u+Sn7JdjZsXYDDffZHOwJxethd4Kf/8T0ht60
+umyc7EP2jTbkUD+nQv8JkfsIgBurQQxc7EetaUU64ma6Icf7vzTLmJ9aevj+fro
xx1M4aRiiDqniMlSm49zQ9uaATQto0I46ZeaWe+J0MFr/Qdz1M7i/05aqrVq/3zf
TuN2g7D0SMT4ri61hEFeBSV6ZkqO6HAzch3qK1kGnlF50LShbQMHT40djQEKgQ1o
NJSbZl4CjLSyPgA0MxwRq9sU7aCULhHY4uHLyw2I7lw=
`protect END_PROTECTED
