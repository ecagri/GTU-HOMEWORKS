`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ab3rtlQrDHipxx97WPp+7kiN2Yb81BwnDPpg1ibfWlECR5PZgXWR+NbVARKXKwGP
MKG66W1B3UsyEKTyQP+PzyGHQegGuwxx6+mGIDVCw7tmx6OmD71hLpX3r2WhfxMW
o9scMc0qlw2CcON3thaqLNGSn9uDxVIPcM8EXps1an0/GdXvlgbv9ylqNQcZfhuM
n1tX2WRGpxN+KKB7asetZHwp4roXqYwfKfWDJIO8kR2+RUPKG+tqf8jEbEh1Fc54
n3FJLi2aeYZ42yhWIpcjxizzOXhEKUG/CeSQe2SYHlyhKhyAy3hqI2x3pqlLWpBW
b1xzh8aa0p/x4EEAUf7XmwZxQB8s67L72TJ/Ram4Dv30gNeVaCtlsikeMFAVN0i2
SCgaf/28ZKrDNRQLUARG7YPwDEEgDcyjcQ4/sp5KLNZSiuT8BK4FrC9wQxefjhm7
jD1IPV6IeLqNF2d3UeTjM6RBtPZRRBOkzPT2dszXu2fADBZBvXkqf2oE2WnkOM5I
fyKthLxe/XQ3QVPU3jE1lh7PaG4jjTcc6YmUK3Cyx4y4WGcQRf/mztDtg+WEWK01
oXlI123S7nbgATmxQ6a6dMxPm4zkZn2Et4UsSW4Ze+pP5sY+PSkKUeJttwJ52O/i
MmZy2WInAdli5p7uV8rAAOOi56K0/hmaBp/VeFiM+wA=
`protect END_PROTECTED
