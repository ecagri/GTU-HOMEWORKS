`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jk8R8+u30RnY7y8q2v4z0vHWs0D6L8xyiKJcdBBcaJ+u4OnOFGVKrTltp/bo1Q8d
l1LSnxdigRoF+u4jwzeghVzfcm3hRh1AtvcnI/3DjdkrMWjH0/FOggugzs0CJeLt
Oxi2pHnb5B3X6skO/bOyFyvSYHxEU2n86czvi3ZNUUwSczMnKW8L5iZcG7Z3Cumv
U56aTITUAOWdR5JdNRRW9O1vK9JknF31Pi0svVYFujeOiMMvPfOqbVayhvfh7lwS
IKfKIcI5YZySnyijrgZjpORr/sr/1BIykNy/+OWEwl+LcoaUwb/DRLAFUXac4/Lq
AWbt32lmQqWblyu0lNdYpXf7UakxvITjSI8iWwgWoEg5rqXDj3P5Spio52ieJaP4
hsvG8dXrEx2mefgp2GyuF9R81fUv0pMApQkZsPT+LHA/OdkwNJwSs9jYkKb5/vYQ
+/P41/p6xRQaTQBcWoAjH2XJl7p6oSFtokdvAupUNnP+qCQL81Z8niYCCVhaeEzc
glGbtdKakj1hmsdbAUHPurrr+m6Zh5EwEAv85rdD9l6E7VNeZ/BTeF4H1nHi32zo
KelfgOsNdXH521kREWbalGye0jlLGB3iKAu26pdo0YVBkGvM9/Mwc1kPqgmCtukR
ZoenRf9URyX7Emoh2oW6oLj8DBoP57sfC4aQwePPx/OmkgaABZCfgw3Y6PMbjrm2
2O8mtR8p05oyAJF2FXmNR1GksRvSP/ipmXHsbsaaltOwKlI1z9eKUtLBL9yKCcIr
qRLxGP/9mXNzw2nt0ZhCY2w4bsOJcUqXsInmg92EY6wcKgXd3JWmZ05sRsWLprVr
sCPJG+seDWLOLBWAL3E3gu2HFov8ydX/B+H/az74Nhg45DSgwC6juXrVBQg9Piet
17axb4btOcrfHhRenpOavOBf1VtFq/vr9e2+bJmm1373hc9kF6W+czMfGxg1+1BJ
0OsrPVWOpaLRu5EAYegvmx8TnSb0hafVhYTsq3bou5if20spYBsKBt6B6WWOUQG0
JZ2n/R3K2iPyqTLhN9yX9cArtl/IUCQAwk4AkL3beG6WbReUw8pw6C3AAYTtd5+6
`protect END_PROTECTED
