`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iglGF8Q9L54yXRsLNLt0IfBHdnlKH7t8N1Yi3qTHB2KmegSxXFukxgIRo3AF8N3a
9F4bce4t2bR2BoqRI+LAp5/ry4Sw2FF58C/keQlpNXr0D5mFvYspeeCRgv/ip6YD
yAdqRb2GgUbfeDE644GOF4FvYoDFCyYGEy1j2tPtdGW/ZYe/lPWenv59eAhfp7dt
cJvmBEW0xfCBIFRhCyugPFKuN13n0LieMsKRHP8UXahzEJ/ylbnfsQVm2mE/VxvY
VCWSUUxW3b0p1VKjKVssihqXH5RrBimbxVu1pYv9Q83HC8LMkrfVCcPxu8eDGJk9
tS2+aNwsn3jQ8VvC8tMhMZcNyg8f7min4FrJ0JgWxCPbELVYGP8cAiEG/Xem4Y2x
13WrPtAD6T136+uX1vBtXlKm5+pDyQY4+5K1JKsaq7IW1QMqrQkEDWD3Ft1AeiFe
+YwF1/TKkeaeUrhpOay0dS6i61I587oG/5EnxdSQGDi+86lbIpyX7AhIKIj4sqEl
DpHLvmBR8lqQtAAyGRTGLa5yluswgoq8Q3KVjFT1G0DX+lTjj80jkLZPoiC6rxYA
voB5HZ0GsP4yfHk/rPDa5DUpjwcA8ut07EkI64T7M6AwBtr7/zaMuNBeQtzTCQvq
uyTzctkfsSBjDS2g+gEkojCrQnF26J50CPPMkdTST+FGsDDkJt7jwBBU5p8VMf89
YmIp4KSBjUZbc3GG+t/YUjdCjC41VBwQGzXFc8hBFIPpRpE3EaeHOZ06aHWaqKeA
6KnMJOI9qXGVbUVnwMl8ffFHoZbSgC83fLPfbEg+i0MaWndoBatdqU0tq/ShiCRH
ZzUUPhgzJqjJwZtM9tEC44aTbqR2QokJVN8IL8XIxAMzomb8JkAfUNEULHpG8RU4
0xxS6f2Kmqxc+FTaas6vfi2NEAJ5nFXhDKhS4NXdRDyT4i9ck3ufj7GXl46y+KmL
GTmPwbJfnjI9dm0Waey6f1wc07qm8J5KfhisO6syaLCbvKGkHuAuDLv0IsgDE9zo
WMYaZfzp4QyvDXu70Wn4YWJX5oNI5jYn7C7+qJRh7IK21Pg4MOYJkM9ixqGxiPnB
TTPgu5RkEmaVkQlx1pstPMKl7cmrINrzFO3EqzSVR/kIdLLoXKsZyJBHEa79oOk8
FGcG2bEKSkgUjBqFjnhyYlz3yDXOIaC/ni95wqV5eSZe1bpuuauERVFv7u7N0/rA
N31TdPLFXkBlBQxxuJl/jUGH+uP+B4f+9Udq3IbY9xACwG/D2/8ZxSK/JzgUWeVP
wTQDoQKRM+BVBIIkaWAouak4swoygU/roHT/hL/eFpN48h3E0pNwjtUiTOjpVuSU
XVXIoMC62cx9WlMx8mSswdvuJ2M41TL4+Ugsz/D3fB+gSICUleVp79WWtobh/uic
HPYPngQleXK/qLugjQ1yW/+FfYH0rEdXMoHZGmnpfIdmxy2z4K5kSQBAE7h+f2Nl
Pdj8Ln++UWUTtWJ9ci1Ua13Y0idxviHaFlTbtGEyDfVUayB3b/XT3DXEUaFO7VzH
DvjgqP5WoAT1BkeYHgO1VETk1VE9FFrfpPmv492F61pH8ggMZYZFqoFeg8IP5KtI
OyMd5Y1Y0Lq7BG5N/WrqA9cxLzdQOAoxU83kjuvsjslxJ+bYk2OZa253uSMsKhUs
UcZ1p2MCOZSiKQxH7u+GWbI/abqeEjo42bO0vR6mgizGCIgMwEgTPgSmmE0E+An4
tpNw4FYXAyld6Zz+Mcd6GDA0W72vtztg+aQA7ORC/zaNaA6673QPatb0ulu6mUBp
5xF6Jnm6MlgS167KeKPSuN99unx7NFzYyjN9sTzHKHWiUengu5U3Ee7E37y3ld+d
KtuINe0VT7mOgK3GS4/MPA6g6HOpvF0CBLCwW6ok3n4VrS+iGQLG0QjumB+JWhN3
p/s5IB+8h9GZbenoVjMk/jGNP9Rk0BZ51m0XCJeqQ6YwP5gQXkLwqkZ4NLa5mgF7
TkEZY99PSLO7fglpY5seUz90/JgkAFSuwJEQO4joJK6nAT0gSsnYUhfl44/rZsMx
ft5dpB9O7g0voIAsO+o9dU3VVUHA+bce0bStz1G1Ya+gH7TA7+8+5qS+SgsK/HVT
WClKmyH/2nG4laFif6Tgr771uNr3tQmrPJts1HfooXqLBrlFx5RmKGESxpsfHYDG
4MGC32iJR4O8cwPf+oBwd2/EZ5QAagyI2zP8xpF1Mxq+hanbZcs31hTum0JEec8/
/sXTYQ6QadqrWrcVg9jMTMVXjvjiLeJ7dX/GU8mN4PK7oIFINv5a4BTAjI3gObOq
uYXLYwtj7S+MmqEm6y+zv/sqGtj2upAvENsgo7O/KpQuApLEMHLLdNLAnlDvIqEV
c6ffhhXv7oBCfFclGgVI2ZmFgBNo6kG8ltkV+5lIwOlGWGdTKaOCxC92EJpOxm1+
6Z64jkKnpDXA+RsUzXlqzGOlh0jupM93XbDRuI+u1qiRL6g8DQCZ/LJX7GybT4Zq
RIuCuNVwnnk72hAjzqHNajHttokDWXE2781pojCZeyBldgXq3zODFRYKYXhOnKoN
UklLwyZjF7PigHnhbMSIrqXqa01TivJr40ZracId4A8h67vAD24DfUVQn8nFiMtm
eataenFLGEw+8EWMsTEig8XhSDbef8FHRs+um5bNd10g+BKjb9oIF1mdi63alTCm
9YsoITbGibuoYobDxytxYecnKnIho07q4LkQud98r6MgObbpM9bceguJR1cuShsI
6BX7H3utnRElf5yeyarNWW2HF9qqRtFy32u2fBTLK+eI47m+eXUa3atcaBievqph
XKC4pBszg0vpr/XBlUhSfS6SVKRO4UrIya2s8TG6eTvQ9BxboS7hzr6I60pjU0km
oZU9/YuWxzGFcyP4KtVRIXNsiqC1OWQ3dZzu5flE0xnLfgu6Tb2FB/KTg5Yl2eAJ
HmNbULAQyEFdcBtrqaMgU/zmyBFjz13W8Y/mKJVAQMUZAONLrhdcrACEWfVo9Tla
+1PLagmpnvSa4ZG12YLcwlNInOTuinBk0RXJYVmlOlTSbguJzjkGZyEaF9Ux0YDe
46XuirEFiwnoqU0NFxy5GSoLUpREOb/PUkPModKNyHabqsIvjaH+Qv/p9pxoO4p9
GUH7STvGb1yBvOItAJSaWgf7FM1Dhz/NPITC7Udj9J4KQtAxxkJ6EihSEUwW7tWE
yqQ2O08eqQi+aE4IQDtlje/wy+q9l8A0cOIOWey5OLbnZrVBq/d4XpzCL+1ETeb3
JDtIv9bW896woBBak4rypYs0YkMpFgwYSxjKrHx5B5z+pt90NPYbb1LJolVwKLOH
VC5MjOutH8eBn8Qwof70DncBRI2vi093sTtJpF3ax0MV2qdiLchqUd1l9LtlYe2n
IUd4oTAZH3pK6/fFR+TpSA02bnmyBx3SRnSb5Gs57dEcfiWH3Htu9LbNWXJdMnY5
MYeQXq7A2/k/j2SC8n5IrSx/pDrhNUd3iCPw4hwDOfJByiW/kH+B4ZLjO2hnf/vi
h4BPvPoGquZkm3+u8BrGWDvXY0SiDDZUfh7VOXVfTKqQMeOP8h/OTPngeLXzVXa9
7k6opJXxDfnBOJ3D4NU8NlubEJNSUFimdnINHeX5cuDFt8CMZ78Sy8eeg8fdxeV4
Uru3iQ7CryYrvbKjcYzEhfttqa/pZZYrTQoCAQNRUtNHtIig5nYN8nVh7bM5c1Pn
VpR4bPJca3W/ElonIJ20IJz1a7wlieQP3qrC+I5q3C3S+QROJFP8pPIwlG495/Ua
fFlRIy65frQ8EPVi2epf+kB73C537QwLobngR4eH1I0KYut2acR50pg4QhNSRVkG
UZTchvp9flKaCsZiBMhKfnfcWt1r6UNxPfGtNwAGE77/rZHxkD9P/DmNDNO1p3Hl
iYSiIH64qBeTqqUJ59NfcYeWPWYHIthXELygoheaf/9T5OBiVxy059XBrXJlt5Ib
HBV2vAEmVdyvCuXpC/yQosP9FYH4CKvuT+CCyVTEIibyd4cZciZ7kG/6CtZutoqv
4+EV+SMZes79PCDWV64NBaZ+dPiUaexLWgmxqPrHUuX8mvxnY0JGv1BuEpHHpQg+
55RB2+dV4BTl/ZnqFNc9lXIMJYbJ6+F/SPXuxJ8DdxRC0NKoUDlyMdSFk/1jyso7
Xk7HZVOpMeaaH/N5TAGsKqgXGWvLo/RsxeOCeHFrdHVRV/9B3m+ZwB/NntRsnfD5
mOVsQd1j1VUz37hYwhQvUOEdfWW5mq6NLlPV0mZcOGUM1/w2oeCWfFsF27rXpfAi
BX6UKZNxxt1U3WpeBs38qgulIY2AaoDSgRGts9FzUb5OJGiUEUOh1/qEE+dOmbYA
fJ6TAaiCjdE1CU2I9PT8Bu7S9W7Ye/Ykn1Lt+ambQu54ren2TLfFFAlY2LjUZuUD
BgrNH3g1YN0syCfezu66abJsiZgiQIb/cm6ama5NmKv4F5sFm2UGdRIA1vJG+EG9
HZHi9SkxRHHwKzP4+KrrACGrF5zM8U9THfCei6kuYblW19MqVNfOGshHokRo4lZs
hUl9gADQ5bj3mq2caqPgjhbzgRbR2IYZ0LHmqIaIFm7j9OaQACDKYXwmlFurANVc
BJEXA8uUM3Uk6GLl7JEvLKWwz+fu0KztlhV8LKl2S6v8bQCOJT2wrf57ax1cbJQG
HYboQQ4C2jVwz1fXlUfsujPtDYfdc/4SH5Pj7M77D7br6l4G0QMWEPCg+cCLrUzZ
gfo1RG1kQ/sTCS1W2I9v1GCWWSv0W3JX4V951JhwtsoagHTdE/g57Ytz5aappoW/
YWuczpLap95+g78SBSHSmgHhm0MKcqxs4V3kZ2861MXi2+pjtBundkHNvLMDiUyc
Ohhha7NG8on9PLk48yd+7fz8Fe19ZMW3e1ydhjHiDOjZEVmDFn1nvvLJeL0wKYbr
DlaNEL+ma3NxEEmhk6efs68rR0PXS9nlMzTa0N0bsvXqggwxWymEXIxQQFXmaZB6
u+m9JGo+rAU+YH9DSlilGfZPHlU6EggH0IeaLVFuUqOgckP2jeLYIGl9J7A2qwXy
wLwS82dp0heVmdJWiTr5S+Rs1PbUH13iHjEYzOgfIa8ly+XO0UZtVSv9KBYrIW49
kSbyX24hW3iSjxaIomHlbE5w27OUFCk7MtgRlq3+NhsjGN41fJwdXe25OrTUyEwo
2RlPngUpcLATFo9xIoqT8c0nNjWh2cXZVzMImjkI1zXy0/XJYeqUzmT0ExwzQsY2
I7eLbQBPTKz8ufiykWlE1nYEaq/Hac9LEyYIgFuyMLuaGaGLfmeV+qe9sO26cgR5
cRmjNw14lcB5PMOZt0WjQ316zwdBWWTtbzPCehjQ01BtAIwC2Oe/+u7K1dwEefhE
87IlvZ1NEqQIeN5pYtt5sswLB37dh5oAm1NzvmgUvfgI2UH0ogCUznT2IxxLrRg4
q7/wVrmF5/E/GUOCac06b7gQZkDLSXF7p7sFhpH3W3/l8P0BOEkKbwcrb2CJGpqh
rcM0WeHhYFhUDxAfNDymJ4ouzwgpObBaEH1cRcyKWnzxzb9zGkHpNMze2mGVr7pT
nxvw+TXVww1DZKV0YcQHf2L8ZwwT8nfOlZjEPIHnY5RnbbVMLlTBS6KAV2olCGFi
6CyG5ixQP3xudYFgGwQXRvfI3q9grl58JuPjrbyQMyIApKf0u/KX9VcG5bxdso0U
z6/U/+n6feyAFPI7QkIFZMgiFoGw50I0p4qQmtc6CUYvv183+H2hpid5RWq4za+g
9MIKndbD0oAmJ2K4KjZAwjMlJiLKmkozkC1efkpBTwetVpESQltbxEvrRBBicRrI
DXKAxFa+roJeI5yRqBecarH7qnkrsbFzuWjkXn+4AChe8UwdALpvFTSGcFqCpRMY
n7lHEja1bs0RguVoPfXumJK4On6T+Q9Amseczglhr+hsb0aotOoFRZWX4Gvx8WZz
iXmASbVMZsArtC7BICIQzC7wV/2F/lkg9zgRaVvfFj8lztBBUnn4Y/1Tbf4Ya5rX
1mM0YySSgFbKUBIJV+a3XBzJnZhCQgPRiqyq/h4tzuUQ7epqjjQfXqiS8X0W+fiC
LKiOpeDQTV37UMAzpyga0Iiuu3Pg1G1is8HnNy311TgWDnHaGMOtPCbvaWLXflkt
FGET9KYTJtrT/UYeRDh9fkcXg3669+I3/ajOasE1Tyr0k4S7c1D7RU8DwwrLJGIM
Ij5gpMUT8oVy1uFk1uh4Bmcu3y58gFQf5Qzl0pfvDd9cxwjTkX+DxRUAFX7GT9WR
LfHNFqfp+C+yo+X55+xrhb9WavX5myUvKwzltz3wBb23Vb2LP89nrI9AY0d7DoZX
pmuh2DIKsRL5HOiiqGty6Kw/QS+yeDWewfxz3CGBjugUJAcCn2/ubRA3yH3J8Zkz
okpb+ABIczKvDO0t8Pg+AHnvXtSplwi2TlOjDBctXvzGNF5rmZPtcyOV65FziaMd
nYDjVyOe8TyMGWCc4oDi/UG1McBThR5gkH7lrqkJr6/Dm67gPZNw9EnXnOyxsHPn
0k7nREerswRgxtnAj7AaS6kHraOkiJWsU585q3bDPrxK3X+PnY3l0qKWXzMm6D43
2T1TaL3EyiPhZyvaE9Y8VliHFipp7d80M1m5jad4JChz2tHzpPL81qnU2OQDdvUl
pV7LiTyf3Fz7ae2LmrDH2nIqrrkdMGkxlr1RJl/ODwkC9t8tlYI+UP1Xzf3a07QT
oWASlX0CJepA2blAbt15vT1zAoLf8RKVkz/k6rzMXE/Gqc5jesirk2Qv7F1dgjnJ
XhFigQAbD6CmM4g9/uspCIi8Vg7iwG8wnQEYKsyy0C2L0wM4p63Jwd3AX7LVTArz
wAZrflscvK5Br2qos8qTjKyvKpQX7bYQclk1vLjEnoul6Ghi3IrXKRczpdTh/vB3
WLVce/HiZxRaGoAhMA4XT2iJ6BaDAfBS7YYe+4m8ftadwo+k7QhPypKZD3p3V6DC
AoA9MBXbSsO7PgMcD90lJVli8QjsLM5SrIU9CIdMvvFw4CgAhV+Xa9GeDG57KOfj
/EU4aQi4fJmyiGs3e5BfdYADXxD7x4QC8hCo2yKWZnnS63jrtoTqCt2yMsNUcLsp
U7J1KjyAQHVYcubSxVpzbe8npjMv+ulUoJuoJ1PYR2JqadhOduedgLrb9oiUR1jQ
+B+ts1D5C6EsFkgLg97PRBTDQsEXonVImZiWBYlGwiVwFHggDbtG5LEU0fXFtMbo
GPht+HfNwpSkiDN0sfJ0EGtUqDUptB5k6INO86fP2vj4eH6qmNNWTAOfeSGA8fbG
mSfaX8jKNqX95VOJoMJ8UU8F9ginAIIGtITj186aU+X1fnAqyvutxsw7Bjus0Cuo
1ytunnptMhG5UMGuO5e5fuCbtCLTSANIMWl9rLQiQMZFtVAkEB7j3kA6EX6Mp0oW
nVGOVeTTdOCyK97LGWEYpP3B+9Sfu9zvbk/tThYUi33IPyz0A5sOigDv/4gIxnuX
upW6OM1Ys8D/RxtbkiQrbcAhilNWZ6Om/9e/cPgwjT3WcA/7ZYc0g7oAf/sS07EB
rjZ9JCySJz66ulwXcCtI9ZOMZ8qmUE0PolXch+19WhmSTPtV9k126w2KY45cypOI
NgUl3H1GSfBkbhNxItnCTQvy+teL3wjUdYs4EHYl8e2pkcqjX9Pq1fZ8D3PHigXT
QqMI25QLF9mE2QC6kA/SVufxF+KEtj1BRvn5qdxosWGLROqSMjyfTG46mWaCykp2
VWfh+ObOrdvBKtL3DMNJ3ylmUx3/kcKGD1R7BCgzyO1qBIe3symhKHbhILIWrswk
R93y1j1Pi8lopPyM8B7TYPIS4t8AC4AxFhgkEUdbD0dTrxzUnK69x54VQV4oU578
68LrkXNyLaGFE1pYUaY+NEQ4iwbXkY8H3O1y9Lf5o61oFNpdEdBmXwDeoMP/1DX8
2+zq3D2H7pIfJOZvHQsyZcZgLA83+DA7GACJncMS5DKZPNhae7xSLpGK8TqoDnjU
8pcXKnupgdnGDqPKeOTX9dBnf4uP/b3BSPu2cSuB52n4OkV4gH2cFQ8tWuNMssAY
TF/QlsBcc23nC2bXjyvkjJSgCsJx9uVf9pRSHVqLSkvScTmM4GtXlW5iqVS82N4J
`protect END_PROTECTED
