`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xz6oTh7bw/EHUFIWNVd7dWO6EjICLCT4giQBRnO8urwKa/c36e5gGR8m+sGJzeIf
SRxtY3rAHryVxsVIHPN/K8+sIZ5oeCPUQ0wNFca2H5d0/z9Beer1mL0nVU4iSgek
PwJStm3zp5ACszPJYH6pF31Kpf0Pw0WFv0TUeHCETEHHF6zA/x6rcnvbz3Fwjcu9
FZAZXQexFG8l93rK1FcU4yYHtWQWNiH0+DC6fyQlMbZREBFRNmx+NLo2hAXHYVud
ckGeVF2zPjKSBISFEpTNWh5qiejthK5gGbytnOLjvKqMh/RTr+xEDWz0vU4pDKyx
nwwl3pB+KeC49tOAyp29twTxlTDSbIS7ZYHdZmDQ8X/dxarj4tbWW7Ej8MuXWMC/
9XeqKhUpvv2tN2BiIvwxAjAdyqV0Psc2XaZeJ6MEUPAgGhEZt0LcBYjSxKZ7blSn
r7nxvrTEhLshZRDkSNJiqYOk5PMqAUKUOtKP/bTPxuAnpbivEM4boowarEeX7ixL
DElS+jyJpi8+c8xnsNB/0bBKffo7KhNm5xo2/oO24FjnZH49surhUIT6ZQSaX23W
OrKgNKn5rgw0LZa11wsQ5crAdUAxPeW57/Ol6VpeJ0HaAP/FyM2hlLEEAPB5N9ej
wkcOR1Bh68fdOP7gM+juqcbcPW5YcLBIdiBe3Sa552OwwbOfgcFH5GodfO8zA030
dZ7mucEoP+vrn/gGiCSznpMOlhVAcjvzLOcGCUnFmaD5r/G0w4vxOKkI4P3Cb4p/
iTjamWTtkKRW5m1hDR39JRpwMwxeCYEKKlysgvHzHaktWzkoJ7FKvuCEw6FE1+Zl
QeOYVE2SE8LRkJsct0nZ2FpPeXpa76cWyYtFnb39Bmo0WGRmMMEthTWNH2ExAGG1
cZ0QCJxxmAjPUxDKy9ReJDo3d8/D/Lgedrrpt2H30FT9xXJtRo6FBQhZCOSiG1Wr
O6ScAVCMtgZjibbTu+3zrFGyftBDJTV5TSPCORhJpgPIuLcID4ZSxXPB9Bh9F0KC
+PMMVradnS8WvoGgHm+M65lkjuUEAzX9xRATGBkU8UkAXjWeOmoTjaqLYxZjkUS+
FW1LJ69bHGcQwzt4Zu5Ua1ukz8Cyk6B4kUl4NH4wKiXrugSCrJ3BYYemDRlkutBu
8QycN2E1L5ZSpT9lkPxveQ9kP9KHVY2LwaOdxQCrP9WanH6GpVJd5cPcRUI5GB0C
CZ9snMczUKoVi+iAp/1IKWYKwXUoSS1NalO0TAsBiWI89Ed/YoYX3npWbFo7st5h
L6Vr1UmKe9cb+XaFTJh+miOlgun0sP1mDUDj4u2VxJg4L1yA2MXFw2kJeTqVCTEo
tfaLJfONu2etsEMPfngeAYxCWDimkZCEbf9FqvlCVW+UGmkGHn38uaErF14GaA0u
0v0g6f3y/321sRzWYs9qiaC7g5ntE/qvROTOwpx7lt6zexJRvfuztznq/KiC/+SD
TCKUHV2nHgth0UF1p/jBLmX5tfVp/iyyz+C++o/CcjSnZHO1F39Nj0wCDwiq5VdC
xX75AFKfcIVnklHUTpopS8eXNqQX/DG0XlwQF2X9VI+0onTVAh/dz2ymiRj0aoua
6mv3cKW3A0SUZTjYX+OSRDwGzsIhdfccp7DkR1iNAC24Skfju2cWlQFvF5IHfkst
XEKbL1Q8KFaI7OQjSgmRe5eQRh/g3GS/lgbrGZzZb3WeACyHT5DRNQ0UV8hvhG+0
Bcbr0QoxIc5yrGirzjsV+Z4NWY70MZXnGFX5hrjk6TjYVhYlCyVwllS6HLqYj+FF
voEFaKcm5NBVexH6ZkJ8If7dhqVEcdMmudWRRB+G+joGsqETGK6wRzwhG6mc0hV9
wm9E0zM+Gyq20EaTdEmo7/07plNvATvdspDcQ5jtQ7/3vBFEwqDYoZb+tR4rfyT+
bnG7cfL/L60xticIhpBtrEJujDuarc4lSqRUGsrkUDPa17ET8uLyGpN9W9sqFOqg
JxI329onOlaAOTBN5rVSik5k3wj+70ZTX/jZDT3kXhefeNbNwCwWw/UhH3GrKSMj
6S0yTOL//fSrwn1nniz8uhdrsHeueC6X+kOsfippqVBgTBMsOMzOjhpkygO+YTdQ
jtuK1s+GAivF94gkwYnBMU6eoSG5+5z0csdG8f2buBKaksezlPgl02yQBJaeAII5
cR2eMrYEZHIhjaMN43URkixOrSDDrrTr+HR4Vge9kDroMviVs4IiWAfVpls1l9m3
0ukDHZkoppnQPVEZyQMcX9xDPGr6BxYCRKE9w3k1wRa5Ui4HpylEwr5XoBT5WJzL
KdUT0PDzgq7nsHA8naqGCjDk/lfmFkkWG1rilhBTPRZDA6D9kTLjsjP8sLL+hwvN
KB55eIDw5QiOneOVMebomN2MM4wulVZFUfmTAkAb7TMm3I5eMUSvLvkKjn6mDa/Y
qpVgFyscBEqpAm90KhVFRGkkV334g2XLGaMpGm/mmRWdFR4mW4QBkZKmap56rova
3YVtSBcGmg/PM48XgU38PwPtZiPVuX55Jv8EAiQOg5QxCSvHkU2azR+5o8+700wx
2boG1vPp/c/p8PyHbNm5PvmmKvs3rpmrRvMhBR9iVM2/ElFbZSfFyEMW593/RUXT
xpOv5WZa2LzXq8BLNUzZr9iYg/+yYtxU9BQR63GHaMgA8PPvBOfBDE8BAgAqqhlf
gF9WMD0dREiQgQhsmRpJpiI4vIDkd6DwUW10Xq9IHt/52M0u5+mO4u3Gnm9W2g4Y
0qsXfeGvZXk7niGArNYx6F0HCbQOyJN8iCrJAe3dC5kQgSCzSS/PSumdnWj6Ij0W
EHAEe98gxOs2yVeE240gxiwDObQIDf6u69fI1qOzrmDVWzmbDNGr8zVVQJX9YYlB
9K0kH80fAgd/tXxU7gs2TXaPiyoTrFvzKg5UNbTtVxps1pBvqBugroQmHKqbba5w
7W8STxYz6Fd5ZZCPMNENvPTVpEVDPMaT4cxeb35nyJOND1oobpB/oIgAbt9t/e49
EeGy6O7AYPL963s5Yed9MDTE2cKq3VP5qLhNVrYZMoTZg+HRWe+CNrR85cIpQj60
YcDor2B8kyhwtWQ6wjKcaLRKqt2ihtDrGtpE3zwNawyfW73iyQX6mm1vatngVlon
SZ9ZiBcICCYaqRVNnj3MV8UFuXKnQDNFs9/IYfmk6+Kb8dEx75WQzCGr+PKevAiv
gBpeuLUtE06Qm4JOWktCmbXzajiAXvToi8RIwTgYnkcfdycDY/tzJcEtTmvPhpGc
reRK2aqkpupx2rFIQcBX9Q==
`protect END_PROTECTED
