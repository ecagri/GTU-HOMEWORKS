`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Pr8jNG+MfXNHCZKGadCLUTiBEP8CyRdhSWtf+RE6E3cJyr9JNFUxFLj2QGfCRy4
CSGRhyAO/TRn7v8XK+toUbea9fD4vUw3nb1ZG2saW3Byi8LbS3KyU3UzJ8VIMUoe
In1raxEN3Xmz9u8euo6Ah8ed9aUC3Ykr8Ea8pd+Ii7Wla9+FKgfdwpIvupy9CsZb
4qakGXtbjqAzWAT2qWxI5i9+nn7KIZJ3J27kK1SkM7mWaeGBh6nu+Nl1ssg9FRK5
/8KgIoeDo+YvBJGOtzH1cDSifgQtIGbC5RCdlmyBSKA/3Wo3i8+NKz62a5WSJ3Fq
gxxVniAPzmaHSxKWtthLJro7CYCGy9dke82c8fsICyWeaBpqhcKTqZPFdXCVTRqH
9yJOTQF3QPWG/z17fQUUdyR3Om1wLSQpSxkphsjsa741KiMBOQnSyL/sGx73NFiA
ni/HXalLckMun8XTFFTLjB/Q4fmDGeJoCn8mD4itS6ddRECJ5coXfyJo2jpT6mPe
uvR28BM57JQ5ECavsvMRiqqI97MPqfKVz8WR/26BBc4ih2DrNhUUDWiAaQPItQ8O
dRlFM80myTZpqOUjIOm9xljhkXVraVHvIxy5lOwO4RWaUcXicC82k4gLgjkamSQh
E6BES5hdttG+VrnLCIvRsMY5mht9lZz6OYcmomXO/HyeJ94fgqsCNqfBzsMXmvNC
pdVzQiTW4bGUA2gURArMZ4RK+GqakfGSZ2P9ZCmqPlKLANg3lQbgtU2XDGvHE5jH
P1Iycu5SAf9koKRhqBP+WgRAZZh5JqJYvEB10fLn3lHDA5K/zAVSBIquaRosJs07
wpVd4/gEEU03cocv2uPY9Zm8AVPL0pMLf0UesCWijEBx31go7ZrWKeGT5epDE2Jc
jIjwt/8BADh4jnXxUos33R4L+UlDmA8KdwXIHSPEFvdGXlqDKIrpLNahLEWhg2k8
zDlMiqaASjfKjXoNOkNxdHhDRoKZmyiISBcngZgtdvpQ5WSbbc8xw7Nqxd+klRrU
yjwxNfsutP8p6pJOLhh3rykSktTg/2ufj5HdcbTrty78c29mLLufOo4RHGMCNa1z
gJwRbReizvhlvtr7PXOmXQZVwwcL+XgjZ6P49w3H+GG45ICUAXK92lWmiUvz39XY
cxGpQNoGyOICvRRLzLUCrdV6vydUiQs6vnlgsup2S9nR83Dn+WLvoQpuLGKM9SYq
SB9+6a2rnCIXgjjxVZPWGMGxhPJPsctevhSCPf2QFaCgcFUPNC/pfzsqKaCSpRkC
3ZQMhuN9zi03/Wysy+JXHYgL7wMZV2PF1PODgqjATWoO7jdQ7moAyN5AwcmBsmPv
qU3bSu9gZVJRSOXRP7HWOgKbgXbJShaJILlzSEqelB02+ETluXHUxcvJ2ZytYCGr
0HzVOGZ3R5iWdMHpWcvIQnVhUyz0rMd8EFtmkTTcuM5J/vVovI5/URieSzVzDC9H
`protect END_PROTECTED
