`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WTbmjqvc43Dtbf5u1N1GI5/RRv0gwns+Vf7ozi83KQyr1mx6pUe/yF2y/sJ6XvUg
9do6DYaHN7U+XEIMu3pnI2i2Isl5fDaQ62Z4OlLOroUA/W0TSWwJqIuVjy37BSHD
V6ZACry9qxqyJKxMpbW4qqGzu2wI6LYv+nqXBibsRrE9tqVeOxRF7l+VbJS0qI6M
Xm+565PP3fR23XLRbdr1NhAg5oTbJL/7H0jf6+KCLpKavEOMiYQRI1TXN7ujtpyh
avLoNbZ4QVP5z8WYyaH3exOUc7uo+qMteGv0Zk2Uygfc7luPdawvtvZ3InzLe0e9
uJZhYhO7DCTwrPKsf39xzVicr445T/3n7gG/DLA4HVN59D+7IIQsc67rELWqi4q/
0sF9Lshv9wAHFRKaZlkrW15Nnn1/lf1i/dx37/8KxSG1zl+2XDeQ32A+iG3NyQqY
6Pw7ChY//sJy8lOnntSLC3vVzxOU66tnRp9CTvc5nJeg8G9QYW/2qzQZaRta1XNo
JvqM994Dp4tDRjBxGZkppwobj2NRSimwd9LnZi9WAXWfnXJWPD9cohDqtWihnq5u
XMoyBF3H8yzY4aNUPEmuEq+kLi6S2npepOJlPdJGVeQEkYmbe3ZzQTh/u3oE8Hor
Tnux58fV7pI3L0hIXdkOQl+3iv7d8Q1fPWvpfhMzwQm3KLVjzn9iIogEaigGJCfN
d+dfeRMay9qOq++p6BMIG1R+jGsvSvG58HoZirn2JyF4xukaItdHjTEkGtrJGH8T
jiBwfUDLzLinh2gDrpAEAToaM0NVAVp/pcVGXWiGZXvvo39mARNwiO/8s8/1cxNp
jkrSsp7FcA+jDnJwUlfjyB/4T0Z1cD464HRUM5SoMxu+N5tiBwqLkKTcan7tz7/S
mMVMFx41Q+1M6D6qEH8q7HAT8UH8XiL9PYybnhpMAW2UeeyPbR36IMovQUcywsvp
6XoARlpdYzkFVCj9bTAlMq8V4wn8k/DNHI7tBNqLJihWbUlNiZpudi2BlhCqMVu2
pwGsexLIsyhCxD888V/oTFNFtRRNc/A1MO5gQ0Og8QdgODflmhx489sdr12c968C
sHQYZFoKUGtWVWFCRiPFH22YdXMm9eQvTtuFr8oURLBoLd6X9aoXsour5V+KI3Qx
j+24/Sp9bTxpkCMrQv3Xq620/1sok4wnb1jE0VcqlT1jFMRgjJsgx260KSq2bvkL
swvLRI1+vOOFXL8yDvD9OrMbiPb49U7Ckd7VMMkKInBwFAIDkuQh+UHKBSZOYi4a
Kj9tpBNAjPKi1ihnVmUF0e2zf6X8uums4pYJs6gdDTlFFKDqoZhjGUjMYUXKEaBq
vKH3374v2mCvc0Uk0XOWN+RkZEfnjAKYpGowIlpXrUN+8W2nR09cw4sxg95L9US1
2xIx58ZSZs/tqZ3DCvTdqp4ay83C7Lk4e7LzPJFlcAluBUGLc2O1kmfIlagOi1TU
z5JoJlufprrGbH5T/UReO/entfm1FB3Ys5dPTK+YI0CuzUJavkeylAbPL92mPWWF
gc+Lw4hHgwkDKbkHOTp3b6G9yFanREH6DsmlyZpdoV6KZWrUZHst9psm9q9OgUGH
01d4i/JFGchO7X9IotrZbDb7ypXzparcHcesflDkco0eKKaG2wHxTtQfOvFLEbyt
VVkQwT3Yygr4CcjhxZGo7shEgbyVtUKMGeTeh2EZ1NP2eBrDTz2ZqiRNA+SYeRQ1
LZYKAVFxJ28DRPIBcE+pHWlZDrJDKyJ6lUAsVSW5hYK0w6K6ymwguHOFnYPqkMGj
KVIoGzOfYzp7o3j95Et8qzLl0X635suxSiOnrJGsHZsi3UU66xFgoa7YHNhTsAEE
5JdR9Zouh9BZCsQLYCcfPg==
`protect END_PROTECTED
