`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yREVZPtemnGYwPnIY7DRxSgzc5jkQ6eK86EWJeaguLzat+9T8qoRez8nJhv8Cfye
ptM2F0YscjjNuHxHDvibw6tTD9HvoVHege5iGyIn0iCLyyiEvJHiEb8+xW9FnGFD
1Soc12WRYZePMNCAd9VCbPbno7nezYU6Vf1I6ph8xKO6RhpNNguTm4g5KkSp7vdA
3v8QoeyQE7MiCd36lJxOLgzM8HfFqEGDHkV9EeEFOhcUA/ifiP6IxU3IPqCRvxdY
BFuesCel0HpNHWpZetYQn9R7legb4vNV02Uv39wer2YazowIFMLpWaAc3Wi9RBNT
xfuceNVXajOQLSzSlM19fNjft0jb2783w+gITptq+qV+gi5wTDn2vBiZdFjKFGmV
EtPJsBxLXyWafpSAKJgRBt2dCldEzYktomriX0J4V/B+UYbJhlHsEjc+xUnne8P6
1PdhI4Sg6W4SqTKDa+eNmc5+sid2K1ivu1uV0dVKsKMoHam8kSmL4y40T0GpBjSV
dg2fAyi3b1AfTMJ9LHiYEMYeJXadiv+PasfJQUR9OlhtGFlp0yZcZR7jg6998i6r
dabu6j88qplkFB554BlFNfkIB4s08H8rtRTfqtwzFAVzzd3LZZm9Sm+tgQHiijn4
zprAs/Geb/DrQkwqoeAO0HIOSnmxgBnrWrbCYVxer0NQMLnKpkb5pyUMx9ExUsgw
BlRuZ72hhlv/oZuChz0bxacnm5y8ceEgpi9u24P6fdSLIi/brd+neTy6MjQv87jN
ExRgV6AN1TJs7+Zb9JDafYIM4Dt5W/kFSJ3YmnTpFRU2FBtpL+Gx8VxB4tvsBz8I
hGQ9ezzfCfXwfyDd8O93+Irp8viBb0cLzwP4Pxesc3eJ/CTE2tIhERZ15o8Fm1vK
UpoK8ooKFUWsafpJcJs85bYmoppcn2SUnF1LG9q7oPt7uFoPCYsWQFbBy4bylxkQ
oXqUyVomUfnTnQmwS20mRp2aj1WHoFgmERELcAvq2vWNwph9KX0FgpwC9bN2dwo3
MYnHNkjLqoP/PEHOgnUji6/1eHe0EoLGHJ2ZSQ41mmqzXwIejl+krwNLYRWnZikU
lzyWNUwUrMx8Cb93IDID2gj2ssE6fgvcRs6TOBQWHpBdJZjEc2DidY9doUTs1/+9
RtPEgw7zW1wMe/Zau2Y9JIl6wemdEGtdqG3O2gB/WYDT+Bc9ERqxYXB5HtKPRh2v
e+nw1R70fnTrCQdVYuimty/hmUDrtQL1hWck6Lzp5AS6BeXV5al5y0rvi2wUt3gk
Cu5QBSRWujyGbp513pDNBthXrmMc3Yw/Mw3FbEddYT4/kI6x40amzHzodhrlQXZ7
gqE6UXj5mRF1h8fwBY08Rzv/3S/c2DWE5RASOv6zK1NBl2qYB3EQ7exL1GPqYpr5
47Hgu+eSxjM/jYmS+tA/DEo3w3YwzP48E4+JunwjHzA+0jcAEVmcOiT3WT7qpKJG
p2hzF4jtP6Jl/Yr+A+tJ5wpJnd6+UVg3SnbLvsZOcXdO6PHupMQ/Bv/eFb3Hav8Q
KwvgyXT1aj3MlxEKiKBW5tuXY3mfPJN9I+ihJwFJLMaUXXKKxIrKS9eEf7vDtpnP
SHZD5iIPvK+ATTqKbOH37e9MHaYcoHNm7czm3hjiyn4b6RXm40fVAeqJKxoKys5O
WwtRPehkaKkRlmrAZAurXtOYzCtsO+rQychCXtNwUPBmYz4e5OfCPt5Xw+9TUsOx
5C5XX10829+flE9WB8Pgl3b5qMKyAQkuUU6krSILcuDkaHGRF2pHavCzODOws5E+
/UQAssr+TSSnivrPaWTOX77Yk4R68HxQsoQkp+1jkAqycAETXJV9N1QQPPqGRRNs
fFy9J4Q/P2dArtHubmuI4Gfjsz7J2lv/pWYSfIMvAUE1LPCQZ2DQ6Dp7bAh5TJdh
bzPtqgmOQhtU+AOWx9388DuS7Zeedpu5xyNl9S088rhlPuWjYm3kHkNSFHCsS1I/
oarED4cFtzYzDc/SBvlUkDkPtjR4FXWMzt8014b109LbuxTQhtdCsoQtROtPFBpb
UXwA/wsj3GGsMtyQgSDbFVL2lxWng8lVGFsJ9VPH9Ru08O6sE6lZZJnh/n8lM33B
f1xb9z57Xbqawb+4oOW8zxpL0hR/A9ReH/m+L0keQPBy4ZPe5gcQH/XJOkkKZRWs
h97ucPYYDYxEr7RbMOCkHVf9qFHH7f1OpFTtl/r+/XIOKtIf6L12H0/L/IHNVVlC
BgZr/wrztbolmrLm1E9V4hRg/9vDdtAlZbW2d42td/3OX3U3va7tGQmwHZFonvT5
r3WdkMhZhqkv4BpzpcQ0Cc80G0qCWC90XUXvryKcEvO7qRBRSh24noOyKKEUIJ+T
Uyp0Z9IsgslH2JMkwnXFxFRsWSArJzKS7IuY/vrsCMgYkfBE789grRCwA3Zwauwe
CYEPGcu88MSQq+cmWzwWn8F5d2iQCLG76jjR6LWtqTckzAJIc3H0IKnmTJ9e8VUl
zX5f49dOEmSQLaxCKhXoWy8Y/5gk9qVkJeFu7tVU3W4dKEaErTtu+t1TA559u7rl
2M2/Std6HJ0s/wI3snKgDhohm3wK5C9RyagNxYhUlUMMYVPicu6Zd5bZvkBFVmmO
lAPyTH9XcXhwVhIeO3np7g==
`protect END_PROTECTED
