`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
whUvWh/IC7YBZDIw1+4VBHSvzO9kmhc+GzrERXJyCbsvIe6MiaHMEjHeH2aUHWaE
WFy+q1CIYx9JPyFu+G/YbCvX9OtOf7/44Dyd2+30TAQzKDlyNibRZVRFGk2f9yn/
a02AMAu8JToT13gRecNvDT2lwUgmWLt/uzNv0HUHosWwnw7VBHiqqO77xgvyIjm1
7Z2uYwUjMLQQbGokcI8RFvk4SDXSMhbhXWYd2RDE90rbIaGRJgoiScmqlIVl1seJ
g9W4/8kiXOY2lJB/B/6Ef3fDMDTZcNaKXEL7DYs8+r6AecFtD0aS1f105e9OeG8r
ARzepDrNSm1oqpIUq24kbT9hLhlBMWYt1FieXqOaPxFowUvhXGHP339qzkKh8h1w
fml5M4MsuKtWTDFGgHKp7Uwubp7E5SwHC6DvHubw4lIq/7QtLvj/TTMDwpLoOrlt
zM6/XbWCGwylbO17TO5tbKBRCQTSUwReUN1L4Sw1x6VeJjc5lpqDC4mI50wa1xEd
TQ5YUTcsWsQzSjDzWoAOrCy9GfkK5O0sVYhD7XQVT/zdQ1x536x+wwHYVzs88lqY
d2UBIsFYwf7cLh2Owb2Yu4HZQiXECwHZO+PmjnfA6LWDxJ1p/42vcKsYwgctGRyp
JYc808BaWwdnnitrK9+IP3GEsmqsMhB0vHbxxH8Dj2fwyCRa0DUYhQVlymTWW+Lv
S0g5BajctIiP3kKasjdat8vShY/H3avEAR3Jcfz5esWy0fzSS2rcGZNjId5Jl41L
astlWT3A0REZEtd4L38gIFGkvpzMr1mTGP8Yh6nEwiWPIzmYN/fNXeFesKWmOKDP
H7Ca5MBv41LQ/zJIA7NJ92bsvAWaTm+mPHrsx7QyARjh5Vt2SuTbx7dC81QvoRPA
o75LjU+eLZzSm4nZo6DIsl5kHdUJA06TTCOqimOSpqrUdebmfo0p8pI9wmfOG31I
9WPr0tUDuaukYYEmvyv/YKyXo9IVA2anlO5C3qSJuC7GCcVDdgDSIw4DpoTCe8g8
6v4qjE+BViz5NFaJwS+f1QZozW3G9W+JsqiBaPj3CKCHpavQ+TnoN/7Eo7Csdujo
wUMg+BkARGNaC60qbScUzIV0AWEvmAvnoqKWHltgIs287LDbvp2hvbxceE1kMcqj
vMd/L9B47iuRrN6fmfLHjfNbFkUbYW7jhKQlxSoA1PtPyoH1SKE1Mdo1gLHOHc8k
Yck1O5wEe3Poe9zd54ke4QO+orkpJ48MWh8fTYpQ6XzdfWpLlSRYzqiR8Fsu/ZhI
PAdZvDyuqCFQhf0KZwfHi5jUlLo/hSpvxhLkEyf+eXLsTWpm8B7attcy91gDogYg
muilUXn0A8ckz3Q3m9x/LY+ZIkE445IZOJztk21M+Aw70PrAf2IY+qAAcpB4erq0
`protect END_PROTECTED
