`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QJd6dkc2AtZWPZRSq8buzPjxmf4jCvBkyPE4jdDdZZ5Q06hCFsxxdEaCI7zJpxKM
cRsYu200jzEU3Er6Wqsxnt6YLcDLw1PEDwNZoHugu5xfNQaOgCyz0/GbOM51wVhK
HP6bMBrMckk70U3JnquyaeS4QCe4JgzFXPNSZGw6Aaql0yvHZFRG/fVZzLg1MsYh
g2//lhlgC4oa/5kGsBptmmFh5PsA/kf1g6XLo1gWFi4VjhDjcg5jKm7qgi883VDu
eXgBOXbbfSq6jUnFh8MzgUAsa6ZPkGfQsXEkeTolNKs+ncewNHuEdSG3cn435HDA
QzkJAEad40M+EfdemAAwj7i9p/hIhQq365q5FH/Na0BISEuYwKI+TPqk/vdtF7h6
gedVZ9KqPuG1ADKmJMXJ2jk1I8pFtnoLsvKCdI7Ih3ItK2NqGSLvbQRnxGXyOsiP
HO8WX1r/v24+u+lrT4zvgJMXSorPupTv9kwWcd+PsJy7m3Ypq++TgGxMaxxpi4HI
0SQywSFcK119DuvoJAob8uIVN2dtOiV6ttC8h/J/hO/NxzOVcOAcS4o2cTd7aaja
QJQM7rCpnLVudbUfXil57ceDMgZ/Bn+ApZthyM+j4kDY9XFQGV+RgSbtaCvk8OY/
cl2xmbhDhJ155lXcn0du6Nd2ojhRANTd/D/5kb9MkBsiERx2k5MCTaXOyz+oYRn4
MYNNJ1LqrM7k3Uo+ow3LPV7I+WSMXeB38majehfh5JqYN2aim6cIdNjYWHorDVt9
ByhxLVk4lWoTYJoGoNvofw==
`protect END_PROTECTED
