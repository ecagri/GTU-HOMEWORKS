`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K9hlSc2nzy9vAd/S0wfq/+FWw0+CFcmVzwOBknh0zNlQwOzgu905ersqIlC6YJNC
zSO+8igWunLvBR4Oqd/a9dBiwdipQdu0YzJDSV2KRGCnintd1/VSlbY3GGiTfv7F
nv+tsYqf0v+qgw2a5KIjl4Qv46aQ2k290UntcFcFjAaVMaBqv1OXDXEkKr/YOrAh
CY00yZmpPks6Y38REy2bFq4Q/P0WpbQfw4J2ZherxUJOjuodCehqkjEUmht+6ijl
0McYVuPoy3WBpq4yknPsImUWFERdxhpI+JMR4Mm+DSwMRgJtn1xXfGfQk2EptPpl
qVbgHUrbYrI0KVy2+k1Nxz78A7cQsf1i/n/pooKsfMbsEEEieLyFDcB4LXhl6mWP
W7xnaMMBrAdtMRiMZyhAbWi2WJl06OxhE3Yizz3QU5+QH0zUDfHvO7FpNf09Z6e2
cJLbuHBBHskNG4lxJgfKKG2nmMlgfq1KZObZ6vCCFz26rE9sYe4REkvJ64kJ+IKa
mrS+7AJs1Suv5yS14gaiZBKlB52p8IzmKTKvHTlir+KI2ulO26b8/TueEfZBnC36
dWN1VOyAjzuD982EzEGUL7MoOnPGMKDVQ5yM1UHIbEsnbZMcQ48LPfG74L6e/qHA
1eHzMgYjmAqnCswTG+bSIqaQ6NMlHwLnfTfTs1TJCt6KJ0ZHrOWnKMQAkJxEX6fW
hx79o9oI8+IynEMgRWRgBV/hyn3TCEnu6zz0D42UmHAHV1L2i4R+dnFtgTfiLW0Q
9A2RtC0/hodcvVORebm9mDpVDDFfRhek0S0wA2/yuTMnbN4mhbEYUVzSvscI6fLX
SXptYDvIGY4A7gRDxSvH5rvgKHQUh2HVY/DFJXKuGUUE7wQWj45cAO7Q4fp9B9FD
Cucu4nJKnrJpmR1A/QUyQh97LffbnlOmzw8xpKDSzrQ=
`protect END_PROTECTED
