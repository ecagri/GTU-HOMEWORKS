`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jND7tTGDdeya4WWDOl1An4IUFiWkOaqcPgCT2z6OSHmzuOaKz+DH3XAsvm/3sSYm
5YXVIi53Fs1nIRhxinhB2YXP1Q5jHNw2vu98aiYFIWfB0sDmXDBHytoUNm47YQCZ
A2UEz2/UHT01arZt2utNa3ywiIXOSN/E3JC7vXLwwa08SGDKTp6kYIfwYbcE+Tiw
Pt+FY7rMasCvu4TdKfQEhYajEp8Uv4Oro8yNz4LcHsb4E6WUvK/Stwyh8lKmMUhg
iHUYVxpMQd38ZoE1Dk6QgHZL4jQwBha3HBtKPbt/opJ+3L/lnL2A2bBIEIwJft8M
Q5e3dg/znULWuCwztCbhGs+pb3bfUNGCDaqDz7Ex6NFLAHKZOSHq7pvD2xz9LP4f
bUSKM35oWRgBnKRH+C3Cs/7XV1cgXEM403O1Y/IoUWlOGr3DRruowOzTrk5LRlos
dvkUvAU+n/UhoJMLEjdA4rOHwv8EsUdTRKtfRHj1zZUtzij/f+352dPBmN32L2iS
c5r5wlKQ1U0Nfn677nr7D/B2wCWEWmxVcvC7+LzlI57c7CCU7oJg59eqntaxsLKt
RlFwE1QnTl3d/gHswUiSPi7vQZOK9h1Hjc/XxyOHWMKR0xeFDdFgcDOLD92BtjtG
Zcs/kO0KYQ+2gd/HfTL7mx9aQ+8aBuYsr9WpqJc7CRJll+jJYwiHW6bT4II9wvgY
gt1g0jvgihGSi85FWe/ENckNTI2JGnAmMzs+/S4HjGcg2UKBikpvbcOOUykXrR4x
tqZzPSJCPJoWCr6iUC5PBMiqw7fvaAKyhNVEFKclSeD7fWzLwA89Jl9aVlbhuaSB
I4xsK4RNr9dbFmIO6FeZa4GeVVOjKu/nHluqXZiPrkh+pckD37PzPJetHblwZlQo
pRowFXAhHsnxwb8PPkEjCMJCP8U8n7/hPfI8+EVAUB3+IZJ3QBBFy+wkQ7GyPtjk
jGtPERKeBgOQM8VNpSU9QceN9O40dX8bpeq3vSqXUgEeZ6xBvjTd3dzOdNj5pwlP
MdO/2cWD9MyPumzhfzXqX0koLZl7S7/f9o/YiES9AsIxlv9jt9PppgWuZFSLzzJK
mDLw+2hKHkHZxZbcgL79yVfCZaDm1E30j9DryELYrh1d/PvqbyqsGzqHT7iFd3rm
wCes+poJ4W2nrO35R7+KdlzJEf1/yBq4II9/voYpMTRuTU63zXRSlpyIiqWFfr9u
HDVoGaJFBFr8kfQA9NiA0kyO812xTaCyou79pO0q2WbZ5G7YDlpnR5ZqeDwjPtZV
2Zj1zhJmrQBnIEIDx0AQ84ONxPiKn6SvaOSW2K3GW6sbuHV358QwhkDn3E6qguA2
P2z1DunKX9JOlD5RreYihjuff7PS6EqeW2n9JY8gBUXJYAb2ISqEFPVXjdy2DYsE
cekID+rcSbdh79/jy0eIVNDiOVcmy/HLjZ13z6dclhQ/RxpC40YxfDnCBtsZd4F/
bBDalT52bGdKCdotxEjHuWdkrfVdy4CIA70MBUvwD7XJjiHOxC0UqibkMhGnsed4
MOp97CNM4MZbpUBygMqUJdqkt/icvfcKf4jmFDqToa7ybw6XCWj7g1i+EUxhL/UO
+OPhqyLqx/M0nDOlGGj8TNCXq/lMzrmr6TU+nQU/BgG500z2mjlafqui43t5nE6q
36oDQjL12BkjOjLNslMmGIKuNIISIstZnuhDYgpmOryleSzC0X8lONuR1mVbmk76
ESQCpmIF8LP+c0N7mleT0v++xhV+IbkBoBAzV8FVFr6aEmmHaSdDiaQLU5IrdGdL
lk6SaAvmNKfDtmhdfotn1MoBGoMauNYRHj8300zTQHYJXQgT6YNWiTEqJVqcnlSL
ASFjUl1s6avGT3vEMAVO7f3Vt3RcvoQNlnLFOU/QzpE2I7jLzDnlAy+JVeIqNbrq
s/9Cxn/jRDhqkvQSgmWy2dMkZ9owkD3rZv7BaakaRfrlhfwdIqsAQKgiRcGNTsUf
fmcJsRYCzPkvHlBIHTE23US80qeChMiOWs1O0TMZNLE8whDVw14fj77PLAfRrayw
`protect END_PROTECTED
