`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IDJ+DgA8d40WNz/vL52Aa+Ed0Ebt5HiH4z/IQauR2RlFg5c2Wb9uPttavR/Uv5Ah
6QZiovoZrPwh//PKiC+nJefguGsKVSCkEWIVXkQ6YtIcwkj6IHsrj3ylVHGjl/Mz
DdFajaXDnfrsR8hkvAGvqycTq+25qGGBr8oHcdsMb2ItL1Pm3Q1V1rf2yOf4veb7
qN8GanE2zv/o8ewFeZUA8V0DvBSKz18U+2xxvqgfjhjhUlOuuC/m3exsmu6Fxh5Z
oxElZyTbPBxqKqYfSGKNoWFZ/Ly3hD8w85c9eej33KjVBDumzoDqvpO14+LphGAO
zg7yfz5W/FNqeLmrVy1SqsZp4G8HVKf82ZFr3eYQBI2uc4ihxzVT/n0YuyMC2I3p
vQk5OPM85oyi2Ly06NtO1jPpajaIx2lsSsJdppwXmXQ9SUwFbrRoDyRdMWjWEOvU
9De8SKFU6+QqTN4lEGrJRrpi8NsSZHkvuVhYu88CIjVnMX/+3JHNQWdRGh0pthfz
S8cWdqEBZSDYxfyYkzcGbpbbyzvCAPTUvr3rdk0d1B+KchMX/LaTJ4T9K50I47Ih
+rs+Eb6pZmYkIcYEhANVdsfzrTAX+4wkf91889aEdtWHvpEgNHSlJ/59trc5Abrf
NSpg/SArgbEMU+AvewFom9ueF/FiVjzycmrIVkXs4vZ6fCVi1LRQFwBrCbJ8YS7O
phbwJiOG3PWzGC5/8dBDGX0wOazPFsTi+UK4riZwoiGq3rexVXQ/eb2Z59r2fpht
30vtzJEV0NNwQ5d34uhYY7z/qyU614GfFNBzHOQ1r0KqcMYYKrKEfvU4dU9DTOdc
Vb7538Ei9g6QZKABJK8jqKESK6t49pWHUNtxCntc8YDXqqvlfldlNQzZ0XsDp0LF
ewPA6uGErppyCbQtpjWTAXos3nTrh67vy5Lc0i8/CaCNhAYZoQ6zPDNtsQwJ/3mb
0AKn+JS0tx2RzrJRUXpYgnm1nva0Rf4wfsvBr136aw1B7Gt2ubOfAnSW+bD7C9iQ
Jnk9JjBE7mdBHORN0u5ggEgeAdAo+qpkMjfAoj1IjmcwdlONuJB3WLD9DD9645lU
N95uKqJuER5Vwifski0geFjc8CGK3fX0p0iLpU0ZcYxyH0xAYGi9qXwumuzkx9DR
M+DWDvtm4UFuuKV4aW1XQRmwoC07XMLZvkb9wgPYGTxe/le/Sb5G8LdAKLeBfkOv
UMBqCHtjc8V8qjqjaiNqKSF/vRKxAPtwJbcVZNCI7ehb+o7O1cMVF7nEt/3YG+JU
AbB485Xzxph0XYYVv7Hnz9NBtKoGVRQt6lPF2UpWACwG4IJ7SfNLQnv6VYbx6nON
yEQEFoW1/i3wKibPDQDmkCNal+iR5yXSjnAaRoobceRwcxwBFW0bn2KLogl1HvEo
AmI9g7T2T3n9Em1vlpbXdW/JHPQdLAz8ofsUnl2KGshs3HA2wD7Udgn8Ixl5yU9U
MPN4BJtocQPgZ6zHwYcL2GFyzClKT0NL4pS4fmVz+Avu6L59bCCmTfR9Q2JgH4bR
PEqUKeTuYRgzkcebK5mO6mMa9JKp35JLhx3M2si8QRQnjoyHJyEAIGiBY0t0pM2+
DjM2yFUkUA0Z1y7A1ubVzn2KRpF+phJfADwHX0pOeS7tqwY+MfhQHPhqbUU1UOMs
XpkgVNGcGCOarSi5oE3ORov1JN16/de7SogG7IU8xg1lVxzXCtjRgDlTktWZd6/1
ShdsLO6JEyp3uTmh6ZLUpElGOBJ8PJcO8d+E6du75ckNrnKz5FnjLE5T3B2TX2QL
R2wOmVwnZzVly9T2ZEkd3hGn4vD/xOLstLz+XauSq10GKCWLge9QH3dr9g6UdOqm
yIBEBaWyrFiFgJQneM9SrNOiNYLSO0Ni891TGoc3ZfqM6/19M62ooqHhf8Ba9dgi
iXHlKz/+bFvpvp8mjiTmjz0aTZ40XplB46bK/Wd23M8r7RP6AkIS6FsHpXuichVE
l2kvDEL2i7bH2wMYo1U6DcCgs4UI+Sb3tYMBwlFivGrOCcfEfPbt6F3XvrRZCTBo
RksjSR0j9UZk6TmRFdn0rk9W+O6/xg9tNdgZZ2X1ZdSs+IgDnZ88CL5F7rLRinhR
7XQ2bui3uR5M4xC3sYEgKFPKy6QVvaNO4Mgoq2BBwdzPQQ1tEEulwV27y0Prc0di
Y4jcRHdDQpyJqpfSIa3OQ56O53OxkTTVebECvqt7VVgLXGTwp7u7gin2chJ0uwAR
61Rmny+tL4yEJO9mU60bYgme2FhWtUUaaZnhoh6CgRMkqLAYZceW2qbQuZHNqOrN
ukvfiCkJ5VB1pyEXPJTtn2yskDfrje6OO43CKxV6939IvHvo3/XkXoh0GmgBbkgZ
jCZrFLFqV95hE+ur8j29dL8S/OuioTn8vKm+B2b40c7XstXJhYpREgP0OYFLgMK0
/M1O+jJb5BtOhf5rEZ1LHrMj7/TY05UCoh490JrA2+rxMxM+EMj20fT4L28uHLFv
LcIjsFF3KEBtBOqEhcJ2ssNc8JurqtqRu307/Qr91838uzZN1aeixZ59EA4/w3kF
LenarbAuLO3ui6oAaMJ0jcWwxnzqfdRcJ26b4FpNs3xutauZu5Zn3w5btXQi7YOU
gUslZnYwSkXAiiprqZSf6oaHcCTV5ZQLBFipHwmzBBAYPhXsxjygns4+hq9ZdPbA
/nuTfgo2RkhWoTBsu9iT7TRdwn3HPBFagJHchlvPQ7SVEb29t7Iy1yMlelwCR3ej
FFQcc+8N1Or+4CmcgnldpNH0Shax9h6tvLjICEdB1D9ZRUyRpvjItlfYPpNosnUX
V2mXi5AN7YzeC+Yo3LQoVXaU+WSFOU65U/qwJyNKf82QJ/9ulEIp7/W+DdQxmpUZ
olpu2tRkJuLU2HF74q/TE13mkBa6WQ+qrfByt21PZT6UoKYBzmDflwfk5Xrs4MF5
Kri1FZWiJX5TNF07uDDpJ8hzjeihq3oT9Qij2hYrUYYZIT8vyGkPOKns7VUSvNvx
st1+P6wsR7m2t6SOr6yKxq6u0woQGsNd2C1WVIb0TBo1uD6mU3hypGULOvWuf80k
3njUEk/K6tYOis9J/OckWz+hdm34iFrlmayYLG5c8qruh2efvqufOjdUI9BG7RLA
OUEHiudThAzmFAwY01xRFSB1pugl16qfEhkryY+el0d3XVm2pn7m76uIZUwGXROY
O1mldOVpSfbkCYGrQYAsVljQeL2OD9aMrxEhfT1t7hdiCPrKexwM9n/CPB933uEG
qfZhnULgkvtHSZJZhxL5q+HuqpgTmvnD2IYAyEVXipW4Yhbvyr0TRF95km+MEYot
Xb558k1ydP3UNLagN2NW1QXiDnv0Lm2q6PxFVXA1Th7ClBdta9XTbigEYfUghGK+
BD0HPR4RBhp6DbVEFQACTei75s2K/7jZRapALOSnebJB/oVuV0YDnBFS9bDbGc0D
hCl9e5rapS/A53bgMM7R/+9lRPBHsCMMNh7o+06pToNloFYSIDBnvZtnYmniDQsn
eHd38kZypnldS1zLT+/kOvlAf5qdN3ILItDgSyZAV9n/CFdGNOqHvmWwXo9mT0AF
S90isvQI9Qdg7zZ5W1TWr4kz5vVhBr44i/LvcxbmGEfUC7v78H44LK5SoI2O++AU
eHlSRPWZr2vFqBnfgCKaSi3/04xrlQcodAFN5P6zFnDJcfLxWaNXLoZU8p9yo0mF
ivWhdXnOqLJ4PjSt2BFegWAvlaIHbDu6gOsvoJ56CofwATc80DZnUrHTwLsd4/yZ
zVZpnFce9Noru1d6/rZBwb/xzdCk6x+5JrjkuoU5AL9hbuCBaAQl95+nj6aavAeq
sBfkWX+zoOGsQHThtZ1hz4JFPaAb4PhmIxD5kDo42wiYHpsQNyV7m5aR3GAsfsb7
ZHaUV1JBV/Lqzr1n24bFABGeuWG6t+7d0pxZyTXJ5izQXKF2V/xRdUwBhk4HUuYd
JoNGf2vq0PIOvUHzLqMr6Kh5uUxl+A3mN/wcyk40bX3Kh7YQoMICMQpwJD2gJ79T
NBWIMtuVsej/+kEbtiX072ZTSRj7uWb1ylJZk5wj35wmuVkII/yKMcqTiUHgB7bn
cMfRiA5ga0sqdmQk8Ytetm3TfAsla3ntoUWkySaVJseF1hz5tH0nueaE3QXOmNuj
kztr+Gz2y/9fYzg2Wx5sBpQZrEreCyZS+au0NVlcfUil8pSvB26gqGgD6/P7LJNc
REkFEEq+zxn9frLP6KFCjMxdkc1D6Y59ZOxnXzCH7L1g3C35b4mCxUJe7hFsM4ET
qQqEHLWv1P8mDs1CkHwyQpe88jf4BaM6jOEfcUB4npAVIcowhthN4+5Lfk8E2J2S
VtiLTjz9zyS7Z+fqtl9TwkDQEFKtUeVXi3GtGe2abZ+bjwpYuZLGsnGr+UZDnOs2
+v9meCmrI5jNf6vdQhYIhuBI3uy3t9rYA9wWqsc1cAG6D8PJ+/MioNDQZLnqiRKV
DyTS6mY/gVa5aEKIoOBySJqbGrfKPzkp64+aJf+pCoVlAjrnm8dG44IoeS8kX5Ds
JpQ4kOVIVI8joRG0ZNeqfcTz5ulQye6o7i787QEc68NsBJuyiD19nzBltmpGpl6h
RdfRetxo1CufC5gCCehQrRUguR8aN3gCboSDTma3NlrGkieww04rRdILWCraEZbt
Bmge1U+R4q2eOwB8wbJdBT99g/Zq1qAIjXOF4GoqCOYyqJfPAl6Ycgm6Z2LGR1Ex
9l+2ugPHgNHHvSaBIiHJkF2P0POH2p4CsQpLCbGg7yzVFqvphAi/viVte0tu6I1A
K4hNdVxt/MxLL5q6fBfvghuOzYC/Nmn0rOaWIkIZq946LQvkk1vF2yVaicM/8GOs
M47QohR96PGVeviOcdF/wbCCozBbHFeZMZ0vdoPdD2YsBhU6alEJVKg9c4K1qyxb
TVo4YVGo0ZNf0nkgauVGI/b+9TsyrDwZmDWfUd1LnBes9DTjTuHIrXP6lAz43hNW
2CgzOk/BV+N1/stoBNHEQ7Yma/4nisRboX1HQxGVUektr0pjoyjaKpphSy2cKXy2
y9h6GSTUdynVTcsoVmrF1VdxtuBclz8lKmF9akM10qObB+BKacJlURoXvPlFQD0O
`protect END_PROTECTED
