`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mixqXqwF53AgGq/xAIwUrUsdhshuZrK+LG928uD7iux3KXtbOgTCuzOWZW/8FJWg
sR+kCig6VK9KA7R1TmlVzs4yGbntCfI5ek6yA5B3r5wvQbdvG8IZWX8ZmfmuqdqG
mvcjAgRJp2y31aJpPv1tOsZx8fXFD7r9BDSWIiZDHxOAYf5lUSOdj4BBMx5jl/E1
wi70vEouZAh14tSIO0P6pXr6mIEAi94sm84yKcEQq4AKuMOlSq8xSm9ujJKF6c49
2YVSZIIyN+iYDKcWncxuhO0x71kZvaHOaD4miu0s/RaVQox+v3hI8l3YAz6vywXw
TNt3u/phikCfzbb9jxS4dnNn32SAHY5YnCgihJ50VIrxr0Vcag8zE6c/6dCdhNjd
wuNU0m4gHoMfGPKcXaEjJSxkXrQsUYPlpBi1ELk21pUiuS2e9rcqceshueXJGFxu
/dQD3l1f178x7G9k0QzTI0QeVbIufeER/zVFxYMkP1FF6fAqiLD1sEoFgHzlA1bd
B9CcsjAkvRpH5j/N7gy+MeaniIO2LShqjp18bRoSKuajJ/8a6Nh4Sa+gSU0dWXjs
GOZQ9/Y07rCuBFsW5FZV18dIVmjKTzCrUZd0w8bIDZnSA2kEfZmfB5NzRz5cdW3L
WBvoupNilzZZ8cUdpmgt5XEhjhEEY/5pZVcKuZnYHuB6hFbQG63HNl92gAUwX8+1
xw2uhq7EBIeBb89pDiWlO8CJElsfmaBcAZhzbmzC8hARIe0FsegjlPyzBl1O1DmI
2nqhfd9I1s0IKK419j+xNVb5gPlv5H/JselD6OtVqoHkef6IDdthZteuslcN7imb
uPXK6q5wEC0sDPkJpWYe9W5lzW1iHX7YpzYX7mBdxJzI5xEJwyMoEC45l+Ww2495
gUXIhsngpRLNCIE54/LlIDBgvWrjq6k/S19sLpr+Lwd28bgdoPvcSHRdZq17OJx3
3bAgyrzClLzCA6NcEfTftQJEMEI1XVDt5yQ/nw90L4PTuZAWF9OGMur0+h0NUKI2
iVDB5fMaitS9Ktjo6ZI/PYFEXZjNb3iWPHBZNt6UjCYzW/Wl19w1itvNwuB8dK+0
atOJ5M8kA6uHZOAbhawSVG1NzysMQare47LbD2H01a3sZBuUMwFIvuqJNwIj8HOL
jnUtj3x89p2ADg4wUwsqBC6IiNL1hEcDM/PGGTqA/l5exhCFkDA7Kkr25XIfZbUT
uYa0NKMgOxjX0BE3ADN17uSnJbS/bq+HaqbKn56BB/XnmZO1Ukos3tsYhlEGMBK2
j801jJbkzfV/hxFxtpYvn2wJ4SsInB2PY2zoa2gkUTMj4vMk5Y7mV9uwwxqlUgx7
osoxeUcvtqLp2OAh9m/4n8N6JEokPAFnMsAbJ3AbCmdhZJHEccJIyfxjvYOS2vdj
UB2HW2X/efpdn6ikiccTb+Kb05NgsLs4SNyOy/djiGPTAoQGAXj4X8SfyHtK3x2X
r/iCiJpNiqYWzIQUVDLPZqI78B1qFlkTRussugHBWDVTfG1J3uumvnRhIhrj79Og
GbGdlyZ2PDvXvw/8OGrl9JqKkI/5VBpcGiY9mZJGjEe9Kl1NAlT9k3L4sdwBH+Lv
nuIaSdl83uFlOKutDAXf3iLWXJaAu5/KBR4DOzZ0qmRLf8f7mq5sy3O5kWKl8Fr+
94Dv3I6b021wVdxekPJU9zfPXdyniRhaghaCrKoajXye5oIcSmNjPWbsBUfqsTX0
SxGqTTcVzB6U6dEO+aXQvGfaBNzfLCmBmtnJTqA/hpkizpmqSW5wX8hjgYZr4F5Z
2Z9dqmZR8WpdI1fp5xj59q6EITb5lKhF0ftHk5XXB6jdJGGhHb0/mR13ufihaOTx
0sNdVRIXxE0X9DmrZH/d4CRWFCDj59WJtAPsAdGTSyjg8NcbvXmgjhY0wduoE34V
zE7W00CvGeS5BpDzSyipH8EAnBUFJTPsqIWxRBgKOZsLKpWRCzG33SuFBTwJCVmL
6RcUyJp34N9R1Y0jeIN6SV5UKgFrLvn/WTUIBb0NJcvCzJ930YVoCZK3cR/gUahO
T4hOkywW5/hqPivg9+Byetbk3i20Y8rhE+JIbQh+H/0B/yHrSpFjm/MqbNTQqcQW
at+xfVdFjTmOY1zZdL8SKjr3eGDYfDro5kMm3ywFFx7ZxwZwZZYbjuY3vZflr+iI
GXhPAybp3a7KG1eZa3rNVUvI6bthwydtR41eX0rBmpfGNk6sTfDKQx7TZVnK8cpj
/bWPbU0Gy6xXmNuHeD3sGHLt2HEqWX8HjDz+VKyHUZi/lVi4J7MOJdZKvRc2koKy
ttCP+KKEsdzPmS67RlmrurZkYKnsjmO6Bu1BoS8wH75ANwCl+/AnlcJiY1WWn2fd
HSbk6cRLFy3wNZyg5BD3nE1jK7jLb9XNr3++1tRSLg6E+1WGLKsI3s50boDg7tfk
mhLhfA8nB6bY79Fh6rUNyvX2J8z/itHTD/LepHUM8kZmwYderETEOfzde++h8jF/
/PDkzlf/oalYr0wlhq4WbOWCz0rIzk4SQEjD0bDkiXd2eKrpk2blu3sm0DOGRCF6
Xg3wiKgeeBntD3LhdyoM9hkerdxQ4uOrkvGYzke4sw6O8UFzQExsHaNHsR0T7xe2
uXpRxrrCAIouMvhKKAEhenpEpUO6pbzqui4h/F5jVGfgwNRCoaMjKPcQfI4oUqga
DVDm9Kxc46uXx11F39CJ5rnvF7/lZ3L/IqMBv8ejmJ9GNJ8WPzmsuA+vDkhFppZU
R/P3hzr/d+3GfZ6DDgYf6BVcMVDzy/7C+CddomUguLopFS5Z8LMLhC6MvRTKWATx
OsUahBCDH1tXZrw4Jr/vDnolKe4Mm6LKDKfH4/DhE8jUNFUoKtAA3U5nLbNl5cYL
0BcI7TGX/ziKhyqjaHsugzem4WffmA5CvC4d2czndV+4PbRVgH7wSUdnYwlSNXG4
2G+zx8uQycXv4aziekAMjF2+ywKeTOmlQeJnj9TJSiAZsLpaMANBKJNOxQKoi6mE
u0WEqR+ZlOeeKaKprrUnFs7okB/lqpHZ87n5VKbQeS2hh6qSKgV+7zdhWC8HvJfp
t8Jj/v78TWAVFKglhJolPtnxO0tH1kUj2K+X7NA2Phjhfk7Fz/DhugZb5BQMZyel
Q/vK7fRsr45TscTbs1wyJWTlAKBiwyHTb+tRQTK0VNEfIiFysZo8VlodkTkHfeOz
Qd4UFm1toTJTRZT3eFMymICiRP+q8lxGt9Ta37yC8FQqVmd8/uDCtiY3sZJbDQFU
T+JNKEtvkkQ2Lk7lLWaTNYdim+ASAbWxnyPT510ro1K0QP+swErt0ypXdvwJlsAi
G/9WWhOh0Wl+kPJ02q5VOBqxUK/s87WuN4CMZz0dICUqh2TVCWZDdNi2bOfd1URZ
CHSqa8FgwW8qy2dUIfi9ij934ioEJZ5aLlsgB3rjla6j/hiTtOZ1MoF8qVMAEDIx
n/MaupinbgUMN6kXJYQdA35lma1jHngLipgcE22ljvkhZ8mmuUadQAFFoJf4QBxW
DG0g4aK6xTK9rDPWpYLS7qcX2w4Gswn3h5R3GgrV1BgmRSox/2Hhx75Fweu5SS6A
LmRlUy8cZ/C259RxHHUNlch5XupFQQxIuYtL+5X8eNeA/eTiLyA86GImTSPdhLY0
VLwJVk9wlDXYDX4kJzYRites2W0YUn9aLOF0dK4UOwOw1dTzuD87qGub1U+j+vU8
HtGTvYhUxiLtfNCmVz3UFLF50sVLe3QTaFY8JlAHz5lWCCMiRIn7a+Hes1Dn13Kt
RVi9h64g6xw6QviA1tiFtnSdz91zjiAcso+tvjAkbk6Ql2DWCsdsvzKMkj9kd5Xt
YFBTAIwZE3XXnrywmTIuHGsxPO1Pu/6AqQ3HWt39hxTSGgYjM/pE7tqb4C1hSwJH
D+JDitGqEdS2ExfTsxnK44Aqyj0TpubkSsbi1IorLrGZ83Rv5BCFblF9GqRomtBg
QwtowEaEtWvBDkzNDAH4xFb/lS59BNlGt5hub0aJVvunTVPzJBp1/N7hAFbjvdO1
3IzeibnAIFncoC1XwE8PPDBcClqLBFvKMDssdjWTZpg/y3ccEod83P0AaIRffPPZ
s17zhQBHm02by+iw5zL6MvE2D/4IdjecALaqMBZJnCOJNbc0cIH7c9l1/j1B+0A9
fgYtUPlauJVc+BRgDvWDfZM+mF0g4BBaZJfJfQWW1KehFx733CbTChx2NKnOFaC0
fXPQM0zFDoGkZzo90oQKmlO+BQ1kaQJ2+fURpNjFnRSrt3p8wLju1VIotFEhtRwb
ZTljuC64RLkxeW+/q9nIKSI2s7VpC3V+tdJmsTM/k/iWkoCbbECVlqJW/4SSLINv
H43OO/BbQluBGHocZnyk9miOh4quh8rlW7UKiZSJHjab8rz8SKvoR2U1gAfaPb6d
EZubNyOyJNY0SHhJtkmPwkMuUnVwmg3xNZJe0MijKwPRMD13m4wK0Dz++KPNxw7h
qY1/JmDDGGIvy5MQDS1Z5NKordOS+3PeDsguCnl6z5Z9ZHAK9bh3yh2bswu+FurZ
mkN4ikpyrFLxpeOa8kF/0kabq4t7xLe5H3EBIID1mzXQFNVoek2FBlfWQvwL96xx
A9VSpGssq7Fn03aTMqPBxEr1R7sDTxuEd2NBI9CeCPqTN3z8SPjcFtRlC9VxfxUq
HvQkaFOOzxdPKbq/ddmFidt07mpIfVLyL53xXEVRKmF6o3YcRpfRdm2yUUGWe/Wg
D+tCAJuopWtOPmLcXmCkkKWz+0hpsle03KOfeM5u2cyqax/N1SAb1TyhfhEI9Ei/
IeFcskji+fAFlo/RM4IfDGWrqveNEuFirZ/5jL7f5QX4d+hXl3MrcmHMD1yBmfiG
HrBPXN2CHzIdKBMuqaWAe+0pYVjVNgN1kEWC4k9GTzigRhDAiwzsV8ChPgxUYuwB
d0ks75HOclgknuubKqWapzRZj00vjjtLb/T0RYeTnPaGnvFJzJgoLb+cUXnbCfjq
pK67PJU833EVyeGYzZm3AMwJ+mt7rVHvkkemQNTh7vSOp4V50pjlm38eK1vgF6TK
5usR0O+aApQT46AXrdsRn5QAvtghguQowMk4wLqnxBtGEsVP3UXrAoHCbIWEKHWY
iYrjGKaki4IKeYS9wICQPiIN7ssenDgLSzvFSy4VGoLRXGYx2TojOFamu+2hTJ0b
fr/W2Hj+fE10kRxdMHPZ8BYu4qLgDqK1E+8oNWlzkAgHPTNmpDdT3RP+RnCKWGmy
n30BqdL0++h2lIbDiUIYIw9ahKkjjWjtqx9bTOdj9plTRGEALM3EqwfYSLBBVIax
YqyvvKqpuoK6yNcH4hVH22EG++9dhmxLgXpgWg/odWa02M2gc+wgaJ5ETsH2Dgux
aLkBIuIjKpbX+LXuz8roHo7kCQpM9bx4bvs70IY7NcXjZMX7NC09kKzUrvRPY0uV
W1pQ3ERzbsKM9lh6JdHMo5cG/kJLNwaWfqP9GBOhHsCUJdoPOBZ5QEjx38R3u4Fe
pA48qyCdHAXh3Eldr/guTsGp2YGpdHv1kqcSkEuTTdGzE5FdZdhNsko78seJzyzs
micbVfX2qQBNI8ToFGXeqKzPVG2i07VHBTBN3YRW+ayHRl9lXmgn1z45xVMzC1/M
CCr1GCr1U+HyiH2SdbdPQUTwhi+gJWnsjt8/UN1dBB532HolYql2xRZRWRIY7jI+
i0jyTw6SI/zGbXtEjQA642XFgKkAZKdLjjJq66NQmLEVK/sDGb8F6jQcizCn5I+k
ex0t4szJ+yezXS2g/0yQWDUL0gUXDQffKEJvHomgGUoySxOZbSgEIQIZ8WL6bYX+
PjNxKjVWOaHk0bpd2KZ7eyNo23moZTAu0glRwTj243jj5D4urfyS7Y+8f6wFOa7F
GFX7/sivkzc2zHVf6RMJMBSv3hWgTzeKg5BUff7Nzwz1h0H1q+Qe13FxxkTzWNqj
f2cNrJ8VOrpzcDYl804DRIsmXgaBOCSjM4EEqBwsvaS6+euSld7B/TKxIlZChsvI
XTD0/YL8mxRiMlK4AmRcSB3WE+T1kVgeeB98vPULbwQ68lwVNfrJKYjR9BxicfMp
zG3iKrsBfpr6IPVUvHI+cp/GObhv4ZUDus5DkXC30MBdw4EIua7KPRIp0fCEWm7a
MofX3awWZukdkdjWi61FrLibsQRwt6MS9lHDkcYI4WGB3/Uep//pZgZxr6tLWeoE
eIp/okCx5e5iGCQoY5chqaEeFYcTZNBIjAUubA8ZAE41POj8xDSfxdqld/7Z2Qld
uLGlU/zkiKBpU3ssx7N/mrYqPi+Op0qFziDeDjSHZBYZ8k1mUqi1DjoLwTJSGIPp
SY9GXfd4jJXtKoqg8M+dRdhS0aOR7PIO4I268nXjYsql2ZB5YQhLlwDl7E6aAfZS
ZsMuQOx0FA8fcX8KzOUSq8mPkXZJvoiSHHcu5UXpTJv6DIv9h05M670n2E5TeePz
g3tchDYlgvvNzD3WOC/khqet7laERrvYFzH3K0ysQ9+RD4niCZy3OlTs21o93GWJ
HYRQmz/cDZezENBnymffT1LZpz4WLN4RvieYaJ8zs6ihrkaQu0DnXtMwaqf17xDF
KC6y3EloMFf8s/OsukqEROnmLt7t0kyuBtQeFhCwtCaHPwbwNVnLwFcNaB6s/wsQ
`protect END_PROTECTED
