`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dpMQVWiG/U6Mm6WNU/L/y+KRvXXgxucMeUMIj6GCEEjpieKWRO1HCC427HdtoWDT
hWVw8aa5jsitd/pMdHLpHYkA/p3fcXAieOdpYDA0Vs3ApKVDCz4TeQCl6a/TrlCa
8pRHDqyEfRKQH/QCf4xnyGUjANJm7YnfNWI3xJbwht/azDSO7qz1YjL6rua/9LoE
KM5NNQ6ecnyd4xuca6CFQVGqNaHoboMuTWJ0RLt2glATz4Kxl42T+OaU2OwjLcjL
nj9N5kkh+DSXi9R7UvQitjR+Uyj8+GhXWxrioHSXFtM+U6yiUCAuF6I4ZMp2ylOV
XccYKuC77ExgZBK2lfB9R80tNMdURu/ouk78mcnpLbrswRsuCQjXjayoZ6bAbLlF
KuMC2vZF5TmP+BrOEf4LBxf9GgsQBbEPbE2Ms3fW1dLQYXUcPk6yu1agldmz87P6
obrtCtZfWcpHGSaE5TEmSHJVfUdRGtV76HVYdsFgTpW1ftlb0LzSPOFJf4NayK3p
O9iqJMpSsNPlJTnhb8jnXh+JlhB7dW7MrhabxWcxFKWsKxw41i5YWgymnMpVz4Pi
tF158T3+pETJKC+xDVeMh3+C70RG3T99R4LfuBfNbYHukk+eJ0auxzWgsdquwW/6
zBRYTAzyTYV3QKI78d6pbS0PGW3B0DxMQLoIexGEAAxNgiBw4OYj5fpjNzEvrh2W
+buK9PcJM4J3DucMBZ1fgfOZWK9ae9mWi7+Vl8sK/Jebq/9nYAH5n7068nu3utPD
J88KD3A+QFPJgIEmLYxdAjHRKiTkXFDKEToNzGVPVYXkKArMNikkZ5P9H/h1q/yC
JYtsTnnMDF2j9vb7rqOua9PhA+F/JDcOUXd07otiH9kCbP0CIZ5VSomFTFCHvlUW
JPnKttt6WAvo7blLPKIS45l4ME3rx6bFKPs3MD8bfDANxb3b79Fq9xR+LNvYwIjk
LbrdW836nJbTWEwAq6jhkBeteLf9qrtC57eVCjyRwHwwHwTh2rjHm5FjKQLCJsPy
OLMW0iRHxu1MJUg/lf1Ub/WBwNVabIjY2nX0qJNkDvFgcN7va0CBpR1KUf2fGi9n
9IcYyv+bj+EHlZ11jksEkwGjoBeeSRieKdtX9BM3xnwdZ5+E1XebvxhDEnAvfnbC
y5zfSxhhanBVX7kfpBZn5lj5+rJPV6gWUOTH0mJmt77iMHrec7JDeIyNZUWUza43
11+OMx3/EQD4hNcjt6hI8gwTYH25eYisohLTF8pCW0ZNPcl1rJbuECJSuLEqAVtI
A0kkpv0C0vW03fW3yOSE0e6pGPuKgcctsAc51Pycz1LZ28cx3KgKDGI/dDV2KEnx
OpfqEyb2KA62nGIYtbXH9HklknMpYIIPLqrBTyANy2ca+AoJqvm71nafXH7F35Db
/u0EYG77cxguLGGtA17twm5NYhshQe9xf+oO8GE9U/jj0sRL4nbehrKAIbRN8Pwg
ZzeyJehzvADodlTXGIpCuAxOW12huEMXO4rv5sZxV7Ij6zrOEonbl0wduNeZxjV3
rUfQC/6KTLPvAOQKjS1M/F+BW9egUzybcioDduI+Zd1FM6cFenKT6ky3ZyH3jB4Y
8QiJzDAnvftO88+wHgAN/t0yltw9tby3e5xfVIgaRc8pi+FTpL160HnZGizfXA6Q
mMv8gEf+d0rvZ8dVWOIbZxgPLHe6AWEDtbQd6ej1TmLmR05UBkMCKaL9tksiiDBC
t2pkIxunwIPBIA0N/pXKmICH1uANg9ukb2WISBq/spmpS/97e+kjxlMO5EX+MnIo
AbRB9+YeKqwrCSlK6If33R77+JanxZ5RfQZiwV8nkK/zHTXcFMJp6Fx4UkTSUk3f
Yjn6EAlOaq2jEgF49ikEkZVDVwKPDdMGu0P+NzvM2xBhCCyFdaBU9RTdmKLzKTiC
jijz62k9g+DD9vwt9n7TNiR9O16kH/AHarqVK2igqz99f1mR192BnESSKQjZI2Ud
45Du4y9XEpBQiLDZwD1n1KJxa1KZcOhNmD/Q6pxNCKODLGiy7llBAESh7kYmiTSE
3D91ItNXME/d8Dm1anthnV3hOxQzloGyX/iz0TAaAhc6sJreM/EF4UgKXxdF1zoK
yo6Myfs1+Dt++MeKEIWMtcyv5BlaX5iLcvakvWy0vSLcj8I3+SIEVNUQ9BQCqVli
6zEdntyhcG/95FPk2TsRKKFXwSRx3Jc0VzpVxABRo4mKQRQoBZX0xcjzSUrv8Xw6
A1qfumS3EatNEqpttlpRyjd4oNY7QJvIxTMODay7AF80jT8pJeFq6AbHxVygHJjm
tue5HwmwqYfvYbZqj0yuByVRO2qvbiBA4XoV7dZEFye1BL6FiKUvrd9obyByFi/O
1JJ0AFhLwnYuApTFy7w2lffPXmqfr7injd/9H8zbOyWN2VCJLkNLRdadyzO89l34
vfHDY93Gg0XIFl1GDSUOwWhNU/qi6RSGdkWdztYymEu3lAxMcTW/IuyHBo/WKRsF
cf5Il0VlcSHVTndK37Wr4H9pSek6H/fxq3fljX9nJzyNGYwTsQCu8tN9XlCO/aCV
LaCz7w88IKvNEGbYFXtSlfZCMpKZDeLgwlbbkoATCOhg6bCjegsPnotBc9zNTO/i
mEwjcjKG1qHVrg2fMVUGLjfwj6YpuiPLFDR+qIjQ6cuDkSz8prX9JntFxdXjj2Mo
5y4SpbGuVNYUWOpr6z5dO1eaU658uoF04H2am/1VMvpl5xpWQ/eKBcSSi0biAnOi
x5WZJfL3WI1KX+Jg5pQ0lHp4Eg/ihMselJFho+tX7447+c4W2xlzKLqHFjIVi0bz
6JMQp2sLjuuS6uxVgRFlV0M3Di+mdiAHYZ5cQXcIxVWUecEsvHsd8uQ4ggRM0cbJ
mF17h2eCbJpAkmV+lp2mGh6A/M+my3N6b6RaeZ8KPRMCbMsq6aoBlz8lZkXcYxUd
++D5p/8E7r8y6RqarjDCwBYn5LXwK0NX991x+wTsuSpS/E6WL4orPkxHkjI+SrLy
KBAVekAs/SjL14IVO6R2uCftgbmtuPAMZi/egGmnVpwb8TFWp4NKG7HuMTf7DdZZ
L5n61aCt4kNPJ17mOxl1/1z4o1vzk4p3nsqDBIXYuUIjyg4C+dEjCWuLmp5dPyI7
X/nF29Qsmebe6EKeFiomEpeSKSBHDCJekDpp8cXpA4DXYHAUeAtflHEHjqzl4DLO
HzqQ9GFHigVjvkF84To5rDu9FiljRuUqpQdCSQD1qUvMQgiACrlE3uiKkO6DNR2h
ZZhn6jaHP9/7F7s44UkZ9XUvbsCOPXnRZTG2m0gGnvfQnxsAiMZUFR9TQ/VevfX3
jOcRcMA8oJarpc05s3KvS1Lvqoye6vQxjRMH/OQzphDBSVANmvFKJO6BR54lItiY
evK4/GI4BvGRbd19qQruFzDMCITq0/GiDkejmSEZuj2jgR8BQ5N9Nrew+6UNSjDL
fVb4rlT2zZwIS+lMwkWy/rw8wHnabzeXWQYM6VRr1MwSSPnpxTTAq+F6v690G/qo
zl9UNCG/VQ5tvb4L0GsnISg6RPdLJ0F+K+wsWGzYqq98uauXhaSyy+dm/B9AZa41
iZdyvQpyupkXQ41Upem6fC38lI1RZ9q4knDf2Gk/dTHKvvOZcfEF3/lOt2WlxJRN
NK+L1HLNp/hkZUwYLC/hGxI4eYk5kRF4MsThsZv2XIetxXgVDj4nRBVzdvRHMu19
dLBzoSDDXe60w8dLsJwGaKyhwIIik1B08KJkf4DWFH0y/hA309etuAXIV2IKfENp
HymQOEoFdtc+g3i5Kt2iWxw7hKuuhGEjbdBiGSlJ2S/o7Pf17OseX/yOd1bAbifh
2oXeu3P3K7SmD3W5xJqO1OonfyiHbkPhCM9CpzqTf0Q=
`protect END_PROTECTED
