`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h8R7/wGR9TVafmNQMwIeeUQSJMUFd8YsAidiiPKvCD48PFLzLZqBLc055rprCsQm
+CZcSLHXPtkjHYqaqoR8i+lQdVL8TY8WDQw2YO5Jtj2WnXqeXK/GKX+T/1ZT2yiF
ksGJO28Hf/GLJx85qOA+YnjbBYA3k+8PVlpeL7aKhOCfl2vUaiCCnCr30fMgydAv
fnajeexFyElhuHq9igiAPZe4Z+/NSzMEQVAGtgy9dF03vtFxE+VoC+o/PSSFxbgh
UPf+qF7orQUjYE89mZCIBid1JnQv0nAGfzgtZr/Be62ftfCuhlAuPFFNcfnYG2Ei
cB2y9aKJlb4xSLs3ez33zhie54rDLZpGHbbcPHS4V4qEb6ce7MMA0jGpyimMTaBz
VCWwkmRgw39bO/4xvHoyP+sgV5hAFMNJiw7L14Sq3BdhzxNMNsm67j5hGM1AJaoA
NtXeOnW4BxZaXkN1bIUC0XRatOIxD+fME6v6ap3mf5VX/rHPI7I8aNUyxVCPu/TK
fBRzJNbQHap37rAZsOLyRlFj5pWjMeBsCl8fBNWwOC+0wUMtadxcKM0FTmJh3aYd
QVftZLBa5ZbtYUC4Dn9Gk58o4NIKr3s1/tlDfLALQKaXxlkINY9pijRuB7QdlqF0
jVEQqge7DYxb6U5KJbuIBv38zBWuZ1wn2xUrSvZ6wj5hVn/N7rq3xpuHdr3Q0tAD
`protect END_PROTECTED
