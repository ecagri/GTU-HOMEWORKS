`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/JImx4HfxbBVcXj23IG1wywIHjJjsUqeRWJsh/EWKmS+jNojVVYWFk8UtWzpHtaz
H2kyWZO3vR247KbNBgnKZnCBYOlmK+xy+TdhaQ9tMDQiwR6KM9J0aUJHXeiQiW9x
tofoKvhyJOYf3Sm8SIulbbsHuAjPrEx6l/uqJ6/EVLvGnejgWWV4n81Tb/qgw9A1
DZL7vlt4UuoWSiobhisgWGqRgJQXY7fG5iC03yswGirPQ57NbR7DTpngcBr13mdV
5ztCjyrAszpgGB76+GR9bsSyzUOgWdNklwCJNKnTdVA2RxbMgVRtYwuLIUkJAReD
U1qccsK02JSTB+b01T8W9PPum+2uD9q7e64BUVQpvf0/DDQWhhhUG/4actnuWy59
lIkDMVNzItr8d5sTsYEgRHOw7hqxUZO0dNMDi3xfahufVZI4G9uMBeY/q5Hqaxd4
JPzxfZMXCcNjm8CBmLyOy9AbUDdm+UFsPWDjifa75+FKvxe+kwj1WdrkwZBu8Y2u
ZQpyDOPBHI5b5CP0J0vuqG4rbsAmCPvlWBuTSK2FvZ7d0fBpIZITmTdosftDxKgA
WrMqKHRJHC6k2IicL9L5y7lqET9t3lgFMGdMR22XKLkxrBRRKFGpa4aJiaauP6r6
WuNee7R7WLr4HOnWafeTJl5BrQYLbe70eugdDvKtGFR/vIkcnNGSdSCebZAg7a1G
i8zFEVnFXwqoQ3k1iuJZoauvzk5lxGYoOzyyQn0P9DZyaYec+tWQ/Ra5uiejJZhu
pe72HDoacFGZl+RvML6Ptb1ZGMfaegDtDZ3XyPoET1C3r/uq0H2oqWNuGXXbGCE1
Mn6/yaags3hM950B4ZaQkj+nQXKQ1V4v15ZfoB91odlMVNoXCGRBJ7jU8W0qjKF/
vw/VkRP0+oeBnXWvq+R9i3B9vaSPBXA0KVNkyEMqmn8+wudm1CBWRlysscXpX8BT
TXC9noJdyZ0o5uUsTy5QP1KrvpA0juLL6AWal4EZORaT7wBO1Q1GsCVewFX93kxl
HDY8PkoYeBOTycnOujSnmh7ci3xvLAoY/fTqwzOgRvkTIdti9T4Mgl/vxebrXvnf
dAfV1DlRh5+jeaiaSrhDdBTLn34CzwdxXUXrIDyR/JIUBrmQJLtAW7zx7qnWX5CX
/IBsVDd0HPU6+L49Lo96ZXvViVmo332aFT0v4prFR0h4YuitoRs7VoB4i87fX3td
Nq/WuGiQvSb8mYEvKuwcWYk0Vl6Cs+PGNmcgsR028NelsGbb27HkHj30bxFzeLNF
m1vdAUGJeGGrC+K/Nn0gGS1EJ41QITbJvZyUUAiz1RaIOcKmxTat+Ygn3E10efE4
EWE1Jnjk8cEPL7DHO2rpMCgt/xpWEtMkqijaBfgNiEXpVSTxZVgu2hNeUPg/awZa
TF6MPhn0veXb0RSIK7jmJmsb90OPDrVKScudKhHxVj2cvjghoTTIRtNJGbOeDU6j
nXmx0my5x+lxuU/NxzlGqtEY2bFhIp2eK6DcM9jKjBKiyv4UnSBmuwJ3mw6x7LHW
su73vGQPTg+zAdhS3a4tKccfxP9/AJO+QvFO+nbN2Me/zFCAD6S/gLq0R7zvEsfJ
FHJrPauH1mZZ0EuaKZsAg88IK3fBatdZ3JZpCqR08sFt8UAX96ipU1v2jDm+pPZA
D7uUl/0A7n1u6JqJx54UtA==
`protect END_PROTECTED
