`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5n5kKSM8Xawu/W656EmFi//vstDG8JDdmduAtY4/i3DHt9xx5Oyq7Y/aVajgYiCc
whamhV3rMzeyWBzNQT0IYyYDqKpUnh6TWgeEGEp+lAJDsyjPoJaRntMOCMDrSpL4
Dq1FUDF5iUOiiUv5VYLHCBQjYOW42+jK6vr9CPjinEGjjouKypdcDhtwEMlNadtn
`protect END_PROTECTED
