`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3vPV9HFg99LX2D0q4U3EuaZRU/b5XIbnFWckw3x51P0wkzEAlJSWDGNmnd6VfZRv
usoA+5RB/hXZJVH5OTI4ASb9Kss/ugUzSHx8YYXcThkzQzrAi1ibE0eT2UVM7v+y
stekzQCIuiqvxHYFU4rh2z9MQJvbx7z0DFxQmEIdT0akbquNbqoOyeS8DFIM+tId
q7XE6bNBaqXenU3CNqJcsmvoJEWAX2daVAESOD+22zCEYMfPnGu19yFMRpN1/wy+
Npw8+fOsyHnG0Mf9yF9sLTLkPtA94Nkg+5waJkJt1hf7aX+94iLwbHqDT+Tf04j1
0An46z7crugLQpbPB+DrDptDguYBYVgSPodrA0v7yQO9f3kCyDqd4bHJAkh4057E
60eQIgcUKrwRtXp9VS2OwIEmFBDFOH/Qz+mYNDh1nTPeISian2Up0ZI5GV5V3dd/
25r8V6XozDCVt8Ge3cAHWlU8TYtVo39n3UWdKbjdkb12xjf9y4+pMakmk0gi9Ylf
f++IMSlNd61fr/0OfofaYDNaiPbah4TtNTAnOuwmqx08fHYaMBa75Z+1Tg5v8TO/
2L030vn94ymiDRDqB7Ho2deVPnjSlA8IM2VQGSysR3hlE4xtlcyp7kEO0QdcwsRj
2u3sKz8H8YLEEySGD+z78riz+DfHw5smvaGv69AJzdAE4PF29rpY2581imfqCmbi
wfkCo7d6WIF1tkkgpOwI3n7+CmRL1PMYa7b8GAtFE3pCxKOTRQYALEB1JLnqvMHN
WEZDnaE3rNL37ODqJI4pwZcAFZvWUHGdD4Y7i/7Z+dd/4rPHqP1UQZpVK2OvhZLv
nmzJdnxKncHtYS3Exk6doOYQ5REiJXA9EHmN4HU2R0TFwlhkVabumjlCpkz0I0Qt
AY1rlqo5ZuQA15yDvyilFqfHwcs+lrMPdJ081+mdxOH83CnhyIbvbBMz1LVGrmHB
`protect END_PROTECTED
