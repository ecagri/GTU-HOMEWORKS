`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VCitYkNJFKHsqsJgBSYTEjiUn9KSD96JQmcM0rbr+SkO3v36VI1zFGTetn+XOo8F
EksJEQImGku9PEGio9K8OKlkPA0bM2dNVOBzCybRlYSNOz8alIdXlfQyTrsCefDs
lnrwsZxAF9tu4HsNw2ABKEpjXkL6b04Vy2LP9aUE483Xl7ntLwciFJEwQXplVzPG
fw9VasgiT8PMbqoO286hj1gUoKiAAq2lapHZoF6btAGYXRNl2mrK+XMjxE0uSsYr
relprm+deXn+Pfgm3GcALYdMungVtX4CA56y1xnVRlGf1ejTiAo2DI7FFCGqmdin
wSoQ9TVIInw3oCn4mBB0FlMLibfeufX74+cK+bqrrfkpBafZaVqkHEzM7iAjDSSe
Y8VnmfBdm2PtSWaZ00k2Zey6xn8IPpQh7bLOlGzDKcn2OGm3lhwgR1fBsHuuqidY
W+I1Kst0Q2KqPSi29c9G88AQYyriUK1qLB0TmYdaD0+uRojJ1g/c7erERpwZlFCE
EobtFHWydtxneyfWQhBC/sZYZPOdWdg2DTOgh7HxHizSWvaohnegXS3yhMEJTpZ6
XkHjPJcQK1xoL1JwoyzDbDaDGmW+eTagGGI7DYZi6+w5G8bWCcEKy8HssuAdrGEb
ZfVKznYCkJ2enT6AOm2sR1LteW5IgoazdtyidJKYZY5F62hWC4W/aA96tYRZFAMG
Gr7o3GwjkWcgP5S4JJJY2MOkeO0RDI9fCnI6IUqj3LUJ2eiFDBiuZ+x+cz9VM/Px
F7hCtyo8FQjPuu0CtoTWTixNybb9qID5ukZoNBWUB9r60k5YpiZvXDeV+G4z29Gk
iSN3q3K2x7FpMcfTI7SY9oj+hiPUrE3lH3PvYsZlH91ml5wA62qqntcBuf+gszA9
E6iR5+V0zSr6mLTghfODK5dHbvfMLRwMaxhdCtHHtugaKBs2xCg0ob4EVAdCHSQ3
4Xq0v/tJt+eya8jq743YI+cmKGGWgCi/UOepFlElDcd2aNFzz73fWiS1+/49uE8I
yRxHHd2Vq3fwcsVYxWReDRmzy6v1WcrRnZ1sEPSOp8tOeO1mlo5n43QxqGndDRHY
YenD2r9CqJb1dwLqDRD/NMswlSCgQ6DWjtbRHfVF9xhDrdL2//J+qMIexemg0Byr
6vJicRXYtlJk3zE4aaQavoyDfqa2v2+AVVc/xWNtuaJKvb35RjuKjW3BWMMqieE7
IRrW2vHfPGwTW9cxY5W6pvNlw9T+a07tlL41YRr/+UE=
`protect END_PROTECTED
