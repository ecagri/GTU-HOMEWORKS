`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IHD3A31SgT5Vz0gJVpEeAXVVKivTZFaL3S51ar7cx8U4Uh4qmGWsIFoyqXswi0Wz
Jms2vVYQ2+BuPI3YkYal7rFjK+3yV8+K3aP69Mo7Yn/ZKF9A5pjtVSdDVeoolJi8
KdAFQxB10poFiJklkFpXyoVFu24RpmLMplG36O1HkIZWhKTl1f74MPlERtQ2TrSy
o9kJUVeDpzgj/cXUzGo4CNXqYhO+SA024eAFTTKFAH5pzcVOSr82tgjkVC0GJJOz
RxTU6DFmmU2kYkRZWsQYNW7Qsce00b092cP2lSsJNkzmeOjkH+m8FvKgJ0OnLj36
z299/IMXEYdl/+VI40Fb37ia7D+hTpI7pEQQVbF9Z+RYYLm3Q0sCEuTrdcorSYyF
jTAVlA5E6jHb+8DiYLw66OCkPkELLEcfjdcaEsX/YFV91bBIgd59b1PmgqyfICiK
ssAs/Read6BR0fQV9pMcKAWKO6aHr7C8zq96tcT3cA/xeuIthw9jRQd/TdcVT2JN
nN1LuLNT5nFgIfC9GMgd3cd22bgI9nPSF2o5vqyKUdO4Nyi51q0xLROLIZN//kC1
pAOwbu9s9U16c5k1X5JhALPKnV0U1820BS9UhrMOchDChMekqXQKm0sfJyhkXPMF
nCGPXLtgK9tBrDZvoNie08mIh1e+mNLO/YP7vJ8c8ThwZ9dfFjVwIubo7qW+cdww
2/3mi40aBx/aXZ2sg9ma6W3YEDRv/xMmPvj1oKn7D4A9pnQABOxsZ6UG32rleEsA
fqh/OYAK+AY3GG3RVIvmUv7tC2WqvCmg74XecS3tXEahwWLnSsEZsi+ChixHuoO5
eyzDKmH3e3mpyBIgJQrLJpy932+2vOlGe6J/1gwhVTHa3hg5LR5V6OC6E9AeyMGx
GVJ6YQ2MvBKz4+oLGqfd5+aCy4r6zBctgsXtWvqeFkN+DNwqcRiwwuC/gHlhuCze
`protect END_PROTECTED
