`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7TxhYvI3ODI+5MbXL0abt36d18LGq1JUn7ZgC4lzN3Y32AAK0Yt7B4CDb3x0mnms
ObuVFo4hFBVAwk0o5JklNCf04/m4w5qkZkwEpppa0Bb18pqFRXp5ebe6nSAO2EVr
JiVHQoKOZZSaTS1HgDttljGWeCF/F3dKNixDmjTy0+29g2fewG3khlUdSM2DGquQ
Tb6oNL7udvPNc7oHZIAExnBY6dBENe2r8LeRK0OkAhcuAWG1nidd7bWLneXdWvnu
mtHBt38g8o7VrDmFOOXGmaGVIMqx/jOJqPKM0CVyiHqLG1byE8rFQPOZY/QJeOLQ
14XyL9Ao2LcXI+5vqKeKx+caRKBrzhWpEuB/pF+K/+G4B+uzzsmrNR1trYqxedIR
LDC8qucJZpWfKXVb1BuEMxaLWtLoQ/q/6dCBUo+qgak7G+OHYU+j0fZABOhhgHYI
I2FHmHIYuukyFzzx8sWr03q6sfenDQsQ1f4K6QxQwBl7rR0GEyDgydxpwzI7r6gW
B2DJhtVGVOQj+zYNEDvVy/vZZoQo6SMXUYWwvpWwR6LlHB+z/q2hRaqXY0x0sm5l
RfKDActRmmrGP63e7KuyjvW8Hv4HezPWf4pOtWgArDYiiPphWsVa/C+XTNUP9fMK
pG+uwycGgnfGTSQU/qgbD31OUq+u8RtFT3HGjy8Nznew+lLNFqXbX9YDAwTWmoqm
ZD6umkgmG9PjWQhusA/DaZBjJ5TTSosetcIUJsUtymOmQOvsvtdX+bz7fF0T8GzE
WOI2lhIi5hNtap7jghy0S3baUXG+mjQiHn/vx/B9kMApWxy45te5zOColkih9JM4
ASSIJS3dfF9W/jXjRBXxMrnCRJ1aKLFlGlP0p5JaJTnyMBeYhliRRuKoQqJ75E4n
N3FyO56UbL4BZTMhCwojazk579nrRCZ8vsAlqFvJLrV7p65CrkBDQR9hI+bAV1KJ
sJY4zkkwsjH8/8bzmokT8WP5hT7LAh9JIBic8M1hzRPRvX+U/MRI2EW2woxCfdF1
WrZQEoz2J0vJtCW5dgye/lNUfErReI7G7LENCNfeqP2JQ0va0WJIjMJEOY4kV5WG
bYnG1b1pzKpIAz0ebHZTrckjl0mrqLrFDVWdZiD23HmelbhLiudUYyjQgIGjNB0S
QmzKpsnY7h+hOg1sWcKqLPMZOjJofh26/wbU0hsga7qeB84ApE6aSRVWWncoF3GQ
uQShKG1gkQk/xGdO7hoqekjp6s6FnXi5FAukiksnHa9Rp74ng5oBmAhoDqxcCwaS
QZ8Vt3vNyYu0/kjdGV8YQ3sqNGbrwa4enE/yCp/bJeolfk0EXBGgr0dwyG5Howjg
/i7XN5z5p3ihQCIwysQXl5jHxZRS3mBYJZvidmT7itjOWiHQBGpwd6zYEtqnJtCo
NJjfypH7su29aG5NHJ4xuV0mnap7Ludd4nZEXe61LEIZocED4/usjW/MxZ6gQVQ/
vwHEZNCT77QFA7Dm5ve4enXF5HgYxMf0lcPbNDpndBk4G+aK3UnHX1eS/m9+useo
Jn+/QwBA8nCPpqVRTgvvywTUqLEoTj/ZFmomOjz5C9SmOS7SQ4l6x8APINGd8AIN
kAuYwhVvHpHE3uCTD1kR6RqCDhiXTBWv0Z4pm1wtBJUEZVDBgjWGFwr4XWH0lk2I
p7pjr9+j8V5vsPCTVbgFhVHa5kBpbuXU9tOVrWodIILJF6rwrvIp6GisVn3F0+bl
cIm9VONCEWNTHaP0qEPwIePDOZlIYbeGy4SGpwk/UlfrZcd2PoAmjJvFittDU97W
ggX2Us3ucyTOpFt96gIaB+ZRGQ1n/2AhJAH7ZkS1GxWg8oljtcnQ9mjW2RnVrpfP
RdZlFZZFXB6fhjpERHQIEsM1wkRq52tLdzk3s2PhTZQFWpM3KGK1ZzIHsSqmI0mM
/Dj4FncI0eWeH9znQ114bxBq41ABCtoCrRkIMbe/YBd0QcnFWgrwASRf42w5t3sz
d1/cdHipME0OYu84YNPu+6uw42D56hzkB6ee21xJpbIt2bUR+xOurQpzF5qCG4/+
sVoYT/6S/psCkyaf5V/RABYqFn+O4Av+b4gswo1WxvP8bu/uJb6eM+fwuWmNrYKW
B37xY2T4mWbPvwN/U3jLmOe+LtaMxcT6cuZ88jLPpg0htXfom/mqsgIwLsgRp3U1
+c24SF+hULBkUVzUEIqMdIF3ONPOSVNM32AbN3QMT3wGbY61UYxFKf68VuP30U9b
Oi3j1tZyDowsNAIaLfhUEEhTa1LvsoL39ridsZlIfudvUcfEKN83g1GmssRBpXL4
8UlikRz4PXcQ1fWc/PAsb2eoVqsxbOHAZK+q3nd6u+1maN9Pqm4Yg4Jm7gyAZyCS
z0mLCXsdiMLdI25+liXIuDgo4pDmxi1S7B2YU46QCJh9k4hsLjTXa5VVEAImysbd
jEBGoVhHBezp3I2iaUsWEbBf+m/Y02xvAIQ+bJRLcXQNpUm0M1VQZCqjGe85/Ycq
e0reixf3UkFGjeAHCXPxR9z5Q/aCioBKdegiEwCQQS0y1ofryLMlZ1e5FBvPw5mV
rMsxPcAlOxXxG/8RABEMtspCnRra2BrappgTfp80wwpc2j7qt5Vt1GARMBHT6dFN
zqema6lprQZd2qma6g4orYiAoLkPgxhLJpvvjVbzJnIwKl63ZnMYoKhvDYc+JmOz
u3gFToviPxMf3aHHqqwu03mmuVq52J3g6aSe5qZbfrm6/+yi3VEKt0OQQc1frEr/
5xhhwXFNZ4IuDM8bY4vF+w==
`protect END_PROTECTED
