`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mmBUQvCiiQj/Iaxu0TiaM2hgcoq+ytzlLcRZ9swM1DVN8/QBUjvueKB/gw2UpCBX
Xt8qTqZYNNmzGCE1DtBbluBtZD3HSaTP9oF1aHb8wgq5q3NkrfNWrzW8OqGT6M+G
J+UMZm3O3s4pSaZ4b4+XF06/nohrf0i02jAxOM0M0FYDG8GZG6LoxWdqAtgrz0pq
dx7bTGrkKL6z6VxVPZEcT4grT+72gmjNj2BrUpilmT3u8My3UUDoNNQta4wI9D+H
TQgCJGeRDkHyIOUX5Hc7Nt4VnJeI1AXpUl3uE/go1tZcPAiVpLo/B6hFrQSnAItg
+HL5Qk7ggEncDFQwp6aDl2mUDRtG5Mt+sI8XYLDFys29BhGZm6wAbjmGz/rlP0/p
81GplDBekJQ03fqRIMTTVl3hFpSieXb/M8e9l6IGWBOCrHu9qQ3yOpHkSQAYR/lA
9h9OXCuE/F4ccX1dQWjaJm7hyL6S4IauzzIt5M2Si0Na9voViJ5bJ086k5HGWpLM
/4niZPzaUBN1uJpwP6dqNFYEFXaQPShtrgYM851ghlt7tIx9pCkxn5HlOW3kFR0b
bF5U8B/LeaMWewxQYGHdhOGvg8mu7X0LVZdaaokPpv8+z/0qLvs0PYswr/wuXTd9
bTH8bZor29kxeuWFbxW+FiXyqhVLA2/iicInHjOy2n6bbVmYoWj+rfvnM0mDfYPA
dImSh1YQiXXMcspK1GWobyXCFHFvyaFqea5dc23fqjbzoLlKBMimseJMU66opLAS
l9nyi6LTOIhE/QP70KZ0i8xm5Xf/voB8pWhTJUicypsCk14afFAPWT+rPRFKTV2r
qiCXo0H7bc8xNKAkykxxT1abK1oQ0jBlEyKloWYfi44Lnjr6plQnuZl4X4ZulPII
Eq4bLrGe+jLcQppL3nxuvqQVl95KXmMM5+rIyMva2485nKYCSf44qi25XEO4+M5K
Rup1gSpEsYT6f2wftUzkoyA5/uX7RTAnb7cy+QacyEfeEcnX4JX5zpgs0Wz+Suax
4wLY6qd96M4ZA3RBvzd3CXwFbxlXpUala8fUq0thldk40WPtX0pQfAx+Fdd7wZgb
`protect END_PROTECTED
