`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MfLq8q3dBrpQHkjZLMWTOV2hMMS2z8j7ujfxOwcH6l5wfjvag3sWQ35zNhtUhAte
kzpDCruJoWqE9vt8TBWZrAV7KSUiz5OF5Fuz6nXSicFHssnxUv2uLOKz7Y6qHYD8
hhR1VZ/E/csgtc9lPUr6MNoP7/p7w1dp9oatolFKX/5qMru0ZzIso6JU31kSxoP1
MzFOXYJdTHHMHY6Tyy8zCfz+B3ousKZTzKAMTBPWQJNGg7JGq9ZgdjK7GfMiYCNx
6bKXL579lZ0G0HntBAOQIKxVe5eDzwPElS/vzwOYqqocapuWyw+oA8wWg7NXJurF
FRzkpkrU3YTJndvxnLBg+G4iEGZgHpkucVfrHhPkFsjeYEZhbf+8jeIqOxjNtWhm
eEWyfyyiBRG5P1sdJpy0tPHLaJKlj+PgBCckj4vtkf8eX9Wq41smMWumwLucc5vJ
Oh0SXTQUT3B2tYqgWdY7jrWXVSHgzoWbUBiQ0H+eXDetrlTRSKjNOoHhRwKzBkNe
45Fjg9GLFwhRFm4a9kVf4u1Ll8YQS28vIqdSVAshgEd0k3tVBh6DIuz/iMd1fiHL
hCkdKjkaQ6F5SUx+0JzI8vPQL98YSBeAxKjlrJ09jfICbpDuSmiIkZpkLPKEOYdz
YWiIehv1MjGJlhjwFbC8Ig==
`protect END_PROTECTED
