`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8YELGQ2mKSBCLSQY0vjZ+TPhb0E6hBHVpxKSfZ8EPWx+KJG8Dpike9kqpH0y/+7h
POcrpg24bwwDOGd4LY9kBmngOuzvXjzIammTs7uu558u1qKiB0RqNbvAqb7lEnQb
xxzwwCJJ4XbvAACC6+TcU5Vy7k8fyXVl8hpnkITZRZbyDMpuHLcKzYAe5PTANl1g
oAaA76TQab8aiv+fzlEI3VIEwtwc8eBdR2WiaQQGe71C9D0xOxQkJUOlzVl7XYWT
opQihKC9p9QyaTEZUkm8EXPf78dCNHt98LzSRzx9wRlmwD8GUVm5o+gcYOO1JmMe
uhom/VwvpKp3Q2zK/NT5hzd1FWX2i/vZSiAAg9B9Zjfc+985vyuCd2UZRAw1CkEW
DqMv0ybgytJxBBdh6++UR41wGOOM5zOwwRAbkmDNFfVVr0EEHIwSylm6RGXsCy4a
Iqz2Lfg52y1OHV89yPsMmWWkbqVohnfQnI75C7O9+gMOMGsac11bAQmEZo6Jjt+3
xMAuvX5ICkH7nvHSwhRzXmyFklNKvwzaN/s14KPqbFBfjPBs0MrjW4ueZZyiUxcG
mPh7l90G61luHJ0Z1UM0JDMYuRBjcOKw6SxiZE0VLr70mzFQUdnMjFUJx4hYfPfr
sTmHSpnHrMwQehFOzEEEKu2qEc4mEWsteqZPS4oyZWeA6arGzfeOGmpLL1UhSoWs
XtnjJxQdwa6LLzXqiwLG+J0o2Br2X2afJaD4Gy4K3Tt26ITElMsDHxKjP/un184j
DyGtnMNHoXZ6ZzPX1cby9G+EOIBjBKgaSU+fLywMygtobPZwdrycTEZT5CJf0D06
E6rUHIBxlzfZefsACb8YWkBOwFX4MCgL1oycay0iPgJfxMknWSxIQm3rSteKeqKM
ma8ILLUquMZQWIHy9LBFjogqqpQQ/jF8fK8cuMQ4E0/e+9OoWryE8GZv7QGOJuuQ
F8jqrWLTdH842ndvGj3oA0pRdk0aVwphaDrVOsuX1cHqlOaXTp/V1ygIcX5YOzUf
PVE8RcWcGHjA2x51qflfTGiTKgoKYPuor8/SVOSZsQqT3TLPXisrqzhUDafav4c6
sZGzlspwEDJWSfKdsRyhk7y50D6szwyMbARoepjM2nYfBy7RaDWrHXXUQvegWk2s
uCQiNkbUuONwLOdkHcVJCdmYGn1ZIKBnE1XujOWpysPiYy/YIG7aCLCeQudH6yAo
+lKEjZGIWNYJDiCKjH0ymjpoVzk/vnWO/R5jj74XcxQd7/VCzlCtwKVrCx8B5nqV
5Z2a+t3FXUypB4wB42pD/lK30bTJwPnCUoMn7lTwnxTvWZ4tvG/RUOS4MHiO7lU8
sZthtYbF2kD7dbEZEtWDncuIFeH0M96i1j1fBU60rJxdi+1Pno5Lm17GeFPirIWW
+5aApq5MXH8azLIDc8PDncrm+l2kgzhzxKX2MRt6Uq8=
`protect END_PROTECTED
