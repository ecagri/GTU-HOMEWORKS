`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sm7WaJ1KL620jclqEuhTuACeLGFMHQry5J6md/bJYHdA/psEZUl3HRqMj6c24yz3
jSy4iNCp4QgJfKqHk+XNhbkMmUEjZKDpF6LLe5gN69V8vRRYjH7ONA0KqfUP5IGN
q5h1ZY1hyZvmWG5PKaMvDyxkUKTBLb6PFYchNkUxnHPCA1+MHD5H04bCaf15ySTl
NNvw0WoawhYUoAaFQ47cnGAptcD7ovHyMRijF7uu6murHMkQ7QdEYXvRaa6FZtVW
FVWTvGh9w9NIofJp/GG3j8uzdsFs2QjyUlJTr/9CoAbhIqPofiY2pRfsp+3BO95Z
zNbat7wKXbxd6aws8c9IomM0spQwFP/DBAHPPVfljP7JPL2qHjjSVt8XXa5yjILe
2VH+lA2SNum7Jx+AE9Zoge5LOtlJBEccCyuPktS+Z0qybE37y7EZCyh1xUctzhJl
8sbtPZ2BkLDAyNUP6uWQyoC4vjwuYtF2EnyEPYGEPRjg05p6PSUYRRaJfTCrCAor
bm44CkqBfeiFNjWIF36dNy5uBbzCDXTKG1fdwdeeP6Y+ZAvpYE+X1cqSsypWL+OE
tgjDr6wQacWdPvj6U0kL1mQzSxW3C4yxtSts6ZmgC0RCzXfCk+P11IX+vJ06nMia
+Ya/mz6ej5b6+JNb78KVpTejLvqKLC6L7fJy68zWS+nDKzAyaJsjhYKGoNBnkJBL
IVHkHqYvRw/J5kr9GGhxbE/2a5nC/ulugNcgndpRaBImxMaOjV4HgWly9FgpT1Ew
XScunNSARsRzUMhNLtAn5Q==
`protect END_PROTECTED
