`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gFc8ajx5i85ShhBw41RxH6ykpY5VUPpW7/7gvHInaRVoiOUjv6Cu98dwYUiXqB9M
dfa+5Z8ukuH31x0cqMMHD2fXg7KGXHZjbkfSfl/G+oUvY0MTosdketGQIG9vmrWp
FHWq/jacKewXHi65vSrNXnmHFqRLULC1JSVFr7z9GJ7IVoGAwSMgYe5JBsehqcjN
sqHxZZJAXL6z0zd/ss8iRERonrf5A5A+bmIAtZwMt4QiJsmtbyV2dIeKHx1abKW7
lkc9GyNuB+93SHqaWC+9133+34+ok287Tuoz4yCkzQsUwhlNVgFBP+Qi8UEhHvjm
pZyyf99cif6C+HMBsqHKvrmy9GBW4M21qDqBW5A2YX6zYWgqPnd0Rt73rIx21G6Z
TA7IXg55D2f9wFBuWHlPfnXW4ioWKQq0gsMHxuQwdi/9tygl0Fz+q1Sh6rPB7+o5
eJol9dMOkjT925VIKGE5at5Ni+DCGqC4/eQJWCZj4EJUBF6Q5gKgMmA3mEWtUfjO
l9l5Z0qxsOtBSS2QEq3BNFTazHWyJpjZCutqIvXaeZuvm3spHF1DeIJxaxBFvc1R
yxGq+/bJXbNmo542/FIcqSQwW/HkepHqDPaJ/p9b8xflNf3qSQ732HLVP4pU3NPD
1/GR+25sMPHSbzfnq5GGCd0R1vGSStPJ9ORud9r5uK1k6LdS7Rvc9BwEYxSX1p5M
2h91AUYNmohKih9EUnvSPceWE7sAcBwgKjJrwiySDrW6TuyZDVwf5qJehWGcOJaX
I2R9Otn847+BTdV5ujXzhVhpQU3FTN2SydbQ6O+9IFSXYuslx3H8g+WLdEyexPaP
HbBhBriJ4JedQQaPAO5CY7v1RCZ0PI+3Gzko6b3zdxv12lvtcr1BK2jkBBOl0/j6
Yskd1wNVCYsS3ivD2BI3QKtzsbYdZFRvs4jVVFNzNSd/omNg+0XXUtKpoIqk4I9Z
Xz8iTJX06oPnTcy9x9mK0CYkgr3sEYvn7DehLYUP6dlzldA7M0lO+U0x0oROsHsa
qckdvJwPQ7m6ruywyfmHfqxYz0P57fn3vXw/LK+wEHKJ5Wa3bvOxg0AFFejAXCgZ
XDMyVHXnxuxNer9k7s6qTB9s9jHvD55rNPy3/qr32t3+A9qOV2aCOCuchZSPeDl7
qZQ7hyvVmMOzC7jJcFZSsQFGZUySR9arEJYi7W8US4Owqr63Wz3s7N5YY36/kyhC
6kq1iOlpSPq0npqGoQGdmMbh/vPQr8iBCY+4NqYLR0cF4kflFsx6G4/4gwzFt75l
xbwJHR5e9mIClMmQSjrMbAZZXUbfYNxGL31ZM2+3EnApgNgxAmSETBNTeVNJZaN3
PR29TPQW6VmWBISHYKKmfhrety2XpjItfoq/tp4FRU74IrXsLAV6l4onv1y14C0l
yCppb9czlklnUMKbGb/LTinUczNmbMH24v5i0+5AV4J/fy4Ys2SLU1mkSort7Cbg
+bt73BT8xb+DTW7EvX3RquELYgK+AVBkHvLkp29M7azRY+yXHl3pMsmPEfp6uUVe
nAHqbgMlxZ6KMBDKcgBkYPW1/oda7kiXhEdwtv6V0T1xISecaAtE3Elp5+G9pmJD
71tIZOp19pwKDuTrWupI4zvEVRzz+psfWiFyv4dn3HrIPisfeLsid3BSaLwuGp4h
9flGdDUjnWjCZ8hzT1ojx7X0gzkSPIhhHu5t4SKiB9jwbNglfp2D1LWq+76TPWxO
DD6nBjk2WDowmrK+QmZer5C5poKAuLF/dB5/k9bIau0v7E8ypB5MDAlxjPvk/q0I
Le0/8hZL9iIqrDV1rod9aFyM0QD15lBpReS23v7Z3Wowa+NH/cBDD7EvaD/s7UQV
PcKkrWGYGVMDjfbHK6ERwhkmD7pt7yA5oCQ6tG8Bu6F297Eo3nM5K4AggjACLeC7
yjyFh5apsWHSPd3OO1rDGUzRvUJ2xltGhxc015mPBBk=
`protect END_PROTECTED
