`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GRK0P6AipUX58/JHBP7RoaljevVj4FRDLlyrEiLrCeaNDBI/5LCyQ4tcKYZQlWgp
mVjwBLuElSG7isNQkvfeBeRSahRphy/SdR7scNqfTQ3ALyKYbH/YSeXmSA+gp7h0
RLBH0ePhnv8U7D4a77jlmu2Ob8QV7hJkAreipuFkuJj8BGgm2GfoIyQOh8LpiEJX
ZSfBgo7/17RMJO6WPgAHbKq8xvuNU5xb5d9/PyGOuXPJkvOM8yCaTBQ2z2OTl8Au
IxuOdNyTXdgvzOigiX7xt+KOZpdvCiz8tDGHCBTL2Qk4XVPDXPfbvq9CmDWXUefY
0tGH+cBcNifHXvWsfFubRqnsUUu1KAAMaQdJeKaj+aBxiZFL7qXEYhCo0OZQqJzi
bLpN4D/D7DPQ35OUTZuJio3w4pd8HCq/+vO3ZbzgTDewCzrfMeTTJMYyCv76XOqk
DAHpc0mpaJ3dihdqdwbOzDMx4I39O7HYuIccNDFTxLi/818BA24ZfaGry5xSafgX
VYyQF6qw2XzqWqFsxAoiiAi8Mn3LyrKajqrcWJZvFPXEzRAKwbl3HOna8tsOe3qv
U18rC7TLFN7Jg0kGwh0oggtYnq9YqLlrCqWcD29mtkC1WrpkuCDWGOI6/QooL+Nd
IczLz9qAA0txfY48e1K4KrYJsngrySstDAhvd/3aeNu/70QvTEz6XMCgDixNJ1Ii
i6A3mdrs5KH99I96LC5mJxaJa5p7O6b2dbpD5L/KievBRB0FoOiMwayd12yjxknv
c5+5Hd66ackDBzT/JsAP3LiheU2b+UlqMPig+ucYQWdE40CVNVJ44V+YmYz612RR
jGAaAkI4lVSd/J9u93g9oA==
`protect END_PROTECTED
