`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vOTdnehihMHxBrq98sdQ5SmFwKEiXA64mIs5tzZEPQpM5YkYJ24Ri+pFVAGJbXlq
99cjjeLz0ebuu62otZtsm+4MwAoiHLEtulomcpid7ofN3V2Zsm0GZORlroPoMxjr
OSPglOqy6JVlcolCT4ZjtBS6C1048cB5wjLzBSkWuc6kXvciD1fH2TDf0X87qFPS
BA7yJu/3RNuh36x599hWlXL9Q1L8d7DXbsAbq+uyw3GM6hbIdzWcIZteIMZKf9eY
PU54jOCyjHJ8yYQijeWF/w+P2Sv9bVmW82K7ZgTNKNZsmHGkox17JHFBO747kYuF
Z1HgM1jlsILIEfRlLvBsxDLCHWzRCWiXsLtT/IVffnMKgDdjSU5FVzroc99yjCNJ
KfF86IIs021Ipiqm/SFhkx71yNButvD3ywT5bzuvpwGSUTA2kpzGBFFOxFykspEF
hEUyxiym/z9hRAbQa/edLKQ3lsfVgBTfG9vED6CYD95RFVI4DvEMZTZ3fyztqbEm
aT3whKREZhOOKyD42t5VNaeiKS35ijJZ6UN64t8RlnA=
`protect END_PROTECTED
