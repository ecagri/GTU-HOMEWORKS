`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c8HplvIGEx3wO3tweaAxBsXDpkoR/L99741FrQFrzMptq5m9dJ3HuXrzChCbd6BB
wgrnpCWz6uugNdJzYxWJGMztkpZVRdwnpDDGCncKXCxjEMR725Rvd6YhiiFgP7hi
QFWeB3hOdQL0qNlK0v4YpOr8Mq73Z5UYPTbFimsJqL/hOL0/AlLETdq2JMzJ4VCO
clR6o3sslTvZGFU6eHTAMUDo0nKE2Yr4ASduRzfRdzzE9UP/yD2CdhUdjaSiFOZD
1C5iPEGofY6ugx3m9m63VsPJLGQVjncsomFk/Z8N6ghppUAj6MfBW44ynryQUCr6
rKgL9nXxG/NfYjcRfQgNe2IBd4FjwEU52Ci27OXD+IxYegMUYNrn+et2Jqs5ENcr
wEylEgEfj4naod/QAlKAiraT5niOavF3KUy9aALzFbuyNeYXKe2oS/SLmomk3HAA
v/g95aRLAWXq7JjAfCub6v9OR8jFyU70pJPRj+nJyXG5C1UyAQSOn+XsRLGiKjm9
YWdYUDNid6sO7blgb8lD3NguYKwwCv2imfT0l9iZb5YVoDywbq8l0kZkGwBT9e4R
S26A+dREqaDZqDtp3voUWbvb61DpzBhsbgv4Yvif87R1LU1OCybzFNzogbAZcUoZ
T/VffQc1a5mjhE621E3p5pKlfuYze3uvA6n+m5FNRDvwEaHuxKWBxbhGHf1eqDMQ
GPATfvLCHAhqZJ4sa7jpZROUHpgLW4dYfZEl+t+vZZNrsb4Pg0/uBdMIXp8Im14D
eMqCqRX46OBpEi+IiNbpI6UGM2Z8sf5bNengUulvUOdixmeJ/roZyPzt8bS65iAT
QVfk4Ft63JFDiOoaCgdvdQ2DeKz7ZooChDNsv58fRCDHu0J0+MtRA0GytzXfGpQP
6sJsbAkyFcIh32bDmgjZf0a9fiJ4/9vDLkkBQWyX2c+V5kltQBIC1qm6sZd75A8X
vbBtiIdYNQzIUqOADVVBvn/UkZybhYPae//FLilVHquj0A97/z0mfb0mgnaGIQwH
K69hVaAZQJyCJFcqiPzyIMNxtC/6jJRocfOxXmW/zQ5QJQs7sSDHpFMLFf3JKu/b
QyW2Ozhx57WQSPWBiogXTeqFd+Z7mpXN4Kw7jmYLKkKfnyDP0+A27tGBdMVK8Kk3
EUU5dime5tHY/O2JlNxfBVYdFe9Z4ktujpz2VvGuQ9lTNXk7gxCGztExkMrco0zE
mJn6qBDMhIGk3gYfw1paCA2ciHYu3qTmFuc9DGRIUXrNO6tWti/Vz5JlTgTvLkXJ
6z9VKgTdZX+SmawIAcjwTqRXdZDsjbba+DQWDlGTPtHDiEKpClEP3BtgMBuw9CFL
x6yLdbf+CTu60Z7L5QytnEUdtPY7tS6J7sZZZ0RSfYj9BWx9TKEvW/yWbtVbe615
57RiOGz3kmXXSaA1s8OtQZ34Ppme/AKHAqdgJziYpOQ4wRDl4syx/0uT04yu/+Z5
`protect END_PROTECTED
