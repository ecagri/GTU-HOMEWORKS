`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rCfBxJOkcBZyCJsdZf/PpJdMXMzC6Fat0/s0p48O8oDq9XgH5OpSfAyHAZTXBG4J
y7pALFtGnyRe41md7DZ+kyswlKlFRptWRpEME+K7uphs4L99xjdGwKMZvI9ikI2d
BZOJ5rjwB/lMQMKJaTSubkkb+YI96LhHU5h2KK50I6NZ6jFqwpGb9+DnJxhP/GfN
B1J0o9Tbjtee8AX21OD+dJXXhx9ufEB+8tqUndmU7KkCHaS7tL1kfz2+eHyCABPb
bYfFdEKkaDlCX6DvwBheFSGSg3EC88+NBVtUzstQzuvJQ7/NuUKsXEMZpCKyIh13
s2lNyGtVfTdeM50DBlPQMpKjlNiKzCMAI3MM27Ltj4YSMkezZnZ5/WSu86jUvpXc
AwjGb7yj3SMb8HIiSyAiMJ6skBlmcamgaCF/A9/LxuYr2cQjeTacQuXC+6vAWJ+N
rPBI2nXxHRmUtlWK/ADLs//NvrNV/W2o4+q5Juq8H7nSZ8XhW4DnhuZHTg9snqi1
zJSYt+5isx9O2q2e8k1Ydgj+scGggBGuksjF0brokiDxHP2kqGgAGRfJYWOwnv+4
DCBbp5lNnIU8RQvMn9J3ldzIXMwXOcYfyV5SHkpHFP25uqmgFKHlwC0yfgftS/dR
hxEg4Wkt76l9hkarHb+jNM2rhHKJbgLbg9V2gOxo13fT8vcE1TRV2G2CIDTVhTg8
/fzfhAbAOJz0R7P55mxNPLzobRJYbEMM27S8UNu5ZsAyLgWhCkx3VGqzwqx5q7r9
yj9IkBL14HLULx0kB9f+T/7VZu3sUG7Lh3T92OsnyHP4b76gDcTygt0grJggKRAT
V7HXMn0m/xtUrZPv17oX/hdBEhETBG9xbzOe8ua0x5OfAhk8/LlnTF7bI/acsCNo
s1gZjQy9XhwbuxvOdFEsrCllA/5fLZiKycm2fX5MRgDBSrtJx4JDgBn+DT3yvmUd
HuNuA4Ink8WVZ8EU17QoDbfzdN4ZG9RnQPzlA4u1AiSaLMSWUZMtLDyNubP0fg63
5cvnkBJQCyOE0MmZXKVPSTLV8QzLvMQrkqI02GjwOIfQ6Wanoy4BPN3Lhkor7tXq
Os2Kpei+qRZbDiwGTMcfCdf9YrVL7hcVl9LmqHACQhHivbuCz37RNQ3r9JfRjjVU
UKvreYpquV2XU7fMc5stLeaA2fVpH7Vujfqn1jj4GL2bXzY0DQ7QBWv7IDVCpkSM
fYrCYep70arF1jTV02Vj+UQ1w9vsLkTVZ+QJ4UNZ/VcOttLl+rEE89bfKjsr0igl
dtKmXCtfW/DxpP/EvyPk4ouxdwqQtGww+P+nLVuhqiItlPHqGo53sKLVoMUj9Aa6
ebhZVv6YImVK8zwQaJiM106xp7NPYARoRc1qHzvAS69KxV8d/3CYP4x+VCuTL5b9
IyX8W2XbTOTKo7ik/UT17ec70BewlfIK0cuQfGxUuU2t48Vi0pIPvetkwPn0k7Y+
TtWMqgJOk1TTspgkGOV/g3oU59Mu07SV8j6ot4Lr8ITmWq/DqqV8bFEMEJHkWoVY
f4C2y6Dr/Bb6laHAkQDiCpfMcKaWKEetZLopnRKeJc2LK3pFHozRq1QnEXPI0pWc
phlCUIksCtqeUvl2881wGUm6vRGz6e2QCmJzGIZ24Q0onts5djujTwoZFcFLCMd2
O0Zsmflm2c+9JQGoFbdRlOxamBj7SJmB5n6bE7gTxEASmuG00LljQE/UlQGQRu8C
i6ZeS3KcaN5/WfwIsPhLJkc7C6DqmUBmFGAN+QGIlH9mgK82yVM9r0hgtJyw+4hA
QAY6I+ZD24PtZyNthnk6uJJ+OGxfCeCQ+hSskJpTQxdOjtgslj8yCJla1s5lB/1j
cFXlNHaneavM4A7RUl9nOb1kqsXxpdkG9tG0pL5e+i5D0n8aT5K25aEAE682TrR/
E1P9owxq2QJ6y4R4J1aE8Key+wYvXxa7zPrYnB7vAn1+1BbVdLgP2PWu3ptxVPOI
8GcHYXOEBf8tDkaBDJzM6KvHmhlUa/ttn9udvbln2Rd+GybxFPvBhERcbf00kvcx
DVT9B5dJfAFME85k4bOq+G3t0E0oxg2n8KnWoB1eIBz2LK6FeNRtkmS0JaEB53A7
ZGkKJvcs+kP2Y/NLvcUNT74Y6aLVzBHOVrVA5QIrcjn2IW8rpzMKRA3Jez4o0TBQ
Cx3r1pkP+681Q0fV7o5+XJj/c+pr6/TvjeWkwvIHFURHW69sU9+dhVricW1at9Xf
JbGFg5tkCdbHGZ8X1UvbSzQcnoSKTN0TAEem/lc6K1Ngp0eb8ZqVVeICrsTNjDmv
L0cex2libMRwIt3onjR98AA7Js6G5aSGKEHQZJCnuuQEssRfawK6GLrExeHVj7Ga
X0o0YSYleSPYLJ/SYG56K/dmohz8yp/RDxZ2BqEP+7v/7Q7mRHbFz5bMe/352vAd
BBmDDbfb0Ze4BZRzB23yIW0J3AF8HT+sPiz4bg1dzw4kTZYdHz346ykfLY8KiKf8
DFnorIu1ioE0CKFs6yfiFEybsT59kqelpigKW/JavbmsNAkmMBqB5ct7Xi28fJj3
j93R7xMFhEWv9MR7J9rwC9nfWWCIRcV8YHY+lppuktLG6MLuMbkY01DlziRHeCgQ
2YTUc154fVNTGAXFfNvJzLEdybWgHuIPUjG4+sgn7etrd2Min4pkTgZFT2SjC28x
oLayzRCBHet/SqIbqs4U0GpPs9ZeYdWZXJAkar0W6/36dXlusB5dA5Xtg82LKbhw
Bep2dZXoQCVcHdMcw1DAXPxyjRnJo/Fup+mdXjhJm133xZnAtVQ6bQaBxc0dd6Pj
dTzm5SiBdROmS+dJBSP1ROw8wxDWG9etH2hi56Xhx3/ypLazCc8cIVBiQbos9zdd
Uj836TLy5Jme21yh+hepqARaYq1WOLT+r2ihdiHbkFl88IyrL+im4eDNoNqUqGc6
b5iPr+sCZnb4o36KacqCUE9zVdyOzXUQmaOVizQSb56IKe9Jk+tLsyd5/V8+JGwG
cWWwF7QTZj31VckPHZ860PWqrxYIKa37IWG3nUMQrsZKFMNkDXfXpb1OGdRyhM6k
xvGyZKObTFA941SQ5Cq2xoXhba4HOX+V86MzZlo+eMM+DweJImkuGNEjmM7wf+AR
yu/MMYPyzadmYvrv/yD7vQIOyQcTBdXvDCdM/rlWRMlZB5adEY1hiMSb6q6FOTHv
ZSN7s6Pg945HSblcIJ2FsyJngEGCJ/EmnLIgNdZu6s/RyAJx0g72aafSP/MYYJdO
Ci9GZEu8MhwdU73fWlQRZeV7A2YXjhTjXahA+U+M78pLtML5hPp3HO9oRE9nJNu0
iHpUzHJRRdT5Qqi8VeExGQmOCu1N2lWBPiBDmwRHnI2dO62/woesEWocvC2PkiK1
CfX0foPI9N+4OYbQ9XaD5+e3mUoYCa5rb3IxckH5zL2xqvI76IaI8wIllraUJSgQ
A7iW8LhiMOKMYb/qr3frPDVGD2ahlmR7xg+Dt3TxozTNXp8D4EIRGDUgozcI3Ay9
ZPNMFUrJyTSzFOvdPAJj9y4dZMYsCq/pEkOQANOL325zrhEO6GWW4zw6IRTKXG5L
Wz4yGPClbltZnbWUmPW9ngOluWAAzygpbDZqO+F0B+LJ2X+vFIM6wr3DcC6/KjxC
vtGfFz1W6P1rfz9Z5OwYRGtHa581PHMAimXzp6xm1Ra5KFMaQ+bjtYbFcHXqSAkb
zcSoW+5aM8Ca8nf4XLBa3MKBYyuTxBNpbRBZz4NYLGZKApTW37sNXk2hRDihSQQz
ll+1Tw6OffHlAp2ZE5UtoA==
`protect END_PROTECTED
