`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OnNVanEyUnO4tPqZOCaOSiY4a9gGCT7uojpkLwJ6R4at/fByee9r1263YrAkhY3o
g9UCcuoXBlaMI5EybUKsupWsPXScbxcQx5zG5PvUdQfr6g1TqKlBMIO147FCIZGD
PjHL5RPvq2mNrVg2nzp1eWv20KIxDGjtQGnJ9/4kqCiF6s6LtNjKvJx6YR9M92Jf
HEOukWDTyust/FgSQ75G9z+GsmmBV1fpfSyUOg703smQJlM0Kas5Sgx54+bGpkHd
sIrEVByRUafXnTMyAQwOBpSAwsbV7KTLaTvJ0vYl2Gvi9Q2T9QLiWIOiQJNW62Fi
P44guktAHwCHQuEPWFBqdexewOHcWiRvsS2RuC/w3InwdE5NdQ0IaKADWuCNOqx8
/qfuC3nv/YrFvHsd4NuCTlkcPAuj96dkM6Fum02qI+uARYBtpK1YikcHIk/blqgF
m1iywpDIRz/4oKvuuPpjIKNQ/S84GH8dcU5EBJkDxEaem0V+C2MU2g5JSvlGCmbO
TowvydLgI5wvZTRkokcb0GvroNDVN0suwFcScF4X1ZEJbqguhemBpVOfgnDxuu+8
y8fnOkWgY6fQNld0OlztIQ5/igmcbXmbeIOvOkFKWrUkvKorPkH03WhLLIpBZlLv
IVZ+FSCmPddhy58sjrulgVLe4llek90n3K7LgV5x+AKF0Iku2u9d6V+qfWWCSVw1
XBWoN8gJ8Ia0cIZpWdJYpamNJbIzlGIuSIyW2lBMJ5MLOrcHk7qWmOHNVoJY9vax
1R0ryYNlh2mNUliMOg4cMTQmMX9j79adOAaTGjkMEtsascVcNJGuU4vBegiv473L
xugF5OhiHVygnd4JPi5Gq1d27LgWAei7krcI0x2XJSBWmIAP3oriXLBNr9R9Jbhe
uy1fffQk8Tv8DRbWsUUMG+kzHJXSONm3htWqpqQ1cSGoeoY4nQB17aDcAuQCxLru
0M3Ju7APMoC/ecpmGLVpxse3DWAkcnhcUF3DJhaJ/p6r22wbbJC4X3PaURX9rIJL
41vshRko3TGREo03wmHi0IN5v0hnrNnSVP26qBOaqZnMRFP4jjEfW+v1DJJ7VDWE
6N9YjjnE7uZNeTQkpnHUtdNT9xPdMqGLfkY1m324zu//e3DPT+IG7iIScZicd/IJ
D/4sWyoyNMmMaIjqkFGXJ58Q0t9OX7fpjj8Qz3Xj6BbkFLVto+eF3oLyeCXZ5qzU
GC8UMgAy3BWBsI8KRyGy2vYMjS0VspiFHtc6BhSInFzHLxyUOaApVjeIoaWTgtI4
gIXfBy/eBEEuBgM+vTYRd75rivECl9yC0mAhyqCSOOE0oYMgbmjMjhyf1NJxzmg2
AZQM9fgHsznz9PIihJwVnJvWLUUMO4V/L+EF+l2RLdzWQ24Uo4K4eqgSZMyqpr+/
sa4SlgxHcTsz6iXngpJPU++bd+Pu+pn1vaJ3feE1V2S1GzoFWfG49eC2NO+UcTOg
YYlEYkCYCLQjn39uypfEjRslw7aus3wsvbh2D/xwt9LSVKSUBcUZRGMpL4BWvSTk
2Dc3tY1C/maFFctPx7wW11Qc4O4wNW3VfEEAljCJtPP4HV5lJG/HtEGN+lHtEuW0
81xPu80dhpzCFA80jp/yV+ZU56BP3xuOWb6QreLVNaZ5HXgYQs7/z827AfPvzQpa
/VxfXT3B7nw69QqNBHVTPJCKPzcyMSbSIuMj1aOyGAsfayQzMgi5Vvr34nsIExZj
v2G2RMpac7+AM9sx4YOt2ah1F6vEodK4z+lTcGhLUZtgHbGMwRo1x/wWKUkbql6v
lMfDc4XqBiXh4ZTNBreq8vIJJUO4GSYf6k6e8/TucAwn2XjST1d80s5pAPmikDrM
VEk9sB2nIyKwww2ARdCqLshB2DlVCLrfYVclaFzUv75+g3UTaG1PHIa6ARdriGwN
o4ME0alHLuwr/HFmCNMxpc/R4yObncD1P+j4VOmXGOnugVkKd+cAM4deiFF5yxhR
Y9XbX29Sr8sl2YTTckz4RbgTzVszJDCNpXSeFm9AOtiGSAkS8M/akhDanoecyeyf
eB7KEHCfWFnFdu0JoTHGe8gJ+ypiWNcApS3UHYhksMaX8LIIJLLozf7aMMuuX9f5
Op9a/k3qhWmf9/ySzH1aNosd1xb9c+UV+VPGw6p6KAKey5leZwp7sNKDwlII97lG
iHCJmodK3YRUTGLdrif0fUOmbUZ0xdVIFHgySQbQDg2+f8fggRPcXwM2rcvMFV5x
M2WYD7gcxV7UhSC5SpCrf0ssUrIaOLYRPurNae0dwBmmpGwtmYYW603QM4qfWX3O
P/p1mpOipcRBjZF9uPurRe4RIX58osRLBUXi9M30jZX+DUvEuXfFp/OaQVM2fKmj
Tx/UznjwLHtB+mU+xFunbYubE5lNjRIBQhVFzOVQF54hr4lq57GglA3PUBbWZ1mP
DnbAnLsX1Xa3ra99OoRQZ9V0u75nSokdx5/siOVOzizzd/HUdvJVts/EmzEQw5w3
TyPxEE6Nh/y5gpDIgE7UcqLJX4aALptxTkSnE8K2VQfceNeeeu8r5HrJtv3nMlaG
6Sc+1s2cfpM8LNrhxaookuCBur/t24leAB4hlZu/55rqLZcS5BUOoCTT8zrlI8/2
weVqsB+FHjFvmRlIFgpKTgakMxeoFFl13FfJSCpr9Yuyh5TGjXOgca8WIKkNnPyS
3OES7UtsXWa1W8Dl05hDtLVWzfQpdHW5n5helAV3WGOpcKV5VQJv4YuixyqB/20c
21YKhzJzna4Vu89pGIg+IrqVWKnjkpoUKIgyOWedFVDqhSmzurUshSl4mX0CMVeB
G9KOok9aBOmTuSta2OR7CRbieimcF7X87hq2sL5M4JexZVDJoXdp7pqyVBeM/5W1
WDunD1FIeJdK+OqxmvHFLgtcoMEuS757K+Nz1+pVCU0v+1O43amsrIJt5AvH+Iuq
BpP2PcZrYv4rOiURauJ+iE+kL1sYjyFV0OjJAbMPmanDh3aZcuJ3hlzp6tgMCqKm
`protect END_PROTECTED
