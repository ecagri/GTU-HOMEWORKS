`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uQniBZOAgsaNbp0XwxUdZGZhjX4irf1ZVFJIc/PQGF5ysjSctl8O2P4HbR+pG2zx
azs/cMnllqNfo+kldSf33AjkGoYUq9kOQ12ax8AW8kmWuJqNkx4lnyYSrwSFUX15
zT2yApSjpmuzKJ1yif1YjnPUzg7xY/MPmRGYd2yhPzAV9cinTtrZbdGn9sL2idqc
3+GsaFkJgeKm+b7siCeffXVxWvPW4ZF2q66AQW99jYc7T4vU8+Z1a7xV8wcOw/ds
igiHQPOV3lBr7ltewNe4hNvYiU2tObExewgEkaVeOwQXRZmQqFZsGXeDY/PzrmFi
5Hy1RwxPKtNumzDdYk2JGbaM6+QeNi4xk80KhBE6O6eKFVM17UnVZf2qg2X7qxxn
7f33HHcOBYsauJ+GvsiddMnlhBRBI/FZ2Y7mnZw7wTLDoZXSyrsvK5LqjvccCMwt
iPy50NKbI8ijuCkDsp/atNwGTpXp6voZ2+6BY00edC95e1jyF9adBNBY2VuH1Uq3
inckwSj7Vri9AI3PnWsKYr59NUpdSnKZaUhSkeYr7Wm09CSZp/VKSDr0UnPs175S
bHkZ7SnOvWKM+7+SNW4+8/5Wnfu21rkuGlrhpXORn1wZz4KSmuobzcKhuxRTAab6
H6smagl0r+qJTQwz4meQ23VrAjGBEu7iw6z6awrf7TFaxz53bfgiVY180vl//SUS
HlIjzEGl/R0AoGfkL/9ETVuTINMfsK35Vg7+jusZZaTiLRkElUBT/kB7rFI6X0M7
/9UlFwcn4lPYPM2jtRbojzT/n054jl2IboGSiQHXEJVWKrLpeshJFNwwI9tcQ2aU
5nHgL5GFkfAdTfPQIkZdovGQN2nQv9KW47Xz1dv4QWfL6gIybjEitYvwDn5nb5TY
JpnhleDxIjy0qT6XGbBYI9/HAQ4aX3ZGqAJcnfOo7a5MJkwzRPTp0i7ZyOwjpD2v
HQ4h/raXObjYCW8HrkfnU9FIlzxZh3xRN51Z7rx/CXGN3PYGXO2CpEIrCCIGPsCM
Jt9WuKnLF6fhWpvZI2othUkfhBBqg0ZIBRBCyQ4MEAOYmYTsSW919uDp8Dyr5lD1
45bpF4cPrlUfPyYm3qB9yT943vVZ+iVLOus1LA+z7rDTZOBDs0v9EesEjgHMuwHi
cNMSmD1pwl1ovgW6z1jSJe3B/2fogmQPbRqOtSOuvovOzy0+VrIcFt2kJm8C2gja
dqOJhTlhK3K/OSmyuspTtCKhLJiCjqh3z9Irykq1beChTC0TBFiLRjKi9DvUQrqx
EVZeZwQY6UEOR3MdKFgYFH3AbAt5dTAjKRE6gk0QtQ3TuNmvNpjTY4yLy5PrdPqz
V43GI8bwBt3vfRg2Oa/OtLEN+sW9xiyX68xxQIA+2rt53VQGJaMQsluIS9dXb/rw
oA2SA/qnh9QeQYPnjgFcxUryRiSOrY5Cx1Qb/KuYx+nPHzoP/FIZ+SRHvzfbIYXr
aA7RgRI0M8tux6rdlBjStirMOgQpbjC9pGisWeKAO7wkpA9sp+EK0RfFneaEdNA3
anvZEkx5Ww5vKsbW5CQdQISj6EIH4/VJLVVhGpCZ6RyliZ46tqOGfyztO9TFWpIf
vqvOMB201tmseVSFCaxs4/iL6djuUBGYQFplRrGx/8NypxeqTf6UfmFNTyRqbLF1
vfiOmFCh5sD2RpWh/fg2E5OaOsWfZ7YRnfdwv5puFgB4Z/Km3vo1IYTRYblKyFcW
mIhdPPTN9th9wcBwjq4GJDW+ff6h6zCuaBAaAo33A+rEC9vrw1zqFNW8CHrOriYV
H55epSv6Arheiu8+gWUKHp/8jmMVTHPXQaJmVYBq8rhzw1LT7qhFJ6RL3qNugvUc
vxl1Ekj5zdpYxGHn/7XSAgk5BfQTzFkl4WuowO/AfVa68uF9UeJv3ASKJ07S/Hm6
P4QXh6TWCo52MxXmsKrzqKzk6Z0Olj5/zIdvC69vRdlQ9piHTVo8FmQU+iR0M6KK
`protect END_PROTECTED
