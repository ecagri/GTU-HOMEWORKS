`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XfCReNmcPwoDgDNP7onDM/0aWdFJyhP3wcwhrv7IRjyGirkiDNMUUTx/NMHgu+Ry
lvA/qUoQphRGsR7I93ja/F4mo/ilfj/KfKVtqkuuEbhwYJRm0y1cpadTjafqgA8e
tbGxjNav+nz8aBeB7v2QNOHOtfnT6rpNUNKzxeBQERYxwxXHnuxLzDNjJmI6dht+
Vw2zt/jyz/+rk/fP8OmgEsIjrMEp6mEp97BmIBJPdq1pwwSZHSMd5o9hRzS3Vr0v
rujZ72O8X97S7G1j5H1fubM1ZSu4yZipKlNrBvnOVecjeCpNXbpBgU5AWw9lKqtn
HQ88P1P3P7y3M+Glhh60aKb8HpeSZzM30P2CyPKQpU+tNIOFf6U/In9RJODGxVcm
TQFl7/J4P4jF6kXdmzo9N/z87JQuqg55m05tZQJgrpSKK9QY13/xhhi7w/S185TH
AkIGQrPavOWGVv9ElXSsgszK4KSxl9rck082paJe0DMl8rtCFDpXxfKpKq0F66zy
BTQ7ytwNnBT0M5WJMmuJRt4yqZgfU0PKtBf3EQJAiewFC5OiTp4FD6yT1tGESt6O
lZu/6aTVklQptLHQY2OqbLSYxR3/w4kufeC5RJ8yzXlI9b8/ZnBdgELujw6eTQrk
Mi5adO7dLlEM1FxuXxZMr1etC7qKVO9ZwQzWXy7a3/WISzTt7puYfFOx7LNXycxI
sbRzHf8MvkcscTKtkh1MVa9ca3sMVy6711Wvjyt6zeUolTtcnNWCKRI55u9i+CgJ
KAsBCqwEtyphEYd3m5LzFPU/DeRYFju8buFyWqvEltLpTkHBp441smFjygVRmZbS
WbDpLMBX4HLM6BYrvKYp9ORL08QtxKmV/Nc1JOOO0Q+HPM3tIwC+sHtQmYALFLJy
wBmWoQ1aUTPaML+1TArx8EpPpZKQrKumu2wNu/lzcbDdk7qMbgFNYfANL1tca5mq
5+kBZDE7ZLEnTbr3+4A0NmJ/zEy5AZ9smRdiY1I5N2Q3OHpJsZ7tgXyh87MD3TX5
bS6ZgdTlGL9f959iubNvp9j1i6B41TOj+/LqpAHe7cLSoASjuhE9CZwMku5GUW7d
NqAqhxDuJ4dhCOM/OH+FWpxhsGmLZgOVsBGKzEiVRTwQxOeVWVEtlWbjEb0OQHKi
+WHqjmcJGFUFDjzc6YLF+bja1DOgTB0OkOza9BMZOGChEyWELfECZ7BGAuMzMxBr
1HwqZn8AkOtcI754jNe2UW0o4z7o15fPdLYnTIbLjJ+3bGmrtc/hKm4sbFBmIJog
2N9Rij2auyzOW3lLFVEYSWWHSNWN6viNGQbuCy22uWCVPfqhS7gqgSxWPw5fMZaQ
cbXbL7/qVDPKMkhYv2wi1mQbVV/phjIJ2L4e/ZZx5ssNyczHyUEpS3vbkoBzGi0u
GKGvUZsvI5toXXABGfa2GB3gqX7GtIYnXJoq5twiCvFLLnxxnfOAqjJ/dMFuctNG
YFrlaAU8g9Lo5h0PLhZUTCrCoR7tDX2M0pAoH2fuT9bvaMVXKOiSOwjsvEgr/fHu
0oEqy3obVMatWjP2gNjUjvXUj4zN9Bf2wtd1R5qwNGLHjB1A+RfYtiNRFDrvrolJ
0bYRHYYNDZE6IrDrBdA83NRKW6xIljwZmS83igny9HpGVpWUJiA4Yi8oaEfwlfQe
VITd+GcU5bReX1H2phgDaYNuWpW7A3UVrIqdoTzqd6/6a9idLGaWdTSPM9lDXTrp
AmFtH+S41BzNl0DR6JPzj2Smw/NO857dfk9kIEkno77ITuP3PIC9t+UfGVw1ydO6
zOGB7LYMmtWy/Vp0KTyAQxy+aQFiLu9rnH5qN7lMLuW8HyG3xp+O4FoOnYuF36Td
S8nVbpkCLTc9KKNlilm/U/dp9gpx+bnpBc/a0MY+RdEHFtN8ELLFP/bKdTnqlo9R
ShH+YDtIHOyDxPXkCSeRRYBJUXwZDMU0vOc1BeBNctoKyodmW/2iXNAFDAi3EVcC
n2UfCNaG/Xpyu4f79dhaZToFrzr1IxRcS/vtUqLuGlGi65epBe802+HioZ+gns4q
7U28nYbTsUE27JK0C/mTzwsQayvvpjBFJOPUqGMg80F+Lkzjc1pN7A6pQgFE4okT
13t3eop9LWkFJ69xExekhqf1qnsGRBo68nhkKDYXoPZ7k6ifbxPX9DRQoaUeoSCW
rTeHRfAmBZ1v+i6wINWgJ7jfFCUY9AxJv0S05oXqZwnhYvlDcOrp4G4DqREk6tz6
/HkWSZMvkHW2uPrLuZ+aRBm//71QRAo4uC4XGXVTB0iY2/nZHMvVZUE4zvfL4DZ1
FDTAsYOLxUNgxIcr2qOH0Qo0pFXQwMIPO8O6j5wwAuYbRpvQpduLa3F2Y+gapbCQ
IIzjKKe19sXArQhzVbtaCcKIDfe5rHv5xi2r/iLfeBmyRy4+HyWGA0hO4QMbXpn2
cMS4BCW3oLX7zHlYK0Tb/d1wMkwnW7O83XOJS+/NLMpZbymH1uIVyjjhfwyNU0DT
wed9aBcf9GNu2qOi326yVQXjDsk5ejvm8qQ+KuK/FUiWlicxLrueUNCALBJ+JzA5
HHAl2ewuEo9umLv960hzzGbAGRBDtq8mxliErB+RVPPySODOpecvJefR5K6TFz09
/EFv5RuUamV1JigEXgYvq35xbHRYalW4A/SOJjXTT8X5Q/X2XQO71phlUwcywFk9
wjuyIleoB8oFChX5VY93Worc8NMXFklSMrlR4ltD92bDmQYd86aahJSXiWnXMPDl
qD+tzA15ILD5Zwhe60N85DxypJs+AOFHiEiZmIuv9VnVYbmw3FR1kkv7NPfxPXCI
QwUpxs8Ovay+CE1dU2dYlgJHAJ4ZEfewS/0Bxt0th5tUzBtMKaM+GgGKAo4y+qpg
jRBfGySonfBr0AfZGEDbg+H3x/KQm4z9t3XVJv/C/zNkHgCpOfdELiS1I9ka7+Yd
bGHvgSWI9cTlegIKYaKSu6KM1swGrZxgUqWyL6JJyipImL/oQX/GN7ic5I/VxkIT
hQ8gs50zEcYrEUB3Kc8MHxOmVESI0eOMMNYy9aRrFIyuykIXDrHq9PF8ZLV+hIHu
EGVVHvuNRI0Lj6c31615B2fCKwkQE8+eQpIO7t+ShPQ7N7l6tuZHWL5Mz6BbdOrt
aPR4fDZIEgeS0Hb01y84pn/TzjrWqf011BsEvzjpjmQeZcju510iPD5PVdecqTBQ
7x7l33Pg3R1wozkehCg7svLCeSlqzQhoS8fyRukN0748o7AWXkWho7qm1RxTan+D
quizlQAnSiIByBMfI+Uu+7QweBAt8wwyrYZ4sQJNxYIuhlppX4MGuyD7RsYTCR34
pl6BfwrnkkG9/TYLBm9Y15TFb+cvCPf63UpfzwXF/GhLmsQbqwPBevrnQYB/jWQ+
1t8isAl/XvXS1AfjZTscG0ZxqyIRwPSe5B8xmyZ2ld9NhzLl9dF/ISBR8tmbiOaz
0A9x/xH12gf/f/k3y1e8KuA67w3gOMwBmAIcIInsmgb854InsDxQ1vilA+OZjNpq
ZHc/tTcLo7I9xk6OIWzBs+Qfujzd59syiJWYzq2OoNge5V6RGjhA7+UijW2yuseM
+QPymStix4XtGcosoQgeqC1IazBF5I6H/CE3WNFhpE24dar3P2qDr3mn3amwy2R8
h24re2O+6FkVeA8GRp6uiMUwHAQBSfj6oPffG3cfetbftBDE7eNgSLiDYRIQvZaM
rlwb9oZKNVJpwIrWa/bwdxyJTwPo8lt1DfiYYPoTSWrBLsElysNFK8wibhFxzdYL
dTGMe3gEiW01kaVSL1448qBk9Mv7/Fud5ZluQxsJfHBLyJyG19bw7zZqetgsvIvX
6lvo+oAAzEfJrajAVzBQcLRv9msx7Fk68lPXVJdloYc7aQaedm6kncQGjk+s86zH
sDeJnhCpO5YsczXkhjqWG94ATlIvXNNOodvcjHw5ymP/DDb9w6r2sSHQ8FkCv1WN
UksWWG5yo3/PGWQMaYEmeVOlimBbPnv2Vuu28CWCDn/7s74vCN2ymBxZP6JNUIyl
rXc/ElO53eHbYmpl2sUsd+6fpvNUe6susuXVo7zZCNBlZi+mFGpk5q1RJK6bldzV
mDTPC+8xQUF/ZPjRYbV7sVfoQKd1jMXLuN3R+aDdTw1c4ryaAnDs3VomgS5R4INS
D5inxMd6bchnTVPuxkAZ5C/rJRpwgG6zvW41Xl1V8jJOL1eLO1wfa/Y4O/TeIaNP
oLlFGadnqPumAEa95HnvOlZaFsa6wcKNFflXks50NUqKmOWr14aKdPOnmo/kM/C3
MySHwkV5Y0T3UkaMtF+iuEoa8UpW4RZCxxLPaRkBwM5nhQAKD6vX0GXms0PktRC/
8x9AT5KLvQ1Dl0d+vdXE5Lns6mYuu6ruYVVJvcYEUrA28q6krfQgsibShPdSz+Mj
4Bov0ELYN8c8FAUihSNh15io1DaYLvzcDCz3PwPCDF8VmcAyDiVJBUygeObH3F0G
Unf27VsFvV/XRFx6l+ckRDtAsCWZTrfETeJkpp2Mwvpc7cUFolAiVXj+UP10zAU1
Tb66s1FDoWQDtNeH1O3mmxTpdAEGH7t0ZpCYAzjSXBneM/jHriB5GGr3CKgxyZVP
4CbeqaVet1paFyWT9JMWZEAZXLdJ5MD2JX6H4Dm9wBsRFDFzTnnJXfubvFo0sU9c
jj5fgLPsOvCvlEMO0Qagosp4Su580WxKL3LT9efo2f3Xo2Npfu7FqOjrtqPSatvu
DDLd8Tqhop1MN6EJhBy0UqoSQG8LucIj3HZLMi7voZVPAeCunnXWrkoLCHkLsW0d
aXZy8BpC2M/AO6TZTkD+4T+0ZBgr9f+6I1KMoLONGK/dhmE8zSumk/E4TJmPFfuH
HY99bW2XVSmkva7d+TatZrnE/BQ3pztwUJoKPODWjqvYul9uQ7NnM8xf1n/5rGJP
UKN126QuZRmsi//a6k+HFFSoC0tmJgSZQhzfHV1qJuvEXjYoacrvaweiIKiPeaY2
uCStf4M624Mw9C/LBgyK5GCMhYmORN32lxrXZ/Ux1uDyUs0pfjfZo8EGYhHbEvii
Czsi+JwrBBX6vUExgjunIrzCJkuyMfKZ9axuYuOnuq6WJOqi4UFTiyy/pFbjojl9
GRhaJfJ8tPqCCoQ//26Ymehrvr46j+RhMPLLtvTdnym72BeyGewv8/M6lotGewn0
ecaG8fNu8wOfYfdBL8iqRMUYzOyosG/AJQE+xmXxeghjbZj7mPx1UQ5Xs/QjA92l
bE8mckr/Xdu7S+mR1lRM3YUINOzMY1oARBrGoevR3kL8N04EBSwg0aKcbe5Gj8u+
WAzsklEeExV7FHLlYKt+7PClvMEXkwZ6gnBVbl1PJUPOz1/FW8EHgLGiIsSupkKh
1t2Kb6Hk4SJv2hjkyHdy4IaWYKJ8IKFPKPtXdmxN61Y+AUenc4UC3DJlxKG/zPc9
SBaB2X9Mz1GXIRofFGoQv1JCG/AD1Fq13+caPWQgpQAlXVY+Es6nIPFKrZHjrQRq
wTogoCGgYB8TbMOERhFveWvYlxOPCx9/a5nrmMi7tIHzuA/XAWQNGsUvhhOHYuaJ
vyts35xGWxZV+i1H0rpIYdTVph3udzUlhrFnOW3TeJRMocpOAxl4ZhHIKgoZ84PF
BSaD4qczgBZdbv8xDSL3aaPU6+uXQsnIwaih1clHtlBvz6CRDQShVfB89739CW+2
BwY6zdaIecO0bBpOZXX+vjr9MOPcPDz3NpCvyPRpViiHUgF/sL7Vmis6QOe2EMUK
RlpFoSuOhmyfc0GwxyFDc5NuH1WzqgNvp5WPC0ZQkisgseyaYHAT5L4Groiu9f2m
5qgwcHp+HrrDT686KbA+ySfEFN1k47tj8UkBke9jEQ7FqU/XPNvySh4kVk/hEWwA
BvKM+QqRTKumt1FGiS26b+5i5t1aqDuC4cYJqja/UaIno920/k1OXYk1kXovUnxB
PxZqYcrJD4S36JAbsyY4XDalZ1+fk+pMKBUP/jJhkY6Nb55vINIBjwCdbuBVKpbH
FFsEb9gW9nyHjbt9zdrv3jFtLmjDalJRbzJhMbyHGBAWw0qZDfK3xxZis1xdM9bR
bjJDI6n63Tgk9u1MOzVXrn/O7zoXakhd0wWjf2Xxx1pzL/3PoQjGUaL8ApCLMPWP
7x/BWQNzaZ77mDiDeTZ78hKMyt7dhTxQLaBlsyhe4Vg9YlJxtqd5+ZijkUymrwWN
7m5RzJq2w+d3xhPa/gDun2svxQLfhSo3FDlYj9K1hYNf50Dlbw2Wcrf7Egt9G+5D
N2e4OXg+EL+UISCx1dLki/8Rd1w17nekKWJWJyLCkWbPo4X+13zSSPzHMf2jSh8y
2ZnoFD0ilmp5Zr8kruIGxFUudpSN39v4G5I/vDrVYAHcdEx6r+uGaF5kYuEDrkv3
r63mujlcI20D3NLGhAOhnoMHyN5j4hvte2+sbabQei5eMd4AMF4QEuvtA32wOcPf
PrXCBzPUKc17DPjkUpAga8Y7x3d1NCU2iQqJrikDyQdSlgcf4BULl37jVhqepBQH
B4bydhrpiACR4IV79T5ovJbP2PkUxMz/SQafScsaKKudWLIfMNkgooS5J7J0UNGJ
cn8UnqWEHNYxhPH/Oubskv4IlYAMLu0M/BbTapNLjzPCwQ/YaldLdp6l+VZBR6hN
I/CeM8W5nRv5LU2HxpsERpl1jcMwe8NYFY0rXImlVlyfQzrzfJL32ZydeUmCA/uR
u0iQLdbu5a7eSyF1fHylnIGOXht23b1M/GnSAUJA5FoNJzrQ5AlG6+MsbrqjkWS5
wgYrr04kKxsy0seq0x4Za54YzwmxdHae38MuLuhh+GmNOrcjlMS2AjfPLjCG9s7F
QcgbESR+fPRHVen4y4WPTF6GFGLPIrLfZG6W+YuW1geocAuQFv6XjVbfAnWsQO1z
+QjKbWIgqq7fBdAz0QGfsyAR3WbieJHlHu9cBL37XyiLpO4Vcgd46bCAIwORiVZJ
VxiC1wyYAeU4XyuXraDx/bXn3q/8LzT45mkzDKTiMo2GquF2cjv4GRoUQu/RVRyh
bAJUK0eccl+XKj+/kVe8subMIflzfFMr/rBn6krutvlz9Jra5ijnuoDkOdSmBHCH
tlngIaq2ifnfu8mRMcIpBewDVR183rG8nd//lNOi8uoAP1TtdUlxjH26hzx9Ut9z
Emp+lXS+lW0xtsbSlmBUM3EY1Qr9P+mAjnaqLyd6Nyzy6GDYTpXXoIPp3MSSuR4U
YleOGkdrr8AONPzAOjnhceAwBgcn4YVsksCQSIjyG/48evfjuwZMQZLMrX968XBI
Nm/0PhVPgN1ayvAf43pWqjYVgEDrveR0X53vuEuuOYvfMLCRfJjQbkAZEd0M6FhS
EytiPkhN9hRbHRr5hifDid1a+Mexv7klKgG5LrQw1ZX100CrCn378hGVzJXkcW/c
ZQ1qHvc36T/DsOjmoVUu7OwNbGFZEhdiv1R6A2MTn9UYcgKiWO1PpdpJtZDQzvqJ
KVaumOfu+2XCVpj2TlDmDP//srBCyYqnCVi+KL5oxZThdguspYKTnAp5F4B2I+eO
gv3rSCwSTjmNrATgfUh1Nc8t/fFNs+UltwryId/hp8rUngiPiFZQXyQ31ciijkMl
BBtKEZTEYI0iTrEOlmEuLMtiB+hcvy+TLbVNkH8eYFPjyf2zq98iKKhRuyUOzroy
O3MPlGXXU6W4Rx0fgvppokpIX4J29SuG7M7+4bhqI9Q3alt6jR5cAAyJJ6KFLhj5
wmdsye5H3RiRxGRtvyy84fAuI3zTNnjW64Y6kJDSsPDtC0SD2PKviPt5ugB2pHJi
uQPKKYZjQvBLnZTLZ2aGIpIeR3MrJEj0ZVsINWSEa8urMunLaDAanL1np25drSn9
B1pwBhNakWQcqlqo54ICcgUWA1B2Ofpns/CWmK2RWnnTdD7m/AKPCUiEDeJ1Tt5c
6w0nwspL6+A2EBAxSX1ylPXSowmrZBDGkLUkyk3kLfjtg0GSYI9efjJXszz88QvI
HKD75815mJzlr9D9Zptnp3vk0nXjp2cKj6TCtEJeCKKe/wC3bh36EahE/ZG6dbd8
Ak/07X7NCNv2edkSf9hJHuxTbarRvZg0MfdkpCQksTRH2RcnQAbOtVV3F3FYQfUR
Z9nazNyTUX5R8msIQHrRrLZPBAonxkez6ZmRvlLDsbnnyTetiwO3WzHcooH+FdfT
E49oxGu3ruvrjV+Qqb1nBmJEOM1dWnHIe7kAlKonMNPyEAeVZiIkTpC8VbgXXrnl
AzG4Zjf/2PDf/mFOPwf+ra+N6RI6cngeFQejNsXEUgcoeBAzGj19lkipeC9bkJar
u6BiuZc4R1tNrqnXhGmJ9u8J5vlt9/9mLKTB/OtdWzsv0WJaviRoQhCYqhMN2HE2
w8uWC9ot8CVUUAztuJOM7ute/pwz5+r2mCfIAD+zV6ZqTuJDhB3J+33I2FlG3TEe
terliT6LmOtOod5EYXJ5clRYXi4GeKQWPpX4HIk6DmN8oQ9D+4JSxNxpiJ5ieXVA
iHCYtaR//s8cF3CeGBHTceWbNgcgSLu3pC/xW5YwQle0gIK26sW6fTzgqQ8vyRKG
RWyzmPkfWC1loLjqTRHAOfDxATJ13aq6u4qZiYE55a1yns6fbbMJ84+OshOm6bD0
9U3PGqG49i0n+suUvKzIdNLObM6MjZb7Ei/CQ1Yr2C7e0ctWI4XSKrgHCjb3Rlq6
jBWHR39yNhlZj8mBW3qVchdXsQPZNWZp5Scbw41cYlOC3ZNh05IvV2yjw0tHnvUH
AIjNnFs7LkpkFpXIWotYWWMMzzVdTkteE9UYoOB0gQ0268nReNtWyk49hvMT9Gfi
svXPoTXjWmItu3tv6JvPTAZG7nP8Gl2t3ue/nqqsBgyeqszVN0yn99hnJWrO9ru7
C/PdxkqwXWZGjA//2zpJZgue9DVncMiKLMUHwjJpvEG3wYI8URcpCkY9OJwcBEu/
RnHDJkRsYs8Edu/Ge8ykPHnA7ArVEsXe8xSY0cAyE+/5WKvEjaaLR3S24ZGma5eP
NsUufVz5750uoCXnUwlmQSa8g08Lx2K5RB2HU534TQQbe87+S7dlBVySubtDYVyM
DB9gbyR1V5GzlFh1dNgtsj0/9RwEI5+L6m59JXEQhOLAAYBUVwTFDC9usAChNoiZ
w6ZtjEhwtlAU/qxJ4KHh5aoNuzG845+QNTDnfg+mZg5XffX+hcnmDAU7YbRjylNg
7hycYEkRxg3/Oqh/ULYDHlopm+DJPIegt6fGryqtfnOe2IqyHolzgYrt3mUFQ+Eh
qGQWCli3RLFcDX9RbQ7LB+SB2RdgyXzCyO0GHKDg0DEUjo9YJyVJEzKiJU/klDYM
bRrCIurydgC+eLjnh+vOk6vZErm6WOMYHT6+7GVuVV3yzV3I2Uyt+JYzC/nrVCwj
DyFM5PBDu8cHgsbHRtwPOoXD4SB1A3zDdWGeKK/NS0G4WMiWYr7hmssuolNhotUY
STjoRVmrv93HRum4ctr1+HqqWD0dAdDs1MMikVfn/gDCFD6XZ/f0WA25QTplSW1G
WFmwALqZOjb3/30IG5CyS9R8HeRTAljBJAvystqraVcfwcnKcT+IrT3W/AFv5kkV
Fo+zt9QhdZyv4xpEq0NPIMZ0sjKbT2Q6npK6iPpcvibVcdDqZU7k2X1IZ0SJimCJ
bntswGgpIR4Dg13dbXNhrxsJeEXlS7tEF73ftl8pVJkiwDXH31zeRKdvm9AnFWmv
zUwOoNrcgVZ33mnvNFujWpl35cm8XZRz6FIlDxDG05NTm7/4E9NVwf3QTUua7nbk
cyWz2gCmqoyXz/SeKEbBj08HzmMrEeXrkGDmRX2JwVt4MTZ08sExJykYJQJANXXZ
At2bnMQPJofsvCjphP9GrIPHSaFc8YHKpmIBMtdXDRwmy64axr8AOLIPJaDvHwSK
UbOawaE2gg7Ym9aH0S1LUBOFtbhZ3L4+/RAGHUXF8H/XBU8cULfu6fTJQGN7S5N5
BQUydSZ3HFz8pnIdx9jlDd2gEnZMzPhOYbYcYAg0ToHRC0b0s0uHGWsi+yGRyGBD
UAKKyLPkvCSJn3+3Z5W+nBzKToWuxtbX6c6s4fXa3B8lEL5+79rrkma1UDjPYsx+
+Wh+y6qs/hXXyS5TKsXTgjFPvm0++W+pFQ/rb2AVOtEP6V9We9RAHSkMM3bqofkr
jEpJyzNJuNU9UHRU0BEOgE1U5RRhVNjuD5J2VIhpksxy8oC7hqk5JqESDMk2W13D
WS697BzPFkHXMJDXoXCxdcC5q4n6BQ3t+lT647Eok/jB1Y52MuoSZ7wtPyV/ZY0p
2u3M7W2G+8W1a3TyWyzKLGk+zdu6nxbWmYhwoMA9IJhVZtsTMdpDdTdLA7bMlTau
H0sMV8XQy2CXuQYfIdR07xrm3vdhWcTnBoELhZmFI1nLb7t/Y1J14TV87WUls/MY
zKMippSAAMtuXS7iRWVA0JaLxqUvrbrX4KdhdGVDZSzRLQWYOggzcC05sBa3jLme
BR9dqrAThnmVyjzI3z5O535+3Y0OQRznR9Umm32c8x4Bk9WAvSnhBx/rOdJmw/HH
fW6hAWIWPysnqk7npxE87GhbFGyglaKhRZQFdhRkps0NdMPUNWioc0SaFtIcqgXv
QUzeJ5wk4gtT3gt8/4TPkD6sJRHOeBSnAgvK1GYftsP32+wy1yJDCLbIXzLWCbEc
rHpY+uFXheXGNAanm/a6ySvWg8zQwMigwwmQ9S/z/zZMpjyfAM39gqqJ+WVVl5zg
CQrHvn9avwEFT15zXVEm7LhUjI+yil4F35I4cRWrAccWizv4wZmp14+jZLhQHT4z
Rrofv5oAlEwn0TztL7Bmohyz/7FMGYq0PLPn37vVORNTA2HBzYx6Cfqmfad6Fl+r
y6UaO+jELEqsaWvd/ShfK8Uvnpr9DaotNJY7joxGJWeOls+wyx2Dgj9U6ssOQtv7
t4btiAiSGwbcKjjFsPPNrnwlEj7OfqcgyOEzpqHbhHVShTqgzHjllW/WAiwEsD9N
f3L4c+bP5jaZigqElV0iPXRBKnaWbCwANdqYPWOHJbD9U5f/dVjCyj38km/Tl8cO
mBBTu4ftJAgruF7+DDNiDnpl3YNKiRyejkxjxRAKrGL4vkB/Dw9AEWjAkfOebFph
ug0zGoFNnoFMrZ9gLJc5YDjheKAofQ4ZjdpCZqxEN7tEA+kweio/NexGOnMi313F
cQ8aNEXNyNteN6BBjuECYZWnAomJmOrw0EpZrr9yTq3k8etfPPyZZrQXoPIvMXOb
z483nf608PwNz4KT2X3fqcIshHGsPAAQ7X9XjqAh5qc26EC+pbCI6QHXZucGR/2x
6nwRgLTlgefPwj1DTKpsBj3IC7cymJUBekCoG5+T+Qwf0dZdu8yb38H71UEU7aAe
uQXZX/Rvc6yBG+53MOqfNVPg7jjVb7tTlLeaEPl+l3vVK1CTBZeBLiFpK0ST/4eK
gyIVvo8DFpOE3A+gdrwvzOfbwOvHK0cu4uAAodLlxGm5un4tDK1v4TSWoaUH/GKT
xula6hTICpgjanPDw+CyN0TmirlItUsbCJf3Ug8cGucviYR5PG25qOe3UNu4VVCO
PHMkKBTWyGw0qRLfZxb3OgXK+aZPsEIo9KGQzKLLsfvtH9Je4hPx8wkupGf2Fz4t
h2W6Z8ILcxSXiXD4iuoHfJTEtEN1+D8DQYpKOLWUofR4+G1vtnRdkVqbLz57cpUl
uTvHsaRGYfNu8H/xZsG4mlrKPupdNefjiVpwPbfOwgo9NGPHvpSaSTvysWY3bd86
Zn8wgOmO1Adrf65fkXEUrTmZ6hz53Foj1OKrOXogU34akoUMoAaqy2yIVqWPLg31
0dgLYc4VYn2rrIPSQcvzch8suYo0cbvvDQwy4WFtinnDRPSsGXJCvSATEJntXnMI
RTWNVS6BZZ+W14wT6ub3VNvfrQF0Zq3o79guEUTJBzgTfa0E8lIK2GOh9pVXQMSp
d8SncQE2E9M4irB4ctnYkQTH6zMEJJNugg4zZUvT8+4RVQbW5UkdxWDnPRRnX4s4
5CKftwibuZoPl9WCz2771MP8g8XZSY/TmWf0mnGegTpTYjkzofxiP/dBgtU7n8aA
e5CaTqcwuCePiwH1lNwI5MBrXJed3a45KlRarao0eNzYU8eORxouqOV3CC7f6Jmj
FTJXZSDviV4KWIy+USQ/wRmChTeLGKaRpPC6Fa5/mCFs1QVEr8/UPPcVkEziZPDO
qdCBzaycJNVKaVAwFkfh+3OgjH2vZMwdgz/hcfW1KYmxZNkCq66jEssbE5fECkV5
p8aTCmwl61gVs0A8W0Z49Ujou3b5WDTN+JAUXCiMae6BEjLoP6fFt6ZRV9Jx+fk5
qVuEpybB3jPXLKJ1avqJZhZfoZc/rU4r01JtTa7BurSbnGRATQplZWQZztfFDo3T
A1sWXfLZYuXJTEPtEgWwYcloxJc0NXvgT/RRjiiZESeYONPJQIZgnyEJAqgjFsYL
9GlJsr7RZj07cJEw/l/hUyEPsqq8nwA2fhaIi1WQKA6rRnX1kQuLf20SYz8chX8f
hB9bS/w3urTsm3sK9RoTS2+b90QtvBCMEECrSaR+Z+/tXIvnVkotVlnCxaAlF5JT
RHQnIsiqlkQ1BdMVRmLDrlOVfMtLTWwQo4RDZybQ8LBL692IBv1USlFH+sFJ3tZQ
z1yReF/YEgl/5witnWVP6Bl9+F5wlYENVBAIaUUWDDvPbc01qYjc4MqXC8HuwCHM
kjOY3SG2KtWApyxF+aIcjkdvGHpA87lstnSPRF6ho2zJ36ww4L9CvO0WnBSSVY6e
pvVTlsDbTG9VKMWbf9DBjrasSsq7txDPYWYJeEMSjgbta9/pEG1E08XRKsTg1fc1
8BUA+OTFuuxjKcdFHipvxNE23QC+z2AlWeZrfURA9leXESbLB71f5rYDUhADDbR8
IwubmAv0BNk6vYduyRIRN99mfF/zIVKmtjTk8Kj8ZrARTncpZzeDqF32bfKQG6/b
9J0hlaSTY/sc6XRpUP5mlL0CKTV3j9jCQFomZwQd13iE5w9WW19ChYg3+Gg5eBFl
TlmxEIy6ZDqsoL4iVh1VxwOuSFAXS1Vm9/9cQfo1iPggRoH9utJLT6F9QrAluo3U
oCuOOFHBb7hcSBXU5SOQmtLgrulPMC8E5PskgPGTqcM/UOeifiPsqhp9yQczsMJm
SSddGsFPbFYvJWUPCtR/xwCwkS//X2ZB0g45fbKIzTQIBqdgS61O3LmGdvn1ycZW
Ded42DZjnEoPm1jC9cgsn2UnBbm5k0f1l7GjJnPC4rpeNBSjpSXd34H6Nwywlhy4
beWcZBzwoMRgorTPB/usSgkp9MUyivI/kBo/a+cp0kpZ8a+GERiXaDTmxGQzMYqI
BPDvzV4nWRAz+hQzhyAANzekCMFrIOs0Okn5jv2bhis4sCvURBWxAmNntu5GqTjK
tZ+T449m69YRHmLT5+62Q395qWIbqEkRFb9eEO550WZv8UP2sCnssSuQ7BXTZfiy
MOOvOh2IV8SpupXLeMgNp+AwS/omyQyTSUQCMUrIzF9NIr5tNdt4q5GC61Fu0eEy
AvRG1jTYmDH9peHrBIfR/7du9qwvEN3QJx5a5X0qdlpiDYawx17CzdsTvW7tJKiM
H7SLhcBuFtk2r/vGxh2WnendZBt4dw/l27QquaBrK0rGEKe3cbQuYZmpNq+XOiSm
kuLrfpMVb0reTk35y0pVBfVCTYfMHnqKIcXxZKtD8yl5J3fvPvhAFzWXGlOl0Rxh
EPYyr02LObd90xRVUTDjBN1ODdXNjYmDW9lBYNnifrsDi7tEdnoybPrWY55wYo6/
398IHpaOItJ3W+v8Zo4NKAAnYF6rFEwW5PLCLzdmCEHtJBOcMxiGJvj/XkMwCCR/
6tqmMqU6O34nXHCai1y0ij/Qd3zhfS3I1PumynlFPZS1qpAw9wsrjaPnA8JToj9+
iLXvPqWCxVpdTMogrHOyfL80c6NNUvZ8O353B9v0//wIv5gFCYkwk2nX3oB46uie
rsiEXsugCLVxm09BjJIvhR4AcRrl4/aPMy/K5E9MpwiMLC4sBJvp9Jqt51oOF2X4
qUZfErclvZ2rkSnrgcfRl215fJQc7sg7AGd9IxgGEbnHjEHr79Rr28f35gXSOvB/
5CUGB3f6F8RyRCeg9Or2iqga1+j+fkVb5s3An26AlVa2ozNEYpaVcLUiaSlT1Tts
vk3yvckl26if/OyvjP9vizhlFEPpWPVIvrX009I0ZcdTAOCXfWz34Yy2cBQplKKQ
X+uwbsrXbVJ0LUeR2ZuqKvVKEt9AYs7Y0K400dacf4KuQdOwH6V6qVSyGVfhwdqm
1VINozTYrHeGhyhB5MOIrg9ZjH5RHbY6ev8Pj5mzWns21eDuolXXENTyVcm6AUY6
iR+GMWKCC801Il0RIhqcOS7lueJhwBVvJSA5gROysql5C3frVCWt6tcRT7shUpEs
oUTsBbs8OwAkB+M6Ubfz9J4hrLteKLjNufUgfMiXqKpcLFCBDSM3YMs2bSUBFUTL
9ASniVonS0j2IygbM0tgv1pZJzOOsDpkawzjVueDXpjMeGpJptdjG+7R944aXWr5
Xd4xuaPabPjy/aA+nFGsjqpEckATxB7GT/iwFSSVp3y4oPuhCZWw/tCF4yUvikGP
RCxLL/ti9cheDumH7wa3AVxX0JELNWc0fJzwXQ8XxPGw+UpB/xfQVoUlGo/OorHe
rMz1aQARMM25uiNTvxJLO/BdXnYPsAh0eGj7eEGP8+Yj3NwpOkZx7RBRUp9ovuul
hOVhNOtzIy8mTUKhNqVxhfq3zwm8fuxx3THeweM415vxDt6TiIS2sqWyaZrcrhBn
zow3m+J0x0/KQ/obvsPKSuuyu5sqlx56OEv32HksL18MSxiQCIyM8ORqeqJS6MFd
M+ZYauFRfhRosoYU4jBaoJywjCjBKpmsmLWRpjreC7tv687qxv4HXNlheBCd8I8w
PwY9OSZXKiVPAtPJN15uSVn2c/2vhdFHk4JVtiZy4jziNUhV2yG5+uHiQFvjcZAW
oQzzapV75ZhIidOUe+J7itHoVA6ukzM3VCrXRiPKdMLEMI8aRdtjIiWGuwgf/mgZ
imtsdGpurkjcTF/wb1PMDe0AI1L7vKU+j3PDRvCwCpK/dHDWuuQNdvMy/zRJon5i
vCl2kgQezFlfapdUBYS95Scuz6VVuD+KtRuFmROWwSY+gE3krLDc5W0V7QLueGK9
AyZnY2W/K5s0GoV6Ky4Rn+lVOawU51rAml8hB4nRFrAqJw4SxzJlier5RofWlAg+
vyTP7xaRT1+y8lOUNodpJ2757dsym+L8vVMe1t0QUchZd9yA/QLstqgY+4HDcAie
R9aMmhrV0KgXg63GzDjSMp/AK9zsqnKlEQveTph1ngZjnzBI7Fhrwi466eDXO+TF
GBQa8qh/HolQpUcMTs9iWQ==
`protect END_PROTECTED
