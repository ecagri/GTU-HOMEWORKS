`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PxtvejQCd2qkerQmswMqsaJDvo57YtCKqo7KCxy6GWTV9+dtE9LgBuvgTqfcLa1z
LOg5GSGYXyhSqQa9A5lz6t6jibYw6dU6Jw7SYdFdKnwhCu/Mkk+WeELvgs1HxRYE
QuiRsbaMFhqvg+HFuSUTVCmjsHJBKe/clhp8kprX00P4tBzeN8RWuNKguE5L7qiS
lRWeDC9U0u8ZQPCd4drG69jEIQNuv7U2g5m05bFJ6yKIhg4LvEfQbGoHR6kykpN/
0WrIt6/Q0/Ud0z9h8uhSbbAEzQWsjyNqbv1hEJSyvwwLuVkiKgZi61rHnoRJ2iZG
2helzy4Gu/qi59jRy+Gc2jnReDXSsECT/NmApkkpJbho6oc9oP1sqhlIwU2m7otA
Xj2qCurtEpV6VHmc5F9Zv9xL9Qan7O49gNJOjeHuIQQp3Yr28D+X8rXRsx/ckOoW
ilfNGRcr7iJ/33jlrdVU7CkLOEvDi5ULzQAUtEJ5bF2h6HkplfhlkqmCPqV645Ua
ywuU9hcSxg5zR2YHQGiebTGePkm/0HYnXRTdOuQiEBD9D+l7CezdcglSPZeuzz6F
G7gFBYX6FiGpzXW7LOzKIsmQ8stU81y4xK8ifR72FQNYN4MkRXPB3gR/tvp0jdMW
tQEzweo+EYeWGzPSkogVZwUXg3F14NZExkNmB7ZyC9K53DbXIDA2Ii62+k406cLd
+f5OILvLxWArPw0FlOFJoLycnj+8wQH3Vfj/naLXchb6/Vx2FAR/LRq/HN/Wh3iz
hcEqQ562frJIFlwGljxV7CxdJQT3RrS9znZ2Jr5Fist7SWEiHn+dj63H5KUELYR8
lhfQWDHllDYxuBWN4LI3jo0OmPalhjaQcLEvM4ZH/cwJKAsFtwZFnbun4EFmIWtu
9ZHarGmnOyfaHdyUZA+KRw==
`protect END_PROTECTED
