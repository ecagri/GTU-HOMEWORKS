`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rad3YApoao5L7LgpGAEoejvSQ5W35BEsHAjXsS427jva5TOFHFcC4FQIxFAvtsQk
E1ZW+3iSccgKytGPjjDQdZCzNUIGU9GpXVdWCQOBAULInBDeSrnyIPiw3G19jhY0
jNsXALzcDT1Id4FIM/Xq16m3DYNwZGzcxtkNeV/DjVF4K4Ur/WZ5o0V7ioowrUwZ
ztBx0MfkaYa6FqRPG1gX/fapBAfqGDP2BmoRA8uqY05oBL12qDh4+CIou5tIhUMJ
pvZxiVA/KAM/kefaM7yONgncsv+m8FRq+S+prTgZP5EyoAcSEXknSaxyjKJ1pM3+
DJ5Rzja+XgCp2wm8X/XYMPUhlnGyi9OzuHWnKcZ1uncUfSyd6rsilWNe2XGRFgNp
HPQKJ9cNM3IRqtK4ev7caDhWDtNY38gW2drHdrDDTU+aZMqvvZQP/bLlG7a3opDJ
KpvkJsVC8fsjXVNUe9aoEP3XeUo1P045wW6deXcjjqju2EZ3VXn56EqV3fa/R+97
12MFmmppaBwi61HwvjtQlq9nV3h6XrGuNoL/xf9HdJjDwvzrnH/bpkbuCdG141uG
mPUS2RnpbSgnXLuYL4TNcHuGl9tkcoMrKSfslTJohrfZ49y64DXII4lYDd41Skwz
uDejl7PIpQg6iZQth6H5hULktyOsRUi+1Bvy07g0Qmi01Z4IL0XpHAIKd0VoY5A8
cURKAMBgyCh9+Ips7b73kYlg/Wi8zrzR/+EtdLnbJUDuuwhxnLRyu9Xw/1uAEDRY
BzwjAvzY6BMiYAXw7GPh0fhADLYiiHKK8k4/Yrf/LMKbyvLYxc/wBYs0oURzxm78
JcTzZNpxc0qXwBYuSrY3X7WyUZ270R8xixaEWjZyb/vhPHAdRO9zeh8nU/sHvp3L
1jrw9hxwofXXpRV+jNdAMOHFKMpBmc4LtWc4/jkzy5++iIiaAbiXzx14IZ6oL0wL
UiJCvCAPEh8D6QzAJztBB2BtZ96+VMCesSXlT/uKTea3pjuwqKbCUhsNUOHvbbZQ
HiFJFLE1Pthom3fQMLAhSpf3iEmduCESH+eYmh3DbAR6LBcxk4y/Gf1DQBVViaxD
GhzkS0K9dfU5fYX5Z4xNrT9yl+Ok0+zbUvqt/EzuJB6wnAFOv9QLZQUQd/cOHzGi
opM3LbQ+56rZDYKwcavg42a2y3zOhe6BMOswVXDdilC8rc4BT1SVHK29/V/IhRBU
hRINiXhm3zWheTPcCRfTDOWnh58r6AzgLnmQ04CEZQOLpQW6YSb1lfBU+rMg7OZO
BifOCPE29Eulej/QU65FYRPFv+rhPbfAjgHXozpO2UlaJSLEfoP5PFG+3jqCD0WZ
jy9FuYK9V+NiVF1APrDaIxiWcMpi9jvi1IO/hwh9f2q77zJTqXa3XqEWHBHD66wA
HGFXnrJ4HtfcUnbjUtZ0GJGv929BDMPCwyZtiSY5vkgkBr5+zId3qTRMuqYgYmUq
J+Hu9GvfTWrjosKU4hQcWSLXvVic5UnKP3DjTh5UKh4fHHwNNTZ64JkXT6eBRSX7
S9RtBibbuOzmLsuzZ6uV282uJXpq/E0E9LcENmRIt1o/S/fsXp7V/wAFtKc4ueDb
0o2d2arVyHWPZC5s33cb2kEBr/KIbTfxus1dnej9KNkLB+bXQlTA8Sc4zIb2dono
DQV87w9smbP4OjJvw4wEyFpGyzMhRUABiY4DcN7T6p6mCBaPzVgU5LsOY/usL2Zi
RCBkpcxPEPDUDhTpued3jhNosHJ483thIJGHZpWf1IXGrxlED4zjDhs/V5JxEZxP
iWVxSMhtK0RIrMpwbNuva1vsJTWKGh7wYCC6Pivn4XkUVgK0ZTXBQGY7/TVhxf/Y
djUyfClUXG4tzywAvNhm0j+rVwAT4+vEoY+SYUcLlJLEGjqc9ddwTilZP11IYnHL
Ed2PsP/XYeaGQ1pe6hH5aAzLcXKBxdG0uZbYvd7C91NmGQzOHeHsyXGAxsSyABJs
aXW4LKWX89y9cq/JZtq114CQI1nTAWmsiFKXUwy+frF0jSDaPlsiYWEn2QNdUwIL
KOXO6ZKk5ycNqHZ9/TXR0TVLpTott/sRh8JRW6wi3X5Mj8bpvcnx3cpPclhbdpSL
v8Uuw8G/aRpKD3xzKi9kEn+XQ7wKyqOo+iMmX0bpFxD4DRB89706WuVHX4J3s30C
b/9Co/33pUCGpe+6K38It4Ww2c4luD2NPC5LS5qupV2V4MwxAqkD6fTIv+oncHaF
pGPLMo12izk5CttYs33iKpZWqTaciunvTqzGjLBOg9KX4pWJAYMlnTyqaoA071c6
iw+qeJLegs3Cg6/NO5pv3HRcQZ86DIxn7pZsmfdxBI97/TiOyo8Cq9bnuIxfC6id
qZoBIl2q/EUknBKcbjmhyfBb8RW4q6o91VkWH6vqWdyJVjyXtG4szLtIZVDmEKFv
FZf2bmh9eMwh1w84zczUbnwlC8eEoMhMFPE5hTnmumcqMpieRiAyn81JfGA4IiW4
nt6utGpfunEgBaN1u3eVVSZUpruHdRX84xiQbaReJkpCTWQ5lhepwSviWXXTgPn8
heAjC7AEPWeWXaxnMyqhpyXQF7sK2QrWR3lYVhs+sTzvN2LG2fWEeT/Ki6j+5Al4
rPIBbt4WsI5KTGlieNR1ef5TWz2cx3fQk6rI37viVoiOpNG7c8dWP2kps10xQ9Ow
r+4bEuWzES56JlpuhpHwrRHYUx+XBpjcH3REhg4/ZHpFDlZc/re2PNj6wvL3KoOk
SSvDb+YxhIyf9tfh/pB0RALnJtg/JunFxioEIyyQdUU7uuN5b9NUqglxJJLxNAkx
dpqavYTgT1TiYVXn/DSNVDH45ykPgXMLqolCJuPim/Dykdc8lOGeoWUQdg9Jzzrc
x+qY1d83GoLI78lJWT98TQwEepJFjYmOQ7SWKaBQ1Mg/W/BDc85jbJ5n/WAuDSwQ
/ZVfVj+DwEj8fCqhsMOTyZ4E8Q5Lw7PcCs4Truzc/lp4761VDsfjfuzL+2U+JIui
JWQ7emM9U3m/WI8hJX/CrOHgKPtjxkfLsqz6hxVmNIAfnre/w7GOhgzS59BZF4JA
8m2xm5KyUxFlGmw0fwuX/n/sT865fA3yeE3EgKb45XLx/eewDBItD7AtTY7ybKAP
jBZuoK9iraSD0A9HtgesEgM6+hDqnpqaZNV8UjlJAryirAmbLpN3PqmnBq/reDHF
2OMFzB7dtZ3Nz+4hAwBdKJ/J6Tx0DQF+IVqpdH2PLlywkvVYPJcClEvMVEAkBJV3
ZRv44O5X6/M2CKKRmlnQLeNUPDbkm6kFZ53IMOeuxmTEaLWMbPS32tGEVY+ev89F
SIN2OnjcBQioTkWDNLXhamvhY1crdOxjVDA0dCZGldt+UcKxRtphu/tdO+OD/ASq
YSq7kl4i6lNL0UgkTouBBMj7ereXcsMyOaKbUlJT02MvFqHz4cakTuEGLyD5Dho1
PISysi6qW1YxGRNScs8odAhb+nrno9GgbF6T22Hrg1EoGjwg9jQSZAGuFbOkMTxH
YLp9JF1CI04zIu9TVe6N7gsUYFxwe3FbtkP5KdOjTSSHOkfu9SklG+XUsZnxBx8n
JsqIfpTC8uP0qx5Y4cmygw6/gxFJy41rbrAPJ+8RDh5tq0thI46oKwBNZa+3BwRk
miXPq5vBPDjIl4NLiHWtNQi9Fz9iOBwgGB0fFkNOVII9/c5mhazgoNoQkACXwfq3
RRldi8/Vi3uidq4JZZIHx/R6slT51WbPYsyn+x6Jb8gDPBQZe6xNrPMa7Fst16zr
zjlkRFaQIhTCjQgMJY2qU7T/IJgymNlvD6eyWbN0DTzssNwPBLWHCcaZcOngf/wp
wC/JIHyrjGL7XCB3L3QQQ7vL0rzqQXYgZ9yJTV6ppevO+vKI4h5Nnw6QotkNojOD
exdlmFjZGSo3amcKX5nZBA+F/pioN3bThL2HrVQKiD5s/MYydP9jIponoi5sMSmq
z0x/e12HvsykL7YAYEIjoE4I8naZ8qefNWYWn12Ofoq/h/el04iim6WlqGzRqL4B
0Y7todEd5mEC3IksHAgpYs12CjvoIIGwQIsZUWG0IqaZxMoSE+eFidHstSX5znQR
GVb+aFEVmj2f+zhANUErbpksDDI3ovYKJt6wtVEWiC6nWbmhFZYLn1uXi/K+zifA
7TEIGFMBUIdS27bmKyljkUEENvCJzFmw3nPMiol++/1x5uZwX5E/v1w5493c7Fk7
LfjhJxlLxWhRqOMQ+l8xc8sQ9b+sBAMusjfUaLj8QPeWsH2xXAIHMPIieBOX2Fz0
/BDpQFbcX9crGqo1311MyzoFe0gduSWUqH2sX1PvB8ky4BFJmcXNLakgNJo7ZkXV
r9Xymb8V8Hd0lZy5zgvGhahl4v5GIAxvWxy8WFI6nYrp5hqpc0nn6hSLACTpWK1B
yS4XeNhlixrpY5EWrg0buMUj++wHo/jSqZQChEEmrNFHYupr+YuD/ZNkSCjGWav2
n58vyziQw55PqFm01ie5NOSW3Feznv0GSCp04inE6lbg901JbzxvBUloBiD5ghRe
eJtK6G2IlusdJEejmW2Bi6Rovh/2YlrZm045DkKed42mzpNgpYyX8eKCQbus+S39
AJOcGr5gabhn+fKkfUb3pKmgvPvtM2oRyJ/lavkcQdeyuO3K04B65iqnFyBcrGC9
qyvZ7YbhHwdqvc0kN1WXz2d+rG7JFlqO40etIGlOZfutEz97OYtvnlST7/bT5Dxi
zqd8HbeiXKW63LCR4zoXZJLMsCUptBS/b47TCfMUPQqwRtE6hnhHWnyXszwT+7+h
sT9Jm832kj0rmT85J7oScGNDtHORpGUFqHXOv1C8jshtvrUf105pI1cZrTvanjAA
mhSHj3EZESye4O8LCvMyhT94bwWt5yECO+UhArbA8kg7yWdiVg4GDpbisrUHgSE/
dnv6R1zXIvmLMLuuHimQmAHif3LWfIDu7G0aqDLSS2RRlUzeB9CmQUCk331TxVhK
m2aQDtP1/CObXnpCu//i3gD/JQgkFUAvJ1G8SDLcVZuMIIPwxA/9j3rZM0tdwYvo
xtTpAq/PV1M0UkhgNPsy3fHEvTmviTz36eaHm/No8XBs6x6R/cRfRvvGHW5Jb5+n
Fvd08kCMjKwTbMOxl5hlNSLkZZalyH1SPP5wUk8qT3uOgQUaJuPnRqBPy+RhHsAG
3gX+/HXsT9RylSgNIOtgW7QGbKncBtOiE61tmjrVCv3mMPoiP0HVAHTgSKcJ4AH7
JfhT0zwvhecelGho4RHpz+ASAuCDbe5nSITE9zvqwCn4lo5KFDAdLQtqj78zW8Ou
LFr4j8O5EaRL/JmGdjwXSt96SYfbeWWPNDrURJbC+UcR1SXZkgsuYjoa3tM4ZhxT
RJPypW+Mif8tgyjqSDR5Fmzneo3rjziGJ5JYEdzJnucwYirJR3FlqVEUe0Cbjw3E
mlUHsoKnaSvCW7ZeE6ZR6G4mjqNhhOAMwwwqfMZyGf4if9EmjJK56YIiqZXt0asA
3c9fxiFl2tVM34MVLSaae2OBOCAblxnZqIzgRW0PamTAXNqBy8B1bChOU4aOy7Eb
I4iRrb8PKcYwi+AIgQrii7KPqj2vjGPZZ3yB+N8+xNb0PyQP740zi1+KYnxjxOh1
oyTdQAdcEQmbWYHfHt2FKr27jPvnG5av1tGGssnCakcwoD/IVn0ZRMp8l65hfMLB
knNeN+/IfqVY7mHBMwx7BQReJrOIVzRWO1sXWG6XZfclxebTSaTbB+82w98V0TQi
b7Qf5W0tcjpTHy4MOqXH3yLa/eokUUvKvEd3SAUbXYLwvfDMdzl1ZDa8aDiZT8Vv
6+47qSkhKJD7ax4mme2m07eNCklvOIpD+ekJxLohYzGH3AOhvGVXuQSTZH1hSVru
MPLVLxmAZRpmrIInlOAmBDz1HGFvSiuBlBzrxWSYc47jcUc1y78c5yfXTFSeVL2m
1sttpYQC0d8ijRPlbEx28V9SgI8/r3xF2CCCcf//b1jeJVH9TRxRcT0IibbXAzzt
9fexPQ6RcdHe2teENeC/0eufUfZi1ZSkafwLv5V5IWrpEllUMjEFqUGcRBQopiuI
J60JVTl3E7kd0Af7ZvnaFVYja2encu/kxgZUH3kYRrkJrdBwJYc6+h6CqIX3+16J
LrEDktjnH8iUmmFDkicKIQ5ZCeqAUlxQms/vBznAa7PhnOkg6fSy94mR7+nOU52L
MJ7xlHIFrJpDNQvmxj6JosRNNpUC6uZWOxDUunNJZNDdBLJD6Q7nhEVO7YM3hNca
jGGdVUqfSegdIWdKJ4FqBRVNYWc/J8YdP2IAIdn+c0VcaOnEqIpy2w8DJmJx7TQk
xkhWDrH+pfzhk0NkN8OkR/sIyQ601dUVe+OCknujgHO1HydkxUATG04RMt96dPCA
JFtqLjvBLyWannukHRk1TZl9bQMdlelb9INAMvPX0QtHgw47jVKnebvUBfDHphRl
8my042o0EipXtOLBKIMv3nLN7Qg7Z1m2kOCAPGGW0ewmPnsNgs58+4V5YQAnhEzh
tQXo5tJ0n8s4hiw8l7rtMni4dZOcbKpKgHfM3lDfU0DjOy1mBpRqlhdyezAOmKax
utP0seN1XUI1gdrR/trz42HGt86KZoarlISIOZ+WeS8vKmvPi7HWARohKQ5TbUHa
ieZ2XDps7dJPrfV8gc9Y/6Z2mcXyeMJBgsouX9JbIjsr1CrZLh2mqrl6BoSqShhq
P1y4OIzGSJwYN1VGF+jTkbsttzT5QgPAKysVhIsuO05bc7r3U4jzG/MJv+pGcgqV
cTdfHU6C2K1TMsoKbRmVOVXe6XKATygBPGLHBLieJOkhE38c0XKlsWjbj5glGtAz
gN4IAq/v3SuPlAfx390fyKzstcQJ2GlM1zSQM0rNZfcT0M7PIxIO/GPYOH3Vprbm
sjicFh4INXA2LlaJ6fq2nMfSD43FpHKJMcruCqJaVjDb/QDNOQHASDJW0QPzi+k7
xQ82khzdcm9oB+gWUWD/F10vOYbd9X6bNfniDCLjP3qEe4+CLIDdmqWA0xjU7Agc
I7dDK35/BatSDPTsMmQupZZJ9pN4C6NwQ9TDgLwAb21qX+JzQfj3HKv1F8d4dNnE
Sk9NagYycWJWyUW8DWgJpxEj08/2HMEHextSrZGq2XTsRZORSkcsQUBPpxAtPzAL
K7h72CFrMRB59lxKpYtobq4YjyH29R2qCFGehdMgDxg+nS4twX3iKi4w9dogl2kZ
1zHnwKDeDua2eAVLUnmr4V2pl/+RoIPnq0Dxtnk1vbiPOkQ01avbaWLFTbcxJvzM
Jo6gLjkpA96gq96RidJvyNjbsbIqsRLl1e7oOlJAE9rhcNp/qhLF8rmz8ZJuL/ci
9kkXEr/qcSePmzT3T+RwEUF9HvtGWF3k2ZvEeqXqD6GBk3t8YFJwUqzsCrYNu7qU
xZ4CmUmGqiomfht/1O5dT5mfUAtFWPKkTZvCaRriQGoWrgn0eh5Mr0vlZd9UOg2D
b8ZIOiMUK1gGj1PzZTQE/Q08WI71jQ9SnCgbDQ+NM4F1UWNvTH+XIa1IZgudDC8V
cULCgq34fU5cK2Q8TTHtKiDvyTPqPUfxYQE4jyGHMmwGW3uK/7n/zPNPrnHgAs6l
BVpqTk0pX5pEfL3yzIbqKMJ44SVBS7/7txmkJe1r3mk+3g2x/TeIe9dI2XfxcGJS
wxNY++Mq0L6fWg6ogkD/LFYnw/3KlZ3GMPIiz9smMWCR2yWh7mA40TTizh0dD73H
X8ynCjuWMak+735zNpBimrESK8EaD52KtlDcJ6DHaMU4Gi38P5zQCmYiZIB9BxBw
yLNuMrdRPAPOATV0jdSfzt7JTJ7x9JwRtwU7LhpqTa3vCUkwTi+ZGCE//NCg7Q6O
esi08uwNKJ3BIC2WZ48lF0f95Lu3/nuzs2Ax+lXXfyN5OmsDWNgcBYaVIH7UC9N0
2W7Ekts7BokSTuRfRMmf6fv3FECUdxn70hZ1j6X1K5Sd/xL6MmTfj1YbtgCxPXSg
ey5qIIzBkNJZdR9/zOlxNyLPc5i99bgLvQ4fySTwee9mY9OxARTfNw+WhDj4RvRo
IZ/HaPRZfg96OIstjfBS4uol/a5cAdhxBf4TfAV0Mw1EySby1Z64md9Xb9hmPasA
2E236V/EwQLc+kT8uo6LZSnn/4kQIux/A+y1/0p++sn1S64pj/odh/9cBIyL8LWb
iB6anTQSdOO7cxEhPnaqH1V+wyIUv7oYgttkBG5ia//pXAECexvr0vfoi7tPskdx
JpNLbC325g4tnEIAL6UoV5i9Qp0U0GoSF5AiyuGn1hLrAonLOcYnSmqB2gyujjgj
vTFipqYelXAkXEJ/ximZOm5wMgOv9qfoePw1thwvQ8pLzPAGG5p4v9LLaZW/QhWp
u1jyD+i/Ea23yNFnlM+vKyzHnBRIRyEa/cvyIC2TiSfbkkEQ4wnjiuITefh9QU67
lewzt/H85vxGq5msPus3/97tvzfL7so9Ve30UIDs7WMK/BZYjleQHtMwdGjpF9Pq
Gj6uPQRvfcWIXvNV2DyFsLZT9HjTHGCDrkVETdmLV4hXl16pOc3qy9W6XGRXra3w
EZiA1Pg5wQxjpewIipc2sUgxehSZLRBPG0nmSl+Ipcfa2icUwzkfsHYnoAqz+Ht/
efVQZy+uFT24caZ1NNr4/jgjBIlyNu0GNwYQdZr45//3AHawp6wyjbjOqtArZPBq
6dgkxuaJrs4zhpANDgDFXdwcD8g+v9Mz7Ih0mBxUfWMzkNendsn2Iw3dv0U6OKlb
u+FsirnqnXMHOWdhaOwFV4fbLd16CyBBYnveezNBkZ8PX/JnBPmPk8/IUrx6Za4S
HzhA8yE5Mh3VifDrh625u0T1qXWI8Go2GUGe+qvP8tk5wA+iOULAbIjS2fBzG7T5
PI8b/yoM4xNTFeaEVuE8BUKHHJF4G3rkmT0H2OPKR2B5Y7f6h7VLAikg43lDZLQS
0dG5yLPzXyFsERVdWyDZC/V0anM/Z+XBhOE9weXz0cxk2liqhTdvfwYREUPMqcqp
ppA+Ye7bmjIajqGjOL77u2Bc29Ry6sJBOhk6XnN+AwnXClaEqWFpvHvqGfJ4DkhY
t6WvwYAwJ+EqnCtyxHGjbWEUzi5IlRawQBtPbh75jt/XiRdQkJ+GpKsnh82N217u
r/J6Hx4DmcEz8OLADLNEshVamrKIJVWhwVH06kxrZiSC32mVSd4slTURvQP44szc
WeLAnT8mseqdLb4ba540J63zTiHKpVPshCVwNtXo/dX1XH0Pn0M+KOjaMt2mgf/i
Ak0xsI92eoIcNn7l1mz65tS1z7wVDvxkEpkfUjTRtK+D1Og26W2Vf2aa0yNHBbbM
XoYuuOoT0bWvtcyLZ3kmCnaNF5n1ipWsPfZ7K5t8/GrdM1tX4ZvDt5dIaVpjgpBe
5Bm+s+wPJR6/cFSAi4wxlQxUGzmDdrPHdzS+P/u4iVLYCaPLT4e4m6ukfx41p3ZK
uGWzg8rf8V3CUCpr2hBfFi4CElyWm+ACOVf4GYtswHO98JC5dVjoBMeWB6C3tzIQ
PcROr36NfU0EpMpMeNr/0rC/ymFdlIiOAilPKNMB9BF3fDyASKpof0gvWrVuoulZ
E0bKGkYmBaG+mutVGNpKbM7pWjdEgGyBXD5uNS3lC4T0JockoQQAEFdU/4wOyKKY
L1RkYubH/WUwj7WMt8n7jhaMFf40UaigOpj+0lpYxzt0mzNpqqSEFvyu/FDySWgA
8oJYJavsxO3sBp/0WQ+3F3Y1YxXzJjUPfDSfY8Qwaixa8Dbpty+sALaz9yjVjYn9
Gk5KPFvdgY337mNKdNYUmvaRt3nIEDbYYv+zIrx4QoH/i/KYuHz3ctn6XHqOY9Gh
4AVkUonta1S/XsGdu1mACk8gKz4XlVvZ56AwNvGYqdxedAe1w9ccWDeGRk9m6Rf5
Ny8P+Tk08dwISJz/rZkvhxTlJjr3H6al8NY+3b06gV6tgGc5zbtUU5iCpi8ILNJ3
Oy47CMr5HMH5GRRoLWxxs7Lc7TxdISr1zqxblyJoK1zr4D97m7Zk5Paag959OAPG
GGug6D3hVPTHUtEPjU7z8hQ7cNNb/2o6fX5GesZo2dlybgx8RJ42BxoyRE3WB/Ah
LO1w3Oh9pnDoxF3CI7yGNsa3WJYW0wdSOMk7dndu8zvN+MYszpmxcyXm0eT7ZEMn
Hx/5PK6B4Z9PPM4qN7QSZ8MF75c/RNzqy2qCEjkNourjpQDeDEp8/xYOjAG0jdkb
jAahcYEBdBeG/bYcByAkGiZWYCCmJ6psFthekCe5LHmT7QN24QL5ECpV4DO95mbx
eiy7WImRduuySo6jh0Sjsadxvq4GdDu9LP8P+9vkr3PLe5fkNxXw7S27Yau64F74
XAJ1uKnMfmvoLvWFnOt9k2+C4AfpBfDYJsKRfk9BGdNg6LZ5Ejtw1kqv6JcNd5ZR
0fMJ/QHllBqNjUrsyymo8Sj4BSliNhU2XSLAMAMESJqIWiCKwtJwEcmW9kDptUa9
RiLMEqyYIX1wIKhVNDX7okgZl+ytQBWUcYtxTiOjUnaiYJGN456JH66I7nG5fnLT
6+fr5JO2VoJ9hAEJu68NzdlQhpBpaVBdjqkJAaO7vJTm5ej8+f++IwCbUr7zF+i+
rlqmgJB5p5rbZwk2QGegKOuOP1Nhm67191vLpHgBv5axvEPYoQGLMVP4uzQD91Xe
G+4wO0tFN+nmoXql/kxCVAbyX5ruvhvZx4BCmnaMSc4FfXATpidtlB5qRJP6gUAE
8B0TX/ATqFfKQMC1AuaBfoZaRvmVETpqMBaUMcgPOuWG8ocXW0JFVqkkDXy9kGEm
6atSEfheGvyc1Ywo7+MZic6T7nPIHyety2/4Lk97CcpjghvE8Yj4xvvhTFKcv+j3
ilqCU/eUa6JEsPBtGfGT3nOI8m5WorFAiSRJdyr+Sfs1J7ZytT+g1tnUs35Rc534
T2wvfCutEosWnm9EOvAnQyjwyk6SGWZNrIIu60BAoSVByWh+MFYxMau56yPD4whN
jE7DDLJ67CPiGWEPax2K7rw5iL0Dss5d2k/UxuhdG+QlhH+zCE36uIbVKtnLnxhC
dMXIXdK4ee5gLSh+hN5knSR/Hp6D0ZHJO54ZyWPPDB7DFJMIV+ntbhlka4kxedfU
CuzDtODVFDSOBVg1ZgCrXFl0tD+UmL9fYBNBjwc4r8HUjdPzTG/yzB3FoZ8hEyO1
G02+csvEfas3/v445/wyJc2SQ2nT2ex8Q7Cjbiwg7qf/lB+4bNTtM206hoBh/38s
haMY5+AMtSAqN6fGN/HUn/E2d6UxG0a0Qj+S9fUsgQf4QJL2kEC+cuddhmfIee7W
CXa3BQn7rLIIWVSmmuXwtRefd0saF/b0l1MOERVQCbQDLahChHqU2RzVG9n/b1tM
ykrEN/SlzXHJlGCsHPY13zN1YFwkeAPx6Zmef0X3IFBLu9vON5FibzRRQDgyuyYb
SlVNgrrX24EW3hPgKJEJbAZFTT371TMSbEb1li3YXZRzw7ah1zhYmlP34qxc1Rcb
Iz35wlap9qTljYyoYwIooFUXugUx1E1M/9RTmwowm3PPUR3fYE3m9bpWuT8zsJJU
h+e74szkrl56MgD/7VW+a185LT29N8D7E5cxLYb9ebd4TxIxy7RXjlFdbCYj3g1/
RBs4yLXAon6nxhTl6nSSgG1I5Hy7y/hy2S4TYAwzMWIrNCMsIQge6tHb1J5FUnJc
ZhHGKQI1fJXkFm5UZLNH4l43SL+2VDvxz1L3F5XOKc7fNdPuK/GqQoUlJCQ/Bk0N
mrFNFir+zlQIRVyctD/OQnXZoiTCOYjJDEfEmPTVihDEy2QSx+ZMudYy2wsH4Feb
ADua+gpqVL3F3O7rhvw9mbnMyNDmUMWUZmWgC0MLqPyJbIPpZAj0447l+37o6x4M
iXDrZ/vRvGbzDXxv/OWCwl/PnlZ5xpxwRXr+Eer+V2asJdQDLbBcApzhISVRgyDQ
U39PmyNOZUqm1/5rCbclrHB0WBrzDgmhacnxmG4VC01I5FNrkRwGXr0adSo9/cI/
HQILAV3BqRR+LYbekgFcK1YN5V9SZwN7jIWUISZ/EpQkzpQWnqWtIblZ8pPAtQls
LoAza1Q14n+1vQ51dvH0fVENBUeeLR9VzDqOkYBdu+/uRHzL9VpInCNHcMUfpmYv
sUuWD8FwV9iqrFabSglhQLe+tmaDtsWjX9VSNxKJ88OgQuZXsESeN7YvfcK7Rt27
El6BS+39Oj/gDQwK1zleeHUb94nB1H0X1yaereyqdkhAObotT3F6TXwJZuekm06z
5E39bQCC0iBxpRd4uF4C5evsxHedkuWfIsdZSmd8u6IZO0J93RDAcCZSO5rOpRlw
R5vsVURC+MtOXdWovPSrInIb8jgSQ/EmcYzvnxjl2VMtFvUsadytd6f1VEgP8mR+
KvifLb/zl07cdCyaiT64K8AJQnXRlbCHdzqHN53pCy3fumEPFbiFaz9FuxAd3Lo0
uwzU0xcG86G8QSArss13ZkqxFJk3Yo+b+ugmps5/Vl/90Fu6TQSEnsgzofOqmAoN
l4HTvUiIjcMLR2NVt726Nqh+ZGsIHSSirMuHRRyoYCYjXJWLtazvD4J2uPJ87RBp
PLo51i+YjwTzh7icJclA88aYt6nUl91pDprfaTqHGNX+ndAfg3WmgwoVI4bnyGDe
ch0++ximR+GE5lOigc+LCx2/n0L4kr6DGjSjfStCTEPvUlcgv8hh0Wqk9ZwZh7G7
fMO7lNXkbnIufwiEkYkyp7RJW5tdcIJGilE8FbW0FxlbQd8xhaO6YVO+3K9xNcjM
SuMpyUfDnPDA7RpIi9836Td5WdDjabkqG3sgqP9L5kWUf1+tGLqwmn4JaAAUn+44
TaW3yfWJvRSepZbfO4WI5MeQIfHLajiApJxeZIFjqTDkIPoHNMYPc5HIf2DMclL0
yEsC6sNqsS3gEeFD/pas7F0hF8UOWErH74g7z+XkFLGI+YRm0xkkVkNvxv8CYPcn
4NyadsagFclTJJQAUKz6nBytNa3hgjqpt+ckXgik9VRLaoYyByVKDda/NoYmW55F
DFUf4zhs6CP3XE4cFtugOKA4CZ1ZfMVywa/9WRWQ1zP928nl9eoG+hwecB1rGyEW
7fSpzQ2I39tAotMEtWfGdChiXvSzZpsm3Wyrhq5Sl0YpDHViELrZ+JV960D07tdt
hJKTV8gBtijeZXpMRc/5OIpIIm0U5ArD/jEbtcF8GxUSeRezxuLo+ZaUKl7dzMw5
QKVWwdtJit3IOgki/reIiNXpQK4hEgufyYLvzeso3Ed2AUNy6KGRMwRLt42bRQxz
`protect END_PROTECTED
