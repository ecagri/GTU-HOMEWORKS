`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
joA5EdnwYqJMQevY1jjdymHoXAWUSPbHR7d9VtDDTf8jLZxRBdko8gSFkHr6oj9P
B6Kn8/+OTviKbO42peWfskf6v5OYczOOck7y3Dpd5Zq/e62b6NZiqzHp3NCNKGGh
vp3T4U5805DoSb8ddlkB0aZLkCbhHlo8GQ/PZezG8z6NUTpSImld3XvA5rl5qVsQ
UT2Gj6w3SaVd8w10Dfi7fVi+rVjMzkHi+EXYNgHGY5+xqdSCASGBGD9vMqKfOXaR
I7EVnLoOYBjp0LcFJN8s/Kf4c1V7fVyLFbad/eoRar5EDu/x3upkC9q/KQY/uyur
n1BpZLlGISQ/55Me8gXILUcwEQSO+mGY4K1nYGy+qCVB5R32SiDYiIqnpNYn0JmK
lTZ524fzswU3CPNwatuuraPK8axdSGtJN8L+9/fIxlXCUt+B19kW0zLpqYYIb76E
gLmpC6j0KugW8v3RZDRs/cg8gdXH6i24uY8OkkP/yTJyEvmKP1jwftGmXBmSq4As
Fv+gaBcu23qgQ/UZDzMIW83L1Zlu8Sp7j18DINctU090NzrA0WrHEyqeBmpXijUy
SEprgBQuixfZ/pzUXmrPWB7XquArXY0GKDEvxb53jBtAulYC0wwnMl41bATHeCvu
++CFDsg3oXR+Q61jo0l1QePyEQ/zQ/T3SCqplCfclzacBQ64p3U5WOPRM2CFO1ib
FV3HldZjwQ2wFcEyEI1arZF0CLRTLmhBdLBDjPzPHyaFaU+W3oyI5IQsXVID+FrD
eiuAOBvzlRZECUbDfLEw/S45SgrCzLE3quWwQuuMbk2GPnfy/CPiiQ/aknd7t5G8
7x1qbnxKLwQT5BC6tFg2Yu7D65mH1pamrcYZbktreeYIdlmvYjkzfmsxge8vAlCQ
MK+3jsalUYe40hMDZI/iXTAqVAK+/Knwv9PUZ3lFOyr+faItI4KSbHvj/JpDtSjS
v/LJMtVgnYe1oa3Plw1aEqkhVl+LMjZ38hz1QhOFUog4nJs7d/GDo7o13FQBfPyi
brGhWt/M6umdTFGh0fUddigy+QOCUNS7VgHBOImrPG63Yt38bNpcfoSPd2SI+KOE
9eCnhhHL9Jrhl0VMD4p5hz90aLucllMo//Eyy/sZ2z9phGYvBSdB6KIbOOkVQWER
Ami6fQbeN22nOGgyma8AjRiAEVaxN1tjypSwna8aEMrhHmXl2NzSnDPmElh9Y+BZ
eNY3KLqUgbKoT/Wyh+c9Wxf60ZCK0vaSwIoRoSD0LRGc+k/f6SP2dn7mBQ3l1vhv
4XXKlUwCG3t1mK10d34TBN6HIj/OWff1faZDOLo/UdOnmCPci3VJuw7tkX8gmGXK
K6F5RB81DZh8uDBBVarRBj/rGJy/fH7/uFDeKh50Xu8mGQcOhkoik68+KtNQxzwI
F6mtLjtxX1PV6FAF6Z76K/qc6GKIBN9SCls/EJCyc1Ld/Mv+upynNpqPWP3CA7GY
YlWOJKMlN7z/Zky5X54bbE3/EDVCNF75W1zkLME3Vmcz7IdL8nvmlpvO0ZPb9STQ
1GGuYaTjzc0xZ7tXQRuti+yfxb8wN4wjJRJAmyOOtTkmzT4oQevMnT63h1XGfOaf
OIiMSKFaSLYwrX4t8yKvt0QR1hXosurItdxWv5G5fo9HbZ8HZpN4rppDTUGOAgAr
frg4gM7gHY4HPfHg5nCrHKZhVyZ1cmZrEI8ScMPVmMecc6eNAcIk8uZ25RGFszcS
ZO0NVoYqeTrB9WOSMk8ps42FSa3JDcUuYzULKFzFoVZ5EXOJ9jc5NARrtevw9Rga
XsqyTJ05s/xNkOACWyYXKaI0GvnCPOhk1oqDjhUX6RdqRR78QLez1xCDbz+9Rq7O
jBVwpiLGT280k6WkNgDsAFXw1w+TQP5tZ77h5ur9U/wItR2QE7cfoJKi1PV/XytM
qoOOyZweho8xl9k6DvTEpXrNfbjtxReixl2Sh3miM60DlDstaoZvygbvXEpMlQGd
lGjbqi7D+4r1sz6G5tStATSY7Iw+RisOhc0eB6MXoEjytHENcvmDyhGX9Ojn2yz1
epFxrO8HZ+C+Sht3Pgm6YOXisb/GMUgPQe6mdml6HsQYfSlaDOTdU/Rq30fdQdoN
VuYvTzywyiVxksSnuvyw4ShVU0l5WhTT34riZEptG73U1TyuLwiEVVQODik48E6i
YTMIikRLfZIPUAvv8ju95x+WfpP7D+0TT23DD4tQzo8DQ9gBnD9JtXR38NPBqLrH
ErQ0UETmiAEjOQACgep15qz2S2YzoQ6ZJyJEHRwJGIfhAe7ascTTW1eN4SeSi9wx
rCg29ENeusqxFJpzK9EW6jNk710tFYYk0l3E6BJ4ZkA6ePQHWC7WSvMXFU667lV/
5t73IqYupUPxQFwbVEWdhvJ9dB81Uu9HduSPCIKiSskBLQXfnpG3PrbMg1JfoqBA
XFW5ia9Tgb23bRHaoQKpj8pP+IGcjIcsFfHEdxUGlB8hAtzIa8fb47si85L7PW2u
YAcN9dIthsmbmAds7FzGyQsoN7oWNxFjrv3CA6KxCfnc+OhFLx0zxANV98r5fKBs
wvLysrtIjuKTXYz1eDQhCvjWj+l4pMf9upk8/7iqIXno2PSQIeqbln6MCGrqYOSU
s+Qc4lqyl/aGqZ0O9ZyDp/qyeGyZRLEZ2H0/VtVHw3FrAge2QduGBa4yP1sIhqiG
S5k6lyhtfUTkuBxp6bOrmxJoBm+FJT+kTCI2yJM1BRQQPIgsFmK2VWtAPZhs6hbc
SJD7SkrTzYwALOtif/cqox144rohmkPOVoqe854YUyz0anHOlkVdlxpj+R2nJllx
T/B6fHFAmT+urLjO5h5Pw5eqPSRQHhKmo9c8saVqKzDA0oBeeEsXu2criEHoS4HT
miE8bM4LLUbCuVVFhmsz1OfvknSxMSeBcp950UiLMTGtUTdPbJnMXEn+x7nLZSBa
R0wNRo7ukpyo9x/E1bgdLtOEHDRUxsNYk91DZ35mHIvphh0rT/O87srFSul29kML
Fh7TcB+mmMxeRUcvtdd8XyME/In3GbsehTox6B4dtVrCQZQbnJtUc3PutmOvAz8l
tswtnvTFM9MlpQXtq3kcl3YqMd2z36LTMSyOQKQ69S7r0EQ4xvo4d/NzpdaVUiQO
UjE+mKy8xcJvmrOLrXPqf9y4dQfX4mjKhE0YvE4Fb/sIpYN1kIeL+3xXcr4RJT1E
4MVY1j50lP0L3qK4YB/6rWT17YkQ1jLMUxdbVWgjleqbbBrvGSgKt7debADpq8nR
dpNJPu5XnhiOpXrvMOlPLNWW1tyQRwrKwV4Kb3X5fwVnjG3d3rlp7TSQbManzwYl
OcdLlG5zDtL1JZqCLpKcbXX2x1Lb3P2l302+gl0Jxh57mTJI7eeSEYsFcGhDqF9p
wWns2wz1fU972/5TQB34wQkmHPyrxZBRuB7b/32/stHA2VtNtM8mhY7BgvcRLuJw
sCxFMYK2T6Dug/+L9A6oB0zTUm3bc2/dAjB6UNJN3awetg2IRDYD1Nt5G6HgjM+8
OHo83iKnyUa1LDYVG8UvdREZV/5BXhKoZcmtA0fe560ToWvQLXF+oBXYJlnuIkDl
JK6cYidImBN7cyFi3aBtYHqQF8o78YBLDrgMy4y1G48qQX6GIe9wVnAC+q1env+f
3cs222OUpIyalw897LkGO15GVRjOnm/yblRyGXgLaCwVqtgPlZwcXUdVdhlPdx54
d4m0+fQrGmB1FzVl9C9dCxGK9ncgGrO+6FZv8iIEUyatwAa5MIIQbiX7Zhu6WYov
1iq+j7G6iitWzSQOnXZmR7jhsDVYqg6NFW2odI5biJJIR8UcwSShm+I3ocPxrRI4
x8QF7vKeseQY16l0dkENjS96hsZqQ3sa6eh7kLtSEvA1Pb422nC+H4wzOu05fYuC
gYuEeYu3nEZ6ZaRhZqdLVRiMxt466RCZiPlGZdMP8ddKLsHG4d8POcgvRb9ZTi6I
1lqfPyKnWfz0TBxF7AcL+XdTxUxaKiUrIDeYmsvi6kX3AFij8MoFFt9OjI43kZDk
kMBfOHi7pSwmZ4vSUtIPvMYBnDJCmHeqkdlC3jhaA92KDOuZ31u5CWaX7bSEWpmf
JQM5+4XfKXoF9U15WIbxaR5Adm59Bdj40xuxsiYZmAgbU8LCrGw4MfbNqvo/ycUt
A5hvL2t3ylx8ZS5J7+0SOLVpZrYeUFd0NxEUKswpI7+dgSC60eeIeq0i0Rfalc5H
KYTvIbytjAMgLCXPogV06Fd78O41GuZ9zVhQOZL5hvYFf2WSyjiz1/5H6pVTKasZ
caMGl/1Mj1qVw+PkW8shBuOxUrVPzxUdPNcbFfRUWQhuCvi5R9FaSXQz1a4SASdW
R/VHZPyqTXAAnuc/HbLtBAaNDmE3h3SUtNIlFpzMvTtKItF8oZoSz3AwITad0++i
nvcoAzyhU3E5MNZmPUaKyiGP9WhCjXWmyYH7Zj6nZd9zfK6dNG6SRL8V3epNnab8
rOdvQ7sg2nZB3Z2E7gfpwmTOmeYiZGDIkVy3VdFmcjMTzwTjEM49L6D5JabPF8ED
ZZ9sHzXdbVLoZQyKPOsw4SzrELfV91dW7eVzykjArdzp8nU/siuQHM2bsPf24tAs
ithAbzu3vkSldjEADr8UOcLpN0AfVMk6ZrzugEW2XyGpNprevJSmGTpDFhgdS9Vs
wSy56bec6ptkOkWsWiK6B9vWreKbH/3epDiNVyer+WKqY3V6QzHi1U0l+ptGf1rR
qO+mZdDswvXZ1waCeqFccbLAECXsCc//wVO8YzHf1wEhZZ0IORLWLe6xNPju+9vv
h8BRdlSCdhdV+LrpAyiYoaVt4XVOKlwOxLia7LBuTBHJlWKg6xk/BZYDLwgUvflO
Rg3LNFd0K3USkt3vC1rPP+p/dbXWPOXy0TAR2UMN6JtvxybiTDZGKQG+wyOPcS8x
6d2Kgzk+mf3VkUBj5+646I0gegT8nKeYJw/0UKriZmOi8WZ8wqSgCu+HtXesHiMr
KGXC9yZrhJOC2b9W0e14qWcRfkDyPmHb4GMTnUaIPYU87zTSvBHD0aXTqvsEHCRK
dzwX0Hei+FCmQ8Mun1q+5e2qzw2XwW1ZgaKWW8lKoq2Dn2GWbribo424Lq1T5R+U
sTGh+sYISANlsFxdnTQK14WAbI/Ck4CS57JdZyDQE7h1lDU9IDt76HA7Y8iBZ4pN
KW7sUZ3GV+lN9QnGQKrGqc78H0GKThM2mICBSwe7Dy5mVIuAL0BDwazFeXkw6/2H
H+zdVOmwCsVF36WPRx5FuQogZn4U4EshBHX+qIaKIJ3S42yqK+CGykYo6AsZ2wbR
iGL7eVxBMya5JGfMoFS1nW8Fi/54vqrseXFZWdvST286LoiDbeIxxEt0Kojgm2i9
EaCktB1ApO1zEKgXdzIw4HIlIjdcNZcpIHPX16NYYijJld8a8H/u68iCIW1NVl4P
y5dYKC8Og1szzPvY+X1Yr2SN1sZ18Auae54NZxoVQMtLpgF38NaMwkdYnHbf6+vx
GPUmqKkgP3Gln338ieDbNhH6zh/qcV2h2XqTS8pAwPhDZ4o1B24SB1cZ9Iq9Z6VF
gWIklbECbmWAH4KZgJGWFexqEXOd/IACfJzftrdVZiM3e5BdAOIqPZgsdDB5elH/
ctn/DIY3zB+GoEl8YVSlBYdOLMy0Qbd7A4yQx49Bt6x9Rtv0YXvnI/XSlxMUBzoH
ckL/Mr0LF72gIJK1BL/1Hpq4W+uKN1bh5ujk1US630svPcaKQSpIX2Jm150YuyBL
ll5OOHeoJ8DLurrtUxAt/tWyrU3z4eisOIWBBKr4OtbsMsv2I1QWB0JSRltq9WMR
GlDAgesgLkP4Q1KuwST/SxSw9M3IeKC8fRmMgqGP7Eb7rpbE+l4A50IWBZbQLAXw
`protect END_PROTECTED
