`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8F91aBEoBo0cmYKhE2O6Ub0+4C/k02oyisrP4EaOnMJQgbp57+5IgrS/adkcSQdT
xuO7VlNfys81RT5Sx/LAIxAC/XACjKQ+jfyvnURwn/YKe5m3kfSQ6ERuDiEfKGM5
5z7En5oq5bIGAqnH96cJ4z/OmlzslEf2rsfY3IbvFM++D7R8bXQXgaVamz2VkWN7
1MZtjqNaSDoNi/x3+iinIXgpeP8jGcQdSOmaws7ge8d4OearyKBfd++4cQUIWYj9
Ok5EpPOS7mtsPVVtKccwn4ehm9Ww0JjiGnLSkTb0IOQnzO3hoUVh6yzj0Oyi0xWD
O1j3ajcjzf94B1kILbtOjWvNON3KY/cUIxotRzA2L4dotzMA31VO2vcxaxh3PgRx
7FkOQnu8Jy2UXKomtZNepFvEahFjMzLe/3/F/hciPaqfmJ19niOvocsLk9OxdgId
41aalrXVKhnIW6NLshcVn9iuwO9WXQ0iuTIAOeu7I0Si+BHp+04z2+QiiD6Qwk0j
cYK/7bovU2OK6DB6kIbj/vGZpZwtZiLa0MdurpiCwYKX8n0ZfGM2afUnr0oI4alK
LkBxaGsEyqNkVx/mDTyBAnSPNRTLKI5/wKfi7oUWvaHX+LyPIVSA9JuJfoY5qFaF
l4URlU69SMynBocGC8z0ysCPRpEc61+55E/EsMxSbo4f9QSkmpcolgulU+EVI/DN
jSrcz0OeWF7dx5Vzqfsg1QCVJ2J5AOf1Rd5xL6kYBhdB878wze86aY+2ldUT/G7z
AASoBx7izSLyS8c4GCCXfCqLc3QaUL8rFys9ofcl4Gpa1dvLdxNVig5Rx9ckAIUe
I1P1HOsn2SsZM7kDbLGI+p9szFYqkahKEBzYuA1lGBHmLspkYowk0RXua0wXol93
087sk6SdaiFTpgfRc5eIuY7Mj2wYdcwcthn6c86In+cF/hkA+En3zdUwPxkXZyYt
va0WeKUtTLgirptxXIiLyVLe2HYdaART5Sy3Ju4JRx7XHv/mmbcEqqxVVFMz18BJ
NKkgyE3diP5VOtNgWQf1nW5HucKziQDRhU8XFWyqCgIlX9bRHlQR4KS7XkWe4Ld+
P+DMj1Dhe/CXYegmIp9rWptXMhFEolCxzEFfkPuerptYcbkl01bQT17zTiOStJaz
esUBmLc95RFCusWOGlz0sUIsNzS8SFluOuI1BrjemQxL/xPlYuyua4HbDQcpfMhK
43Low4iDSV6QRInoxbf3NBw0Eyjrh+lIytyH9cz5D2hzAhvzvC6VeCjxHOmv4FLM
V8wd5zSlEZbDf3rsO1JcpQmUFYk+uHFlMI+8WboH6BnOJ3jANM3q9VYuqdI+DKTf
AuD2H/4EEQLZQxdsQ8yJc33+oD2XFPx2rJFk715V1KDl9qJzt+fQhuyW/iYaoYmV
nibixO/x8VZA2kseYJE3lP+qKpGSik0v9mJgPN4BXNWvywujt4OAGpsj2eonch8t
NKKfmdXkYosVHLU1gH4JZStqIBL+v/zvz4MPfhZKX6op5EzHapWB2gEf36Xpk4l+
Yis8unMetYz1eue8LA0ZHd3q9I1mpQ4h79gO1QvaOELVgn82GFUZH+IDlnVu35TM
N+gc46SeMC7mFSiAWUKmTE8ecj+tNO2jE07YNDB/1OD3F7MF3tewKd3Xq9JhkBwB
Rhh7C8I3CVXoR2az4gjjwsG+lWx2gqrL3EOZyvvrUlMH2z1pVNcU0nDNAT089Dfg
dOObrGgzWiNmR8a0gY1whbhbEagfKrw4Z1RuV8vhq0ZSPBYWEJoAFHszcmdO7ahQ
hTbVSVefrCFjgqbIDe3qdY0emiwVXB0Dr5s8mttewE/jqrcnTRsM5Xw5tXqaFlTG
CyErMxyMPcfVg0CY3/rnDuPQpeMRj7SIYcAWGuTBYN/cQSURS5CmQa775C6meR6a
iTWBo7Fe8T69IPcqh5dGir2rBYop7F4HicuLez1jeuaXS2UZXpU0h/gZ/pXlMIQi
OXzwKGR2pq5MkWx5UIwlvXwwl70XeLcXcmJgF/ug8dcXmNrA5t5UoTK52evVZnUB
ev9YL+Qx+Gj6l/6W7ZioUzV1T8yUheAvmnvD/OwHmZSFqhEU5lIlt/6TA/oNjkVn
V2Eo0k3uAJ/6DwHP5Jka0vDMzSI+RAwAY/gq7blPYAVq3PP3Kqj4lU9Lhvur9wD9
BjOHqIhyb1i5OyMz6f6SaYe1aTT+x6UB5TERyV4YuHwFfjFfz411rY0zuzv0lCSB
fGhg7mxRVvvC6DjwLvTJG9yygCslo44/G7u6hvF99mNvBfB+TDkicUNkIr23k+iH
PcPDcVGpMx6lPVRcnTLdN23vi+k15LDEk33ZGJ2eJLkf/CHemtYV/Skude6vZrKB
3Xz7lC+SqbS9YIg/LB2Z1sm+QOP81HxHoOJOICt/Ue4JirNY/nuXetsXhsoJOD2k
vSmb8TqfyokejsEK9xXLYfNUz8cr+/rsz950ziWi7zaBsipZWvyIJpFZtoIe6soZ
+VQZeowOBJaTLNVzS/VXR36ceJaDaFBiHX17fU9oCmpt0lFEy7VLLv/SU6jmtWSP
0RoSumf9tE5GghZ9JZ4f99CHR+jXr+SWScsGbv+y96hDDP/8L2f6DNmWc3EG3yge
csQNAYSHNAzhW+bzKAvIGl+QPSWo/Q89NuOC/x03WW9NO4UTDM1is0R1NWPzex6M
Hfs/TiUMKG7Y94xohnt1mGsnSAVt86M2JXpA01dy4IS9qkkjuwIRCs96nLePkJVe
5nIAqD9t5ETGXRXHFD5hev9KbuN+VxWQO0BM8gpYP7vG+fHhlUhCRKf46GtIKpmJ
Wl2LAYa5teG3juwwlBPFVDso3P7Zicj2dJBaAxyl4wpeWuZd3PceI5If5gMIRSNJ
AEQiXT3ngJ7OzQZ/DqmvFemV1d/kS5NSR1RTgEfKnO0h0Kc1gQKfyh3Jvu/kYB4M
QUhoUM4XlYfsD0p/sVmwdH7B+zqsbZpCk69uYGCQhFPaHJDwZEKz3lVXPwhQnTtM
LXjCeGltsYf7ARCIPSsKyv6arHpCGtVRiY8Rjw5LzI7GB9nVQfciNF8BUlW4xLJQ
oCZuFLW9vUxZ9qXOnD0nqfzUAtqqA/Skmw8NrkQSeEvvemkTt9wJx+LsXDKCkDh2
y3X/oWhTSLdAZTakzpxnTYRgTL9aTGy5vfouRAzyfTF5yo1lSWUKFkAxNd6QwOng
vN1i6aOhsOeGdP0LvMxSaFfh1ejHrbcUaqIcFnTNYhKRNEZqUWD5Nr3uR8GVBOvZ
Fr/dtKWae9uuLiaKURj6s5JcDugapGHYChsfUPzz2T/xnEb8azf61xWAl3TqFSWm
HEJgOa/1zMQmD3AFjS+oDo5yU6B87MXGDTL0X0YyrrqtIwfjxmkpOPrTdB1DVxsf
eTRD0qpmHJvoyMVpVJ2Jb3NQe+ZilRuAj9nM3iWrzK4SnkAbrGFmcxrpfxxgZfpo
Sh99rw2b2BxbGjWpWR0wus7BEDdJreZ5AvSK6tG/tfvVKLa2nGfNRoaHT6m7Jz9Q
kqGhuj1f0G3cBOR9EpdyZS0J5YD0VPjCaIkjyNuWprDnZD3u4Odp8nTLK1RRAKUq
LqjFgQXijPyeKi8G5ykM1ALG7TZiH+Gc+fRvM3rFfq+Nv+SssPlxpFlhOW/2cgRl
UcaM+6DtkwhKNzfCUlhmfAAFK9WBRT4ayqRlo/sQFS0nfa2cQ64uzgbKBL3hLyaJ
o6tVvG141+Gd4VmDUg3bNWVlJzy3Rhvka+ksrqNw1P9U+MYYIgYYLT3wT9XLliiO
TB4HTq++CiVxoK0tdwOvtlkEHn4crkrN1HGrwyel+LfhYOJzOQs9j+T5Ol8GW6yS
hNG76MC58AUN9n0illSTzOpEzNc+/UxgkVGJVghw4Z+k54v0y66I86/I4+b7L0K6
Zv/INFNzku2WJgC5T/AaPF2eJftfLKfCUZVCe3TDE/6ARt1VYkxTwF5GC0DcL6yp
N1FbmaHu0L6TnFW87fYDPaIblBDhGcaO72pBS8JITM7tNRQRg+aPAHsbJo7Iq92q
qS8OlS/TbHIOmcRdzsdkDM0nvLrvjezLSwxWibsz9cMYkXxrl+LtUmbYYqT6s9QM
adH6a/7FZv+WueNGXpZyrmAYvKwQrBrGY+VCXQuz6B1BJRDF9AOmq4IFN04e6UmU
uJKVThw3AXIjdKMvTehHhRVv8FcNuRc8JQ3/NYh9P++aAE/SWScEMN9Hlr5H6gAF
Oq6+Omsx4Wra14S+2+1Fy5XPzPuAZur3CGYSoSMVzGaXhpR4PrgePGGpSzcOsU8W
NIOR6elqxikMp9xQRCd7oqWqtE3OsXqERMxK++nSoXAN7lTSt9DKwFzpQXzCQGpv
Zr8FP3dke1jevzt/5D9RZwPmRp6DmAvxlRYGZOdYPVWgc6B5e/il2Df/2VUep6aQ
p8l/N4SXgTsTRIq0DC0zqfXFDKdayc77xXXZdv7HLqhTIwAGlT7jo1lbx+HaYIWZ
e0jaJXaMMa1d9YTdJSpHz/i1nDpktC/UwqxEryKa9ApTHkOtLe7wxVwnIWc4kmLR
ivQpMgRFKchcAk8cjg2JDCG0aKdYkxAIhzQr7nwnM9FztlfUqzyq3I/253/eyfaP
`protect END_PROTECTED
