`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pLa1k8FMaPU0KzBX1FCGGyYxR3kcOBdzUzNlHxCqL7SM8uUMNk9A7TK1zttaVQl6
7ej7fEK66FkQi+pmdEH07tkH/5CLz26yz9xPBGT9qfDsCbi1Df/7CcNRk+k5d05S
vFLpjvOjXVC5nNajzoHW82/CubwRF/XrjNdiHbF7HpbB29rlW3XIucKSyhW8OMAB
I5CycjXUAzZN/RQ8AzPE6o0uOR2Jy7x9EHy0qKYZY5yrnwgiZHYqIfDN6qsfDaFl
UMMm/hHmshBonkQtiVbDMJVawfdu5kxxSrULks05Hbr5pEmO4d8o+Aactv0vAjwG
+3rZHCS33lzbu7k99O6cGArWSnOPpgFxmmo22rXRNc3NGwCCmEHW6EHls2M1/zDo
qI7Ojp9NB2xrRQ038WYU2uK6/DHvXWa5JEavog3DLOVWqH+D8YvERI+0x66/yj7u
XkvMnPunzwYSbhHnD3rZS39SfaPQx9EkSXGdIKvebbs=
`protect END_PROTECTED
