`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
94XAMK/1p3vxoKQgnccKuoqfmD40RLczqd4fP5F0RMxu5GgN4lLIl8xQMcVaKXHO
UBeLcOvcWRxvvoO8kXihNVNPC58ssqFjHCkwTFBZvRgdi8nobpP69RfF6/3BdXY7
x2kUKjMVO9/Xgf4TFi7Z/yFlwXN57heH6c/7qWaGGeCrFlbfgFHTq/eclcDFG/1f
DBjefSx+EzcWfmdm1hMkO6oUIR1+CgGtzEXzeCs02J09BNw/dNROcew5bHOTjM6e
IyaWIO7sHQdDPlTn8ai3j2E7Lr3nZKMELkNQP7pvMhmwQua0KAqqslCqr07M4q93
ba+Nwz1G/rWO6BVRUMXh7kgFPNJKDBltGPeNRyfqsi/IPTfMkOK4KLNWpGDpD3uw
DqosqpS+66RQHSWB2MV8LItCybndqxqdrVVZUHGmtlwaGsCRAzhb07IU60RgESAW
wMUDoVr0/A9Jt1R46zs60+1BFvvYbZ3FTmEnHnKYFR7vmjpKN/OnymHElFw8W4m2
BXqd9x0QjqUY6t+U7esgTcW2YA33VnEu+XlKTeAAD3sYHZQSDWtRgmq0FfneWNke
dATSvxujZRqMOn3KoTvOtCP+vk4NcMJK3CMNXCrff0Se4AXL6RiiGms7DybXGGET
TxzRHCwvAsa7qb/172ct45nSMCZ02Mw1VU54+rczIygODrj5r88+iswmHQCZiSgI
AdJZJr12U3YnTD9uPesJb50Lsg2vAIP/HGoHh71NxlUkpszudLrO0m/VqVCrv/2b
43TiJrW77cMLsSiMVLH03fN9blR1BamNCZJJUHxFXlMSanerump/KuIL3RrPJhT0
FiXKtJzfJSU04dgrC3CzXyzQTWZG4MJlQaeBQQWy/7B9XZYi/mOyJt+85xoEJyPj
7PVEPLfY61rIxaPX1WkXzzJ2M39IHUS+/1BvMuz9WkeHFkL+GAJyzckX0Nn9wBxQ
Tv7nbIKHjWdwv80WyGu388JzKZisBnIsTKhX9p2eeF+RueJblBFvnTGZFzX1wzxn
EV622EQQssF/tHSWJ8GPbia9/FQ8bZuJ685CCpSxu06gsSL6M0wwK+3Oz9yRGbZO
JtWYT1CZETlf0qG6Pm8NUYcRWh5H5qG3Se5kZ47VEXPBcVVNRf7p3QMGpqr8dew2
8xZCWjNVKU+TUi++DCgpEVEsbrB6I0YVFukvqjayHQ/xPcQdlFOWYmWZm3L6wizS
Dt/jBd10acEIGSslhQwSkFZRwZpeLX1GD2w3WbYKVpMsS9wY8PJJzuc0lbCs2IEk
8lLgOAr6zqR6Shict0z2hyymrBTNgiLPLDpGquEamQZ9wD5JR5GhEvW7q/BjLyIk
zHr8QxENeZgiv/EA0+jRhbJry5MdjYT9wDaj7ZWQEXWHNO1MLILYak3FoOpvHKUL
arOmHDoKZfHutcOC0OQS7AKimt8auD7f5HkWWiJeCJKL/9fG1pR2GgJFdmhrCT9N
1S0w6H6IRS9Q1bkl0qvkWcyQCBuC8RdKl8atg3HYqs6cDaGI9tXp0fHQqHUI3DMQ
7R6dpvcTO85RhM4qq7NfTZXR/K8Um++6C59Up59RbvSWMlZqiaqvp5owhqgqB9J0
cNVWsUdqfyEqkZ3OTXtBuvA8jUKAmSoEZAKSngCYtWA=
`protect END_PROTECTED
