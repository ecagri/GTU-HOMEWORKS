`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AxAbfGTAz2T8542BQJfoYh1kGMpUta5ca8Dbl+3rtEOZe+9cY68Y4t3SpGFRp+EI
ZAoTn8jreEg38GmXX8O2biEemjUYAT9LF+ZnGxHPFn2KTRMo7KqAwpmI9dIA5zsA
4xetEoMk1vicB2YE1tbblXv4NpMPQRrPclTkquNad/PqSMc+h4Eg1BnmU5iy37L+
Tgn2Nv3hH33shtEoAsZ5FGjOGMO2cfJZv9Qd8CXGZnSv2GO/ky0YvhRqggkiKdVz
399p56Rnq+5lr4rmLopozc4fpxj0hDBddcisPnlCHJr53/lECo4vkwHqTlJldOH0
YTbY2XOtWTk2BmLtPZYlNSqmjqI5kMPq/12hPR34N4yiuAC6n2zNUEdfcBjPNAto
/V/exMvDMucOF3QRhf+sSIpmmYrmZ+O4Fdm1Sku/2UsVyEg2nptIQYhB1ava7o80
fAF4jZHS7QrDb8q+VC1jJ5XSFfqIwEOAFFL8v86+6BMSeKIRnGFZq50HfFAI5S+Y
F4rs72kNMn5GG3lzXsOrSeRiO+j4EcCbgP22HSOkahUe/g8vqYxEIVvIlgvhN/Ym
wAplKJcl0u0HdW7E2JUbejPEdJCnHSf4M9uW4N//F1ENl5nWRW/xnKfod2Yhraqw
4/fwjlhjz9inG7UK+ldsHNjz4j3sOnmy8JEaWTrBUxWjQPWmkGLFK02cYR0qaGez
aGBsYCTE9eOZDp1qZM05RdVx0FD7EVNqovTnqQjglLMNeHUPuGiOVXyenZXVuMcQ
qI3nAOHenWC/ZXBuBgqEyM3Ce1dx6zXsPCOjXVj9+GI9M2dQh7WO4sQPe6LkzFbF
ShmtGb6SEMLiQBaPXf1+DR6kw+ekLtwB4PZq3YzFn8logBdmtbr1XL6vn7IbpiuI
5h8M/3QVKl60VsDlq/r0k9zdC7O+EwLGDMJyvC6R3gZcwFXag3LhUdSez3q9TBmg
7iN+DvLZvfEFgqwL+3P5vvskjcN/fP8/S1rPeSNV+Bszr9c4jXDgqHG2t/52FN4m
8OP4RYwnmEstEOl4qoDlWgyH7q2hNAyPkD0+t0aZAUFyidebEwJBvcc6QsZgj1FG
MaX2gqT5zvT7v51WAEtdv6LOSstGiVPdpDCXCRPzElu9ssI9DMLBfhgN2qaAlS18
5eN5P0J3obt+TD1zasDIvmnlyAeVAGtf25NV1qo8A3iX/wL3+vN6YFPJMQpvdyGw
RB9VPz0fW9qUjhSdh8k/Ky8HJzbZL+u8rHdt9QvgxucjVs661f8xeEoWV5AoiIvk
Zwydb6Gwsg9dintGHbnnVY01D11r03DslyLimGeWRGvtPL4tqmnUN1IU6m1fz763
BqYjBWRA0AW9kXJiQJ1b57RmNCMHn1k3ocaXcruy5XJRLu0F1x8lKitJBksMRzAU
pTkt0jWHig8cjfYjXkkipzKCOAmbkmLTuJwpD/WtjQtNsWiGOZy9qei0hIe/8/HU
RiopdEk6pKv12nxYJbU2z+Ni/BtE/PHwE9ejKrPPWoIE/wfRWzhSAgbUofsT4Sr3
`protect END_PROTECTED
