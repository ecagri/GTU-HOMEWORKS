`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9OabzrpYgH4/VXPyaeReMQdWZoAMlGJ0ykssw27mLG/ePOrzbCZI7fd1efAgjYAW
YgReXSj6HNsm6SEFQabooYHKwTCn5aQ8wiYkidBJCBX5M3dHI4z4RaTIhZy9onop
01QEm9rPIodSCyFbv9uJKbPBclkRO1tbtFCNL5ECiFdBMeiJXdtMCSkP5cGDB6gk
s4tlYfoStggps8b8U/dHFUBaOJ2jZaTmW5oDznpvZZzB3R0Pybu8GvyqMMLiHD+1
pgoCeK2AA6IOKgl86tnogTDUO54HJ1bJg9F1LkjH3GtzJKILAG3cdZor64h41keB
RFSv/c7kKvU7sMRboYzqwae7t8FBYHuhlW2dM9B7h13WPs58GkEPMi+X6ALC+oJ4
1+ou06udYeJg0P5pPyJ97mC1EXY/4JAoEgvV4+l/iE0kEuDCX9oLbIgw9CMcfUB8
l2XETuz97fQu3h6LaYCwuustlL57XxDTuEdy5KjiXaL3eDATuIC8HC8/y1ouCb3q
XL+ZzMgM5QlDe8UYBbfoQ6DP2U9fGzqg/py1fBLQUqyb5h3tgtXTRIRfzQmx3vXN
2T/TjENR7CcV2rJe61/LvllvKVELYK7RBJ0gSFAOsjTEw9zVhuZDxfu7WD2Niagv
JrMjsOj0isT6BkRhqpE229G56EMq5/Gaa4JmwUbMfzTYyRoTJBweAR/Pw3/DxidY
LSsoMsLdBDMkHfsL0Nq0UBUjlrx+Q2TUxCRL3wOGcTakqf2VeC6GAHdqwSCRfkM/
Tenah3n+8xGXTqEvUFtaZjjoN33ztB3roFSYUO6kNOHbDmqLZUhDaWCSIoF6KO6G
nQ/EoMACFuUeQ3aub2wlLlMcsULgcgbFVq/MtlZma6+42PLaGpjpue57n0ULDz50
RZ+t9H/QilZzS7kKaewgon8E0HddQQ8Efb6NjlWlBNqFFU1Ei9NoYtEU7cz9B87r
1R8FajXjhtuTasVniiZdTyUcgBxo3ysEv4MLeoA+0sZnPjTXeHW5xZemlt3osb91
dh8HtdvhCA7tlTcQ0LPzDnQ+3GhAjX8o/O5up668IjCcaPyY3bpOPE8MA0xOUi6n
/EiSCfehFZZE4YrrphNTcb2SaCb9Dp1k4utA84ClM0zewYppjNrDGSb5stdk+mD6
jsbx7B/qx1h1+ib4WYhoXrMB0LgaAVbXPHTXwKMiNPwwTls7ijm3ec77N6bNY171
b11ZOrtCLw8RUl2kfzlW0v4PGB+Yj6iM+fSQAGzRBlaImi4nJZ2Rj4gyKePwJLcq
bdetHsmUmlcO6k+dUOW5vFXxteNcbzCngDsKTeemuXvUurKqrWE3HQ0CfoBY8UPX
EIehEe1NEYVkKntdSENhvoK4iqdqPtY30neKEtoy3np9F0rUuTiT/9lYbgNwgF03
yhGqyGTVZbqbc8n/gJFblQrhY/EOk1gDt+Y0WmChkVVRy2apl00OplJ+oWTR4hYh
gorlbzhZpyHLyOFP4p6O3VfrdFRKYzCfyL5VR6hk++K3cpa8rRpfFYMTNVgr6t6b
WQDBKzApbjSiLhJQici5Ze90sqdJss88FjY8ZwylCyLxEGifOek5LDFh+jB08ZfE
cGtN6+7XRp+UNFmcJZO14bqODm8MWiUfMN1tNbnLGUyKeupeqWkgKWxwz2spoS1Q
DX0ghfybTt72sOv5Zd5dVyGVI9NYp+BXKS7dHWYs5XvybnvodMv5J71ExC0vpRNw
Kpav6Y6w5v/Ujk2hAOKXamn2lALF8mUqct7rgPMkJ+yAEwJA9TaZQGu2bs6Ik7Aj
9GYlmNY1l3AXXUX9a8//pwlccPgkr7sGtZ7Ij78FeKeNF31vR9611Ie2BRMY7tve
3CseXoBe+/CHHfPIWnEXssQL/KoWgJxRObYWsriRzTZ26k9iHWnnyLVao746CnMy
fo1q+NGcehD79ry1kcCN6Nnv2gdaHRt03xVb1fmnxJyWSjc/z+Rkobyc1BroQeRx
Dt778m+pm2v4zl0YCc4kqBFNlSbygYXOyhM5ZBEtgfo27DDsXVj7V7wlQLVcRTHk
zLlHYuJNuudh8XlvhyYx6VRgbnXG3i+NjpVhJ4wq6ysqY8/7qaAjyc+oiGFEbje9
2mxSS3urV9nQCG8OfnERyGw5hx81hALchdqW7XoMMnC8VfIKEAxVNzvJqZoPIztr
NAmkH3N68OPNP6hZg6k1oGwJVO7AcWk01OJsm2VplGk81ADLMlqVrFTqaFFIP2nn
Ffd+FMaeCJbUhKMpUakbCJmTVPM8gezCgAPUEEee06RzWiNilvkaplA7bfFoL1bV
axO4TFXLgCFvkeBuZ2w8PvyxoDWFNlvWYXsK7S7s2L3VDUNnbhkeFRL1C4JECJtX
itHyyd8fqoAhMjx9xY34KsShFiY3PhKAmSaYQLghE5x1i8J9+LCciEY2Xlp0oUjm
Oe6shQ7APvNV82EA+Yla9Hp2E4bWzPuONAy/z/X6DFyhJS+AI9PxoocJeRB1eabN
r6r2WEgOMHSvUslE6/k1n8fvE0sGyXAb4jtbcAbw/nnTIaQXccvbN5qwANVZXDi6
tJQLWdSmpMYpKGfIGB4tPFr/T/+eXe1zKUts8NNzP3ELY5cIVr+siHPRbYa4mcf0
RiQVR5+62WYXjsmVL+GhgiVP6o99tcEVqu2g6uiEDkx+bVGDfkMVy30ReZVwwa2n
CEgRUEwWU7ukwrT8YfhgqbwtNEYS80xeRZgeHLe15Q8ECVaptP8oU0Jx4bS1LYgn
xGCWxnYaUEJegGdmMlIY0EL2hJyKXHIJ8sWS7SfrxMba6nveAA6xj+JhSQFnNNRb
JkQWe3lfLSz83kTrBelZdUUog3ETBdJaQvnLJFfsjtyp7YpAib0PNhnmKMlqIpcU
9Z90wL91NkOE7bEMTcbNPFE8c+Ai9h9pGjn2l2cC5G9ANb0l6PGfIF17Hh607yNi
Vtdy3S7D6ZwvR+ozrqiIYVZrjRCqauhRl3TpSXzhlsr6gk0RHY6WHHUTVuum2Flv
ZfHmSW50j2kkzgY6A4b2Fa3kuo65OBm9Q7U3GfckQJCE7d9zjt5Yp3cT/uxr3nyG
cTcn4LNBYEZnvG/9U325fRzTHyr8pPN975AqZKa9iY60/3vJdK3caZodYoQdl4lm
5uu1mG2xkEEsyr6HLWtiUbRlKt/o+ZzWsRn22FSFfhujPUVDgMv/xBdf/kTrQw3A
iXW3UxlXjLDoIM+dr2dVeghZCCZEJlcGSqjs76zKhdu/LaGNYfLiKlxdQhlOd2bj
IhmuxOA8jE3u7sFvmrVWl4bphMnTTec/d3mF9JU3wIsraPwfexph0oyZeKMes+lY
/DVjfjp7+371rCB/BXd1VYTYgbVnx+jDulihD6FUwZl5UMdVBuMXg68kkdSWnNDJ
z+aSaEM/rSPu+31tHi5WI2LasKyRePG3NvVNiBKGXZEbtm+rzkpSiUv2kFIRX5ZY
qOaBM08USrn1LzZPLi5Z0g==
`protect END_PROTECTED
