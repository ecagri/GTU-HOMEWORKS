`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j26GIFUm7Pp26K8A5GQYw+/pMtmkIJC0ktu3BP9LYB+yOOofbzq0sZcnEXxMkkCz
5UPf3iYR1qp2uP+cm3RNda6lV8Ew2ilEuO4yoxQ/MD0Jd4M5m7oxwmztvahLXLSW
v/jK7HqqwzpR9+4Qu+3MZZeb2Yql2joGkjEANTrWUV7nGH+OGC9Lak52wuaGowpF
HMYhzEw7nZ+rs2cUmD98AWIAMMrL2KhxeNUr8jr4L5vjTxa+M9Li4bO0eLTFx8P7
t8+7GVJMUq9HXdSt0F+rhIVb9IBiEqoLPajNQqvxWV84/KY5ORzbwZeKlcvflIDH
P7EiQbFoAZERdDeNTRvpohsn4tkLTfx+64VL3PbJGVwN3ovF+UbS1EU7IAzn6JkR
Khi2DjKXxMK6tgx+1Om8witPkJOT1BcfbEErOzLDBKJe9gYuWmRFUZVgAJYyqOfg
+nxXaAZKgP2QsgquxgzMmW9oGF8uYQwA7KHptDo2AKqug+HX1Nfew3kMHxdT6mBC
vRXBAgL26wLSVzxjNXXQYAOim/O8KiThtrX6pZlb58cNumg7sLEuvsiSMRjZbgD1
noUh4sTdoTrik+ROD58G5Afzm0MRZwB/Zh6TXmaVH++bxbOmUsVH81iWRHA4R1oF
X+weeOhZ5ryuYsEvf+Sq3+NkB3OMzavSoayc8Y/v449rJRY8R3jXn7SRW6cxtl8l
ltWjQDcfYaLfcjXNWqE+iixNCEtiQt5AkTJBEqd9gpL5uKEIJtXalIgWOYGqskyH
z03J/c6z2Md8iLVGGCxv95NfSENSmC20NaCKsY+5qDbQd8sG0++KmRbX1dqQb7Ug
CE4flikE9nXUBBcpGhCSt8Xmcesf8w7F1mvK25BIiYp4RZPbq4ocaBA9pH1A4ZN5
5dF4WtuTf8L+7Rqat4JLSya/AfArtrfY+Ki4zwhUOggZ95Z0TpnHgQZRg8kI6M0B
KX1UernYnoAxswKHb972Yr3K7vR7XdfR4uhAmiPSDZdmLLZHVVNvlJSjwcOU9JqS
IGV8qn3Tz4NCvRDWcZ/apBiA1TDM62hddsTYwxRFfYICN+uxvjYA3TKfxYzjtYuR
mKwEHqVRITYnJttrbRY4WC/9+IpHIWpkcafqShH2KhUm0DcQa8AhLka06GlnHmKc
ByLOXXOPKsW/CxDRVg+NlDZZ4xCg/2PyCY3nRC/qQaBcZuTYm3s6zkeCgZEUsSUo
KihHWcIrBWimIyNEZmIeRs3EuTy+ELCqCzqCnT7RTDaJjkUuRy95s2D6GWCCZRCg
Ai5MfEHnasrbMRfVht2z+okryqP5g7Bk1HvMEvjoJHXBvNrKhJNybonY3ggM/YnK
NG5NtbJxVB/t2I3xsKW+N/B9OLUNJ4A+64nh2Xw6CqwtpX+zrXDOTOOa3J46gEtC
n92s0EeRfQW9HBPs/loF0skVe2SKbAOFeK//BuUE8svL8xM3qN0+2gp0OqDQUPW5
v4tDmIapRn7r1Hle3TomY2Tb8yQoDObnMaurHIKCfdQ=
`protect END_PROTECTED
