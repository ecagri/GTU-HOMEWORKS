`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dqVd2f3cpw7I+QwJKuFm4wPUBca6Lj+EOCw/fd5iK+k5PvCSKl6To9uA+NfZJMf1
mYqVIJf/5A4QNDMlalPxKOKqoq0psJvIHzy50Gh7hANuK3IK4IPuqNYdtHz8UcX6
ua0RQSgTElxFkmBjonoge+QXqVVXI3SV4IMc63iMQkzAtTJqxUH+bVomw4NljsmN
5mpBeh0MzJjhCZAhhU2rKD6vGCzAaJom/kXmACev5ie1OvNUuFVDCKXsrCN0W6gk
XCJ9+4LOZWDUaN3vxyS1zpl3J6eJ3eYysoiPN318SUkAhqwHXnZry/rViOydn2/u
nw4EHVfV+oyxF0BeGbd+iREspzT1cy8DvHJ5HtVpAkUS3cKWWMPRrXH4BDW6JCvS
dVp/inw8pVLbQCIKU4kC9dHj5ygnqrkQ7fbJ/JmMgWw69l5ZAVjVlkOUKy31OPiN
bg33Nfs4SgfeMHVTMGwG6nj8EaVOpA0YOZs7d9Xkn4ktOQcUeS4mEYSyyNjoxfak
YIfQlVdB+mK/wwptgHTs169mkdJKPtuap4RYiRrY/eMGRg84eu2qPuiT0fTyxbjn
4UCupRLaUVcbe5L4Mh3OnPHyefPoofVeK/oGk0SiJRR9ufftGAeOSywVbyXNRVfn
RQiNvdyyFzXHOY6bGkypyPqAlvU7ulfdpZvkccgol7ZUpO3aHTmolJK76TTxhKpt
psU1aKq4HW0aRv1P8/7hog==
`protect END_PROTECTED
