`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DYH2e0DamNw65r7r0+SKgbMbN4gLuqZiT4U4/H1E16b8Wp2iqktTJ0VqiaOOFjIQ
EokIYu7ZRw6yqvKCpKQQKjf3kWDd0jlmfcUlq696I5WnZ2ivM8r06EiYY5/s/QDF
2q/C3Xjkw64FcJEy1wKk+0Z9kNnYO6gkdNKzm3QCQcfFfJdU/3WYjWpYiYNRRvgS
j2uD68yjMljC8K2JBzpVn4Rc1YKtjkD9tk3GYW4RQch0pWeT2Qak/QI6eH0NdzEi
rCqkOE8i2/tlMklPcqGMe8vvmpquzaFwEJ3MpaawV+MUMwFNsQVRsA7mkWMm8kbv
66m2/FxA+LikvMQArcURlCWMe/b7dkWQnUa8ItQCoRTrDqbf8/bWy6yAysMA0JbI
bQ4aWo/n4ZnwdLjshkHX+LxWKWpGR1HvlHbs04h2+EN1PLS3XpWEQf/MsPL/48sv
/wnYxLbcP0eSGaEfoLbb0dyh9/fiBqpG2TcRIp6PGOQMFwN+vWgE/0edCJBG0aqP
NvzhxoKP75FvF7mpmetM0+fkN9X4KldeTshe35UfRVaLlRjiZkkePb2cqNy9g2JQ
whBSKaQXS4nto+Cy7OP7ryE2N92Ee6ULsORCgprlAo5PVTCiCjGtb4p1ZRAaVxmP
5a6zcsP3JWSN/Vm7NV6GIlwway6RpdFnoU6F+9XM4LHJ0xC9xzUSDxkJvSz5qH9M
bTIegXVxoRCla0E8Yt1glDAW2j1m60xWAr3CK6yDYBFOjlxItV4H9u0TfnD5zT6W
SJ+2mmoa1O0NQmVl9oKXJx01+KJ+IwSL2NzqIyB2O7E/JekbtLieimwz/3Adm+gr
t2FQm4xpivyGp5y30f5qqV6rvJDtoAo297UyNH0jdZ14iNINlE82eIRNJLxBpg6F
Q7iWxJTgA8MoURqSHa+1HgtuFph/uHSd6CJhgC8IUvfXwp3LgQMRi2Rh3Wv0B9AS
EenSY6iAtQ8CI/nFHehKhluVD9bPjEXL3uZnSVkc4SxLUl/Dhkpk59+pCjEcJ5gg
58gjQYiD0EE70S0/MP9sZ+R69cV7pHUsrFoVA0554n2uA7ZD5I+KrzyvonEiYEo1
+Sv1sDIjWeF/dtEtoLQpDrwVJYi3ygtOiHlss8C78nv6nZdA6dEnM4FvYGDRK4rW
NaFf+eQkFQP+uicUt59G8jlxEOXNF91Nb3O4bw3qgjmRnVVEuXJRWq9i9b4nPNyA
RZWX/nD/n1tr9GYdXScpwVm/PtHYP/h+DqWetYrL7tG5RAVJZaMMNQyXt3cqU//K
Z8uWoZzMP26TLY5HD6JFnVP80yh7h6EZvpe9w/9U2fEzvQsUVOeEqqS67lbZ1lZT
WwSJMBONVaptdYSnn6oVnaRRARASHkqyCd6rtvxcirs=
`protect END_PROTECTED
