`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BFUEN1eKFEkFC0yh+jcS74wiZbnoyPvWDNt+vuYHC0WPdraLUNhrWLDiqNMAOxGm
oU7E6ZWVmXuviFoO+t/ruidrFrUdnV0i1wHU3hJn3CW061aUNRibna4qm+wYMG3H
UUtXo7eRbXtisHDLmCiIpUaAocBS9FteJbLq5CUXaqH6Di2ikYz5L0zIpVfno8MV
65RvhaLppp8MEAOs6hm+6jQzfZB0qL1gHGvprQ1XPOBUqkCz5XR1VKMcsI6g5WPp
JsVlUi/vRNYnQiEuJE0kHzr8R7aLw/SU6by9Ylip1YvBoaO9GQomTY6Hn2sACLef
xWxonppMvUhuY3x8ppsyeUPt3s0w8hKwsD0ej+Dpm8Zf8nXRyYNe9EYyOvS9IM+i
nRPPeHQ/ncL0HEfcfWMhpE1cuvt//iH3JuegkkfVreNd9TjGOrU8zMuduc1EJE8/
+Mi3iBGm0Vl6C4xQqML8jQ4+IbK7k1NxaEppEuxLwq33E4QMwqRdcltJsSHSBtxp
vKC0tzQ1ezCgDQJG/0aAS1F98oL9a1jtjynS0+4zGG68+CV89TImBzV5SI3DWNrT
IBPAkQdHPLATvHKd/XllVDoa1EjAZuM5/JHP4m/09kfq7Nt7Syh8xNfhIvRcdH+O
9vbw3PtWnfagAZN8An/YDUS9yVXPM91FlWACQgLwRzie745VcCX8TB7ft5uhT105
q/PsWBx4Pj1GhmQdDbDvxNgiKrwPMZxp1nC/HRjkJmdO7XCECeyu4b+mUFfRUTsl
NyO4Aw52YQJs8OvNOLHDZ9oesjW/iEkmQJgN7EvHx4G5FW4fXw0WuAFxXU+1Hjq4
xq7OPCNbpJ9BO5/9ZZwya2lIjIp24rS7MKTxuj6RVSqXJmWVFgkbH51GHD1eaiX8
/Kf79poxzA+yJhSR1OCorAqz50oktX21I4LmKETTEIhpTf28FLf27zG0HvryMkuy
kXJXcUvycNAT2lIkSL641RLn/3qdM6k0q3mAsMGfJKY0Ng0VdrgELDnV0vc+MyU6
DBBvNN7vgaSvuIVquzX/h3yTH8XPJ/7ikuhBEu/b5b2eCiVCouRfHkAQPJZ23gd0
kO5Gd2wrMvz9991Wi/c/2fQwCkXuotgSSSbpZONCeSipT6+py9/PkqTnAdTneOx9
on0cQmktfvYbaVTbd2IUj1sb89c4rVsoGHOqnIvZJ1KMsR0YIr9OsDL5jGJzm9gy
33RWkxieU8FiHHGiXBTYq4KPb9Oq2NkeCzDJVUmXd00MXFlR/EvhHmLNeOouJn8I
/BUcIlG4VWppyqxrZEsL/wN7uR/9ON1FUlm/ixKmXM7PZE7qHkWhTYubrDhYOKma
fwqc/0ly9MhYS2jCMWiUT0BaLvJYwqU9gzy2L2Ag9xOCLgScpLSme7URWmh3WWrh
keMuVoIi37vJB9ivet6FLfxNa5HH1dT55VQuG8mxoN3Rp8MjsF81Cle8NvZpv16E
coVLp9MNxoRyiOwMIqur/iOT5lFxArPi5aP103xQVt5I/7jgNmnmsm/HdKqbgkLk
HRe6F4NGaSemtmkx1jk+HfCQk4whD6UoEOXojuQPHEQ4aV6hxyZM3nGd1yf3bUL3
3OMLxZFPN6nVtpVf2Zx21ucVFa72pQk1GXgX/9z4Pasp+pzJhzJ2yfXR7RRkxDP3
vXl8/8Jl+EXTGHEbR9Yd5jLP2Lw4eHTWcRxXXCMI5yV4Rr/a3Bs2g2W4lTCE/aQU
HS93tHEZiwqua21Y7XdJ4uMK//Wmjmd35wg/y468Hq+Rddz86BGCLXeWaXkUfTmN
1xJBDQJFg47SQwSVNHy0mZ10buHovfgexKCnU4TiRyB0U4HCNNWW9mcnqPvmlij4
Xg1LRtm78GqocmzWx5ZRFmQyUADBhELA4yovobMolJkEf6se96lhGFSLVMEB9MaC
qGZhXeVEigcZf5oRPlYEBApTPZ+Oq/ayffXz79nM7QuvT+J5jkROHg1uN4wdQo7d
S6xziTBVMJ/iHgfm2lzQze8/Hb914ABAVvCTVWsX7WmggewByz+BbguP8DrIUQvT
LsyiIFcLQ0X8L2oQsyaZdMYR6yQoK2mkRgHKKWZcxkjPt3nBg11PlbsI3DjofBpz
vAxQA10+C4a4dCSeeQ6CZI4tq0Dh22/YmOUkIEQvnCjCCwvj1ebqTVgy6cmHpcQe
WUt1AjbKC7KOlDfrYeyN8/0yjPBByTilXkUGGck/K2NvreIeOOqUy8P383Fm1H53
JSOckf0QS55RGaLSCy8cgulPMZaP3jAZeRwxc0saqpWTBPw2st3UsO5IWIBgb1Rj
f6LDNYNWRRV7MpS1hHlpfXLSzQEhXm6+KZYLDVfbmqVbKF9UHD9GRvpYsK/55WTH
uOEmh8CdkY51zqMxIJYzS2+jjc5penM+HzhXkg7J+iL65WMVzOGUvE/mhBigBei1
bnSHl1zDQuTJgyxOenWYLzZNCOpSOIR19+6rQyfO4fREXRlQ33BWDzvKJ4eKKG9s
tqK9rtkOWbbWLLFqQ+EBKAF2JAqKf32Vsdn7jXM0yAxsaJiu6qcLRojO0aUESrJz
h6vYgyYx5XNzMi51+k246y7MemMmVBDBprkQO//Vg4bLl21vauGML1nOg6qxE1zb
0N9+Dymdel5yCO8JteUHzzBZwcJzA1KA6GmBDPCcejA9EDZnOU1sihB4+8RFr5iL
pzsbob1z+ra8m+tKd2qS5ndjRY6+jQaiCEPvxrWxUbLkezQwEjQlKFY7TmWwlHNu
kgMSPCvK06gS2c6Lt9S3OKAT2h4NK7wAIUMPx20QBHN8ImdSGXlVQZzA89oE8KZ0
EfVak5ildy5gfx5e684KUzZB2yuOtXg6a3B9/gLUaWbZ/9uJzwJr3JT7+f58DKgB
6lioIB67TI+5bGrTVmzeZ5wTOrHPcdPYMOaIVkH+Om8ESlZDNx+gB06V4UkH6XXf
0gdapncWLHCaF9LGjcfa3/bgKlTl2pGTqzwChP3FlMfBbsNkIuwQ7WrqEcXxCZ3Q
FVMhcIjzf9HtVBGqVNdMOYnY6MKOupqQ2rb4rtMWBLVGZ7IQqOvPutWgGKwl+yTx
jod2yis1bqofPIHLjUn7bhkg846poxIFbljrCCheDV7gJLbkfvUQC4sZSYfiLzph
iMt4KkrsRIEXePT/kC7e7DRqxoCeedqsQ8jA1w6jbdtkuC62UEd4iT+lWxAJ44jb
WAjjogQRmgDDaU8ffUfmUrOv7/q7Ipa1PTPwXDjuYHPaTVt90IWsXZiDwwH1gbih
XL+8ZJl1/mmztc09TVwwHiUuSorIi+ZbfMGy1oeScVKY9ISSnX7arzvLdJ0A5Nlh
n7kRBGh36Lv83+HGz+Xd8N4mlTPQuHQuOmvUmCZYnv9JQqduODcRt4wQ6gBHOchx
PT73Q7bzjVNlTDrIt04kz5HFzwp7Tdp1u2kLlo8WMDHoPBNTqFRuPm+v4/fF6MU1
J9kD0Po9Xkl/xzBvbwX2C+kF9P8IukyrxBFCS6NpoutuT3BvwpcN7NqQzg764K4/
URmxGjeggN2WvO6aih8topjsria8A4VE7dCHbLWYY/chVw/5JKjZ//wfdTQQ8PxY
cTqHi3cx354GaOfFzhSi7je+Gb+W+zEKUwfwfeiIe3DyVd1iel/Y6jkcY0faeG0j
GaHaXloQ9A/dOBHyUNqCPwISZVHSvirn0QpYMYdgsqFaAqkHH6HJCJd1Ih44in/U
p0kMQ0VUj+S4aLWyMJUPou433nklCM//Vj89UCL6/m5VTtMjk43PaxhPHlZM1HJG
6Re8D1xul1Jcg2EfESkZ57IXWGkocKWi4JFQ9QKaytfLL8pwlHTAkhNsf9BhXg/t
jiGwF21y9j8uBMwVSMyCK2h5wIXGW9ddMiOnrGEV6L00NH27mg3iGm1qXz9iPduh
pNgQ7Spv7EwlTenCqk+VJ7yWt/zfV9jdyrd+lu9v7hSj6NEhLGdKy9vdjvGLx/Q6
Q+gQon7k8cpuMA3jGbcqC6eQQIyUCqIpWtWu4VDzDE/FXbHisS99se6MFvDutV4T
QsRzDlghqf6Hy/46NzCNhDVO0TaQc5jBdzp66QRaoEhdEdnW3ngayINZ7falQ5wM
9fn/+3HmS0TW8GiUXn+F3qXXE+WPs9Y8Ccvg6Ygtjey8BAOAhCz20TvAONfo+OSi
E3RJU57+cKzpCEY+wHZV6eTIMCLAbSfk8a+nj/cdBbZ/dxuaYRZwGhDu8yrFegL/
MdZXSRFZCQ9NPPaW9gx/7Z6dWTxvWP/0+6j1C9pLfVfvWUlSXn5OgBp5uaaLF7tJ
fESEKPfVfmxxe/9JZFs6BjUM1yK2jG3zHZPdH6D0bWlVHQZSQCiJjnykoQ+koHuG
CzWA9/L//JhiXyLJA5nJdwq5HkBW4rgMZk0uYAUKkqKQKlj+hftIOtKnWgfGZEQI
DZWXtgEYmSi8Dqd0cbXXb9zhx7M/ZYGk3huGoRPe4WhAt0l75qLIgjt+Fu6KQ68P
`protect END_PROTECTED
