`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NIyBnK9ens68XIzZwj3U4vOh/VptYfY1Oyyv3FTJH5GncEHE1v2u4OVikri5ItRP
PBOpACliY/THKLHTXxWzhIyH1LfbTFT+fOBhkUWI21JI6JRwQtKX0xVc3nBZUyLu
raLnH3787H7fSasO82V9yXdGbivkGI4Z5evGpwpMuLH5FEfDE1HglvKKmT4FwEpF
iZGtu6JycLFUakIkVNTHH086gtYKhaWahNZfEnQO+R6/BsfACOCOnKk1QSjU4YXW
RbKCxMSxqOKOhHQLkCqNliu7InXYVaBBrligkP0zzvB7jEjWOVzLJNwnAjCWxdT2
djSAs08H3R1Ewyiii9vYpQrlv0nNWbUd0ZYVq4Bf9tA/FkKs2w0ZiI+y5NmLDS7t
ttAhyM1FtiLg+bGbhE31oT8QzqrwO/1TW6yPA/i7+zsD26bL/oBWFNh6XZ9cVl/M
+bcJ44dMJMiOJ51LYfRJS6ek1z4ZKnb6AS9L4NK+ufPCdbdLXGkmpzNt0fbto9ST
cC8p5K0CHtg8vFxX4zMWhmWHWggIR2sCP+uBi4JJzNCr5ByRMU2YpZmA3bBWrGEP
XzmYA0V6LqOu7MQnr5vA3eePgG1v88zWDvTfvu5RXIJpro8muURYxNa3s+s+5N+5
IZ8d4fpu/GY8Q7jxzTRJnqpQLqHyo+45z1/3hgA3sKwuz9N4h6QXs9HSu9jYM19r
I3tSRjhCd1IkqcA53FBoE7eaQCKZSiREX/eG3EKdMu7M7TPg/I/NC7WRpfd81Sq2
7DS6Msb7tPHwsaKdcq4EG3ICQ5aM92qSVw2/zVq+b5dbGl+VRRTCzzBo5kGajDhr
ASyPGrCFMWJ9q4wBvet0PoiivQo1AWjqHR8F2DpiKxtvTBqFeOHVR7Jo4aEpd18Z
xXqSDDXYdiBLVaSl27KevXBKJxggPq4kvFNLmeNzYS6jg8DXi0RlEiFdXZA3SPJN
2SMzKa8uuOJAAi6dZElS8bwPG9f++TiPBYTK0Diyu5aPELysOTuBYUNApjQxdS9I
mhu/soR5GS5+i8DjRbuJMsWiWMZTbZD2PsRFgyOY00/wGSQuC0w5OB71OkKfg6BC
QHGPSEOaFVfYttNHxB3OhVIRxufl2qRExX1PXd5euFpvityVy2dBOYj8JmePikKN
TulVZyqTBOq76F2AHVpUR/IK/afVeqFOXZvBOD5eeR1JJpitj/63QG90s4ruVxhg
YBH11d6o2nMiB2BK0/YsbGDD+X1ZnuEkKnqHsZERBt10RbQLl4j0kvV/OLsCFLLS
vQ4HeV2v2wfFOkrXji+H0hSz7y8u6NMx0idj9INEZtfpAFyXZ1PDESS7Bo0YJSKQ
P2q0eWBPlxnZl6JFB9kLp7QpypK2crlKyhOhsg9N4GFPjoJVL6JcT+2OL5/rfKp6
4AwMNXHlsgvFLi5ut7BZw/L8iZU7YXeaIkO/8X9FHGtbl/DBI+swp2PBguO0YsEn
aEuxyrXxW86zFu1e3m2uoRpZ8yc5yxBTTzbYvRl4mkZ0xKKQuWZsEf0oPC+EEHtu
PpekYUJZu9xKbVQ2xRGulI2inOT2O3fKkTwiFcoiabyB6mKi9eXMLOHk5GsH+4le
p4L/kYhsSbQiF4p44fp52+xfxvtK3+xrHupTS+pVKVX5glQzNy6N06i2GAjsTJqp
IJ84olarJ4bKTw2OWms6c4EC78GF8a/OxRNsU1ZDWi26Zea9PJ6gz3Zk88Im/f8D
qPfMvkQ3okhVaAMTFCu5ztmd561Loysnsf0cT/7qD2HJAmUKyGMueUYGl82qVJFJ
Tm2wXplvibgC2xwpQp/GptNIe8q2B7POpO4kDdtsvQfMSbXPEv2nxKMGptsVAByB
dd4K6+g+uEJgRkFHE53ys1aCv8aCVlhF88AOvzq+A1UpDloXgb+vfG8noCkneF9S
IjNPvrP+WnBjoHr5nrnEe8AOi+39owwujY6vUY1zZlnx5e/CrJikqQtg44CBqXZQ
iqFmVW0tZYMzDUJUdCC2i+9gp736c9e6easSApA3Ta+UaH0rPoUUtWyMqDUqulmd
eM1x+zr6rutQSGcAxtyTunHjLFBUdhwfLNEIwq9guVF0acW8Akt4IVrLewMuBhLy
ibTN1lNJcomWuGtuLIYVAQbrpqC12unO6w/C4V6dc0I9kZkAtAWeOJaz4fqRL9/v
g1wmq7ISSt/V67SszpgaZbVdMv3CtmsiSFeCt7ZHWzaziQUOaGO0PVSHhFBt29Ab
x7zb0lUYJ1LRET4GV4AwiChUuKbg1ntQ+Hq8+CGvSr4HadCSi5C8B28rrFInLb8h
F2PPfBdGItB0Eo7nZ2fmnaXhmBBrFUWk2XuGOK764+gsuvT19EAN0w/5akx1Krrh
oVxxdwJhnbW3OB1brEN2FGL0chXqdjevi3xm5YHGhC7bl8dmMzxLAdMFYO9eRcQz
Z87NTrIvN4eYGe3c0XahGDIQM2giuDbF3IM0idC0J/JVNb1JQccV927vKiLTD8zd
Ng+IRS1NkPR9jMn6tce5DTAOsqQuLMWSDzMrydhArQUt1HH9s7z09YDKRgva3kOd
KGOnfCR8VRtMUwxxz9z1376ln0qe0oZeDr7xOje9qQS2jzGgRNX1jTWzvIYTvdQ2
/j0OBtZRGAGIfymvRYHOL/jjZPOtrQ+S6vMnIGiGuUazmzEgkY26KQiAjxsIK0lo
rxIzFjg+2fFo5p3mwuqala89K7hcfWEElpk1NZiYBmKMGGMJVNPtpkqoeEm0js8/
MxVD7rF36sefFNz8fIg13Q/jozFKsxBFsaZhF7cbxKGfnK/W4ODAsfO8NypqZewT
788ujpKUIy9HURhSANyfXy9PatK9DcLkRR8r3vpKcIW8ezYaNwpBnROPEhGX6GV8
Ibe01iqUrdg4VVUhIsyTtDfTRaIPCQW/hqaLnN0sFNUG8vzuj/mP7EVoVoACOFlO
mQrDjn+GdrhmhSc47BlguijIB4YWyysfT+oJqrMET41KjNFp6WLXFYbdF9Iv21C6
nDfvwbZmOIj2AUc/pmOi1R2Fxijf6gn7Sjhz9BbsY2hYmZVCKfTH2gzkltKCR7+p
e3HIpaoc9d14f//Kxv1PcZqJc7RrOZTw8TEdXa9OliCPnuYPbHrPUQErLCkMNXtY
z658aqtdFBXn3lEza70UjaaZn/o0zN35wNMUDE3uwscIW3MAPZrthLrNZlKTTXTY
cuDDMKL9SeWRXrzB1jwk/tSZiVN/BV9z/N/keLCBYNk4gSh44+sdd/GpdK3RuMlP
Tmxvx9QkEWU7gk/H811Y9b04KQ+VB7IgbO2PG0zqEFbt3vL3uM+0kAEcaFPWEEZh
H9RpAamJDwLJNmz/Q/QzO2bAv0hcoa8FmcxNXFeWVha3VJMdiFppBzP48NbwGTt6
Mp8xZUBkmX5qEXAEUm893hzpe5319/d4/MfOOZwyblu3Sw7zRtO4tw0oJMktbZvB
XxRplbqC4DElOLyXDGLh3yvVAx8kkdMGz144ZiD8Oa94U7tPC+k8w/9aYoykHzLz
`protect END_PROTECTED
