`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mAs2Bl8/HFa0/TSFdPzw90p9yZzq0LrEUdVFGbzV3831HF0CHYzP9c1PvdLtcIQ9
9tJDGHid2TyzlbRfZg7pGTMx9jJ6SjEOVVGUbJZwA+iMneCA5M1xU3EJnFvKLELL
WlB72kMPQwLr3V/BO01sdD+9CPhRTvYJi+j0gfYGD5e/HLT1DaY5OH519eyiKlT1
HbtiqqrCtsM1PrTws6ScEklz5sJ65BZxLrP2XEVzs2Hucu7LAAKIA25KnYGQnUb3
YFn/bm1zS5Xtr5Zk+kApHTtzKpTVpFopfOIZD9Nfa3h3AowOorHKbKUg2EXdPhF5
wKfAwzztNvsHRkC0g/rgGcMVzTJPoCnfbwxQK2qc0R16EbzrsO+6ZwrZaTRLrgwA
7i23xf46PGdTG9IcTMHCV/2Kx/xE6dEg9CmLOXain20ZFdKTAOXZs2F/HDLMgKoz
A6w3mzciTNBfB3SRfAlRh7Nrio5nRcja5cB8yFfJ5Lj3h6JX166mBgI796eGbTLd
j0W9wLhWFDzOvI+Z+501cCZBQl41Zr2k2BjJ61TrHhxzg7R8J+6c8hIPV0ZTM4gK
5O5vakRy2ljDus5bT+ZZxk4Cs29b89tBm6XQzKRcYEw43l1ISfth0lPYM2Z694Nv
ZoDQIccRSfKRJmaiRz5nrwS7rFCrQ4OFKNhEEGUCfov8m9aodNBKLjuwTrLmFaEw
KaHd8R6kNWMDlvRVws0WR0H+9sruSjAL/I8LW+/+tFJdf6xCiIcCy8qDia4BeVmp
DkFW8msgjkg1evQrIgh3xNTjJXqSUVAb/BmTjl+3vm+eZXfVPoaXr9NbWr8TZml/
LaqnZjGBmXgD4MoZRhKPq6rgk7RGQEna2Y2wRZCFERvXmSoKcJIPq4tg7WX4qgiZ
eVXpwNVN7by76LQbUEzI2raG5GvJUOJWFFkMEMdrGep9Zl0oCRwo5EKSPP4JJo0Z
W5xHhTkNJyZoYQGlDnLCzSnc1gyqVJzDEzqBR6X3fdUjqW+qKu1/HRvdwVNZ5mN8
hF8G0fXrKU5EJ7UwoGs3ttCE/33gw6xEYHYN8ch9MHErna+S5N8+GArJPaUnVAx7
53j1iOnNixdLncUKSRkeGrAQqaOi5OBqy6JKdyqdezQyk2rJmsTDWuPE0LUdT1lZ
nzl3VjUshZz0Uee4NLX9tFc9m3S/IyVVX/rL6oz12lQeVsR2sM8a300/V02HSH6c
14C73UpIGszTBuOMHqf/kyfL5s7cX+FMpam2J3BUlyjJ/+RgHwceM+xbm8ZIUVu3
Bq1rFkbMqeSTyIMubJrFDgqeQjq7I0uJWl+HNIZCcuzqnsKL5XinBy2fGiZpYTOM
vr/nIoER7OSX71MlrMtNgND5oU4ZJZmuyBuaYBGDdirkzuGtM5OILw58xqtaJdt2
jHJJTtXKuFHlbk9l6q/mxGPXYK7dJ2xupSaJtvmPXe9GBYg2wddrPD1oJxau0+A9
CxNLseA9edJckjhSr9VGN2KKwYTPjlzeHwnZlEn5zmDpgU/gHzxyHUvGgWnR2ikf
kCRA34czKOA/LWsJwajoQJ8RWfbRF0wRHGFPLIBytQGcvDI+neQSr/K+G1YDs0Wv
UwIxAUgkiLJBqqQSF8WATTuvc9UChPLTpmOokMeOoxJ5INUyIrStYzHUjdWkAWYc
Fa4+J8A67NxoX7u3AA0fdP2tPTkJqDIxuYuKGZdD0qjrDR4tm5W7KX0v5N8t8xUe
QtnJG94h/AqWFD4pLigdWdHzX96HEo7qlTMeqETb6YYlZVLyd6ylUUhC7x0PDLdo
bfhuIc0Ye+NwdrEIpIfHH0wJIPZhB+6SEJkyGEXRERRjM2/lhTpUKCClqDEWyry7
FC9h1nrQYgKqYE2+QldFF8iG/+tSCiNx4rA9fTLgNvpiskqPr/CTS+aCI9IBvYNR
MBtcubUgg3QPihueXoETZ5emYIhxdh0Zo0OS1QM8qzQau9XCvSSCIBSTZB5DG98H
0RRJrZXmfRGbgoCEb8Hui7WpJMbDfIZIliTCJ4sg8jYNT5Cdkq5Wl/ijpxQaJgYe
YtO7ge+1pPsY4dwTgJwZIsdm3Qj62XJPqSIwAkIqWtQLXv4Alff1nRDGo/sMcFWv
rNA6bvhf1Hnf+dtAoJR3xi3dqqrgOqjEviBFhuVi6FJjrcFnbtPhcrYXnyiRzrWg
NMHGdDeFQGayuyjyGSoe2dGOULU9nwhqvqI2d+1fVdYlRcs2eJeXHiXFw+ozEtF0
jsAe5fEsOSw9DjNbFnNCGYTyYCpIGxCJK+Fl/A+xA87YG/7PFXiHHMyjk/Q8KnoL
tRExxGMs5DotO1F8Xtqvw+nMcR2l05SVMNebT2638PBNF8OUSCt9T3AB7hhUkWsi
oWfGIT5Rh2XGL3IH7CzkNlmK4eCnL+GO+7cLjxkEKmQgldOvwOisxIOWLxAzwdnq
`protect END_PROTECTED
