`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
stXXapbpWCTBsTP6m18+bUQqsajeJnATRRaADQj7Ef8y8U2lZ9REEfWcjBfkIimv
AnztXJiJeA1rwON/0a/kqs/o6VqjUg5ulmCdmHHsKPre7Eyb0CqATIQE1SZFlSmN
mzmuaJwLc8i87IsB5U2ryDPgTELljfKyy4BGpV0DOG7WjOEdH/6X1eaB1t81ynmZ
IR4v6eLGXk5Wdt2uCPBkO8nWMMxRdMy03M4f9P1cvKVGVzIfEv91HUT+tdoPRcT3
aJ5fREdh+8t7SWOFYqtrZ9oqyp5dZzZ4gcrgfHsbSoZaCrmcTH2tRA2pPTm/K/J9
zV59QZJib9672wk7r4egZse/FiTYKYYFyyYzlUSqg/vYyLG++m6nvb918reANnJb
vbV14hHsFRksv195MRcTJZK5wEQlvqFb/mMLHWqSihmxJUeif5FX/WE6aS0j/pm5
cSf/kMPmjdGsAfiWxO7yueyf/hncAPKsE/olMTe8wi00/NFkKzkdHSMHBsVSXIMZ
u+Av/JSBxGR9bv6pwQHp3PBZDd/pIk7AbSiiyonk8eCNmuNNYMvKFkBm6EXSnQXj
BurZBGHqX+9D21stw/v5rmKsAMcciV1784GnqSE1NNf6irWo3xp0QagN6WIjeDDZ
JrqVFaoM3KrTosBMFzqMx0VpG/hy+8O9HVSqthjTRzCws4BaUAqw5uuANn6+im+c
S5ysbOW3TIy5nnOHpnI4LRjq76iFh93NR8W/SP9RqFSPRhHxxWbZ2gmxlNbX7A/5
y1iniHTnut/P4LWCiaQ4zCVYhTdZPH3U/N96Dw0mkDY4LIfGDXeuEbwUkAuju6cP
pgEtM5oXUkMnrwVDoAwRwdRY1RFM7/qQUyJMAMQyQr2aHt60A4LabWiKBQjH0Kaw
1+9yRvIpJKvgPEvGMJ/6jNL0PhJsSW/oPTAcy5k9rCIbUzta7j6nJeat498EzdL6
5kvtgRX2hSzTBa9vtuNKwJWc436JE5G4zEcRYd6HzOdtUAvfstjSrGj2FE4dgxTT
ICe+JHHlKkr4CpMhdnDTlLYa5DG/tVZQeA6wjbtRBi27tgXn9bhHj1eJedrNlwHK
+AMRECUkNn2ZVnpvXMNnCKDVu89lVHZLntvuFSUDO/Zs5aiuecgNh8MDBYT0Moxr
bb5Yfq/w7E4eI870blkYVjkGGq+deWl3lo9wXPHhdiFt7UhfNq831Q9cJQYNIiOK
2CMzg8qOikZHgl4RfvqbK9/OW18mqUrXYPtYYjEXytOvbqo/zgT3VCFXcEze6poJ
OBVXGgdYucOl3ogAOox6cHKNr5mCsgy7tURBPBzZR2s97ouHjWiuvtexpNMj0pWN
/2dY2KpdQjz3Gh1Fyg4Y/6xxwq3+fHM24OT2qRrympvMpQzYE7wrdws1RjiwmAsS
pp5PlYashjSOgpZ5/3l1rVB8bOuBgAlzDMtRR3CSMCiLEa9av75xTDWPV/vgqRCb
fKqO32VDz1PrqhrAudyIeJiZo9HVAkSAzxU4x1VDnWNarFXYt7bMm62yVhUNt7iN
2B27jDpsoxna05k9LFsSlOZ1qxxJpG9vLlI+364Vf+d9Z04AUweZkzq+UKbejedq
tfCNUfA7ehQ/RmcroEl6IqwAzpEQkUdeebjurzp3kI4v+vWGyor2ppONDwoRO3Ne
/KX5wKSstzzXZgfa7jDbXORNbVh8yRYWrkDIquDZiq7+N3bT7U/N9dUalVIDRJFA
R0IQFqajf5d78Pxw8dJAgEwMd02C8vj2NhoncZpA7XgzKv87jUQy5No1E+tr7jVz
rp3+/qXHrrN0PExcYFQl3OsqHP5mRZic2YDwIn81UgmSGWIZtaTsriyLvksGGyKH
X4NpJRvioZ5iMAkfU+AdnASpiFqXdi7FnLZ7SZA54THOaHBCyiTGkyN312cDvYw9
M/eiDbHBxqPSkVQYNgO3MJWW/rE/aPcHaVusZjDoaZevavLNO/dMisnjM3QzaB0G
2pdSPBo6X3IaSFS0aGEvTKRvRj8glPwWvyPePXsrrM4EJAa41LlH1UtpE1Zk0JCF
JDmXGnMW8qUMUQ8Wh0G52U1wWtqrOtf++7/HUMjoBLXWVqSOd1bV/UwDWhrtUwxH
npXIA+uZuz3ntRxydr5qggr9UR6HZWaY9ak+rH7Jllo=
`protect END_PROTECTED
