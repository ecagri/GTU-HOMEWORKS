`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YIAiRSmQWi4poVP3LqpTXYeDaIqpJCZFva/bhKJz04SiyOwLbhLRg004k7esN3AC
wb5Lwmo/QEkJD2l/JdqI/tf2dGMv1b5P/X7AHIdfzDEFJcbgxQ4SIbwFlkQRv12p
wjLt2Bpah6KLUSQJDU38lwEojca1LAg5RutbDeQNK5rSlzsIfvq8tpsZw9OrArb1
sdI8gWy8HKa4jkMa0F8WEdNp8sB3VX7/RA6skggyPQX+WgWV/CJo9otaMqT1ALJ9
DAGACKIMmmpJZGnv+RgLo2AcFzSA0zU2ZbDsQg8LOZwlq49shOEsIL7ElGat2pOl
nILLfw2vC2XgkzGITAe7RjQuAKYpD5o9u+QjsBa45+SNiA3F76Hk68K/Gh9r2MTG
Rivxs6ehevW6sRK6P3bfPoeHfjkQUg3Kp6WIdoGvBphZWsoUENB7yhuZICvpXJ/v
ajOQhYhGnMVkPO7zPnMSBVIRPnxf3doMqBEBkUphK+Ulr0EG2lOVX8bDmyYdO1DM
ZJQLw1b0KEc0octN4F4biYmzIsznVNDBBkZLju9o6Gt7+Exyw5aIPytpLOpvCtZW
py3gDg6PACmGYIGLcJh4qlEnQOCxv0HZwHbfy5RJdu38S+Cmul+GT+EO+wzQrwFY
oqVbgt9SqMkJ9P3xQf4NXH22Lkab7FcrWG4JS7gGBq5x7SSjLxQXTjTTOtI2HWYW
`protect END_PROTECTED
