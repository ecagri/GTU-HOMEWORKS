`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7TACbRNnSRcE5/GNYmcU6XQycIyJhwQcW1HpiFwD3gtNPjO6zPYS7BiiNjegMhrf
UinVqYkNifmLBss8z/Yn0+JLUZw7HteB6grjUd58G2N8WpsK7ytmhEk59k9NK6j7
pF5aJEq5HD/8q1x5yzSVl3sg1xWqI7q8sbkWOZnKdrZWMc+2MyiW5WEMpv2iVRp+
M4lFUddeLNfBK16kaJYMEDTwmxuX+7r4NXBIGjVGR1Vi5PlWhZFNdxHxupi+EOXg
9xF3OASdyR47aHJGsb0YBsgitTivizTbPmfDRchg21Rgxfuh82osHGPYjbzwR/S4
q86BBv/zrPFdxEMVoicRPCxT4TQOvD9tVqs6qL72vOjv9/tCWUFqM8B4DKpqOaAR
WAjP70OvAKTd6wLxxtmZ4FWBnKQ3fPYw+NuKFlJLRHBXK3/uxQGaVIzinHfXVISR
ZRmwzBM4H32/VWPbUYlgyw==
`protect END_PROTECTED
