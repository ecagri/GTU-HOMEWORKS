`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AoVYbGB6sUnbwsNqx1PGCKGMz97hGrI+RMJBsZPoAdJSEowFgkvviCNeZsA0ET6l
2TwNi67A2qvq69zl2Ok64dqTaIp49Cw8/lj2HTa1+6nlhzlTqXX44z3rjxdSv39f
r/2nEVYQ68Ja5PkPHwHwn22HFwuEYwIgfjEyUEteWu6KNqe84M1DVJIYHbxucvvI
MKGot4iD1pQ276+9fCL8tSjCQ/noGrQITWluysZp1fIMPx1n51e6hgFc5FrLFUxV
0vXI3TbsXKjKjaT3E4TNBgMfxa+HVivplY2wi7q5iHCmG+7OG5Absl7htE3wJLVj
jK68Sj9J+lZltcLYfFjkF9FVKEx3BPqTG3qdGh5kiXR1Td+ZPermfj6R1k+h9Bc/
JI7sKmpXiK+yOAPIQ7WUxcEnZLkAGI+eUoZumM5kSEIn9qJut+RMxKywCI8Rgk8T
icFCR9rHQzRlR2tSq+O2W7BzCIi2TVB+Reamy8wVe0pTR/kJB54JwEiK3WiSVX8V
pNe5xxAKZI+HkV0C5Hgsh0srCS8jfi8bfxZ/UPSUwRE=
`protect END_PROTECTED
