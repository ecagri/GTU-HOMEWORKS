`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZZ1VUgVCwNMJW7M/xTVl5VDOOWHkpwdFcs7fQgiJHiindrTD0JWIpA4gaF6Kf+eF
aRhbXlzoVDUP8sQIOwVOEKOeqNS7y3hsfZ0bxr0ec7/tVqw0JUhdFcjip6JyvOik
EIVM8rwaVvwP7yk3YeGft/cqn9aMkZp4CokaR137GXoZ4bWYCNAUTy5UwMgv7W0h
j9cVqpJ1BNNkm/ptyK01pKq8gMXI2FJA+fVQfo24LJd+cf4JcvO7nok527nbV5tJ
7B7eJpuU3FXjPLy5wRLoBA8lQeyGTeDbgWLlOdcQjSqcBEcX+cod3Gr1z5A0qqP6
uxePRPZU22htMpWWACrDjLwaSNXRRO6CNfQVhyY9oT5i5K8+S0oFpxQTXIU6lgs0
Nf+7zf5gGjCVSZsYZR9tYWFeLEWCYo3UiuWOGg+QXtR27B83jurwSGal7ba449ig
7OzDc9YdRM8dfcL/46UKOc/ZLGB+tR2SpxvgqU8QMsWojVPy2N1TKfqy3iUZW0Nm
RQwBVkXT/dCf5Couxf5Kb3CK97atCLNnzwC8vjJcz4XEDo4xvQ5UYxyfTfDI95KO
gmR92xPAV+45NLE5aoPRB80vIocLpfkCeXdnIrEDRmtzc3dJq/g5AoU9XbsBKyi3
u3olohma0rf6yWwR+AQdopewlpdd59fjdYm0g2Q2ibBa4rtCzB817VhFf9IJsf12
1NamTAuY+XdEHGvwQPmF3pKZssyD+cKnq3mxPfXmmXBBNFAycd1FlUL+Z1L7ZQln
4ySb3dUzGWKQsVOU+SSLB2uHoIOJTFfYPzFaDJEQ0LXkyxq3wB96IV7/ryt8tUqu
+o500Zp431/qDIL+PoA9/a45vgQ+RhBXCRo5zJVIT9VtdQunDCKpUq9v9/DyeJcM
+EbbooLGVH53WniE55r+qCb6+DNMuZoZEa/fYeTJKmqMZk8LdpHe3wXVcFutAHc7
MoEDM5qk47btwU9DR4ee/AcnMNSOZ0JD+r8NYxwCTjBs0wTS2x6qPlK4E3AZ/g73
klcft2qnZwWWycYvwXjCJ5U4TFTnj47vc/q00VeJH0fJlV45tSlYWnVBO4j8XJQT
Xym7tFMHdgNUsENa3EDc+AT8jN4cEnEMq82wzjL1v+fHICyhdLtK0ax6lmwNj8zL
OuvnG9nrsv2yRdlIINg/fzdhYUD0Z/I8vISE6q1yTfHjK2/GY2zY4/DB+6wMAZir
bUF+Ee8wu5+5UwiS0nIV3Q/4Dru8MwcO0gO/UhTD3/dMsvdN81PAQls17tmRPhAL
9cktilSLzFMlhIsmfrZYeq2Xzj6iKcgXwbDSxFzxI5YiR0qdE5+2SzvRxLL7O7c3
bBDZRx9erpRt7wlWkljkVetNEQlPj8X3O9mtwIFVY2Th507Ta8eetc3g389Vf0hv
FGcv1MztTNnwus/11bfB8B5dgyD5G/FQyw/kuNoSwYk=
`protect END_PROTECTED
