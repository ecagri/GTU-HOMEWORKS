`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lOuC9ZugViGmh8PZVL51NfBkgC6bp0op3B13E8mS5YceF3BkZaNplUC9FuLak/+c
IYUlcv059vC+3vnWjxNH+wCQ/PjkdfZS3iogjqWHNHJeqv7cjFbDi1/vsSBjGzF2
aRATJYrUBfDi0JpHGgcwt/fguFrG/QW4FPuIw52E6T/Ulhlx+CB8KoSTjcF1AupM
+ZdIKA5XykQ7yuCoaKySSvR/jyLVM24P0i+cEENzXfA2Rms6hPog0+ngxznIAA5z
1T9OTLrfwdm9ZYYG7fo6+SRPBVMMDCu3DUQnkJ8kzSKcxJXXrkL3v58MnT3Y5ODi
XFkBdL7ZMAiePukZ45EMduyLbZm2ASyu03bdaCn/Zp73kk7sTuoNCU5GnsIi6ipR
owD2I64CtP344IZgV++pwXR5yeF8NIMIzGwk6Eoc8fxQB/jB7PDegQLVRVZHh+aJ
W/W/z7lqP8PYSoEei4u4YddDRkdZ4CRfHhTWCEg6TF0Ex6Gv+drRCf7QJ5eL6Ofz
iEwOKp4bnBHEf0qFmJ+KW+2kORN9slRcZLT2YHx1PpCo0Ch+81O52MRtXAEhiy5c
4NQ3/kwBpQx5Cn+g/VQUzZXaqQ5MYmT6Dbw5s99TfnTUIEejfG0a8wpUOP4fZpUU
p9oO5teK3c0Ug+1+qjCqsw4tB+kRynVIPEQfRNn9QXUNkrR4MoIO1Tnj87xFpFsT
F2jhu5ZkDlJ8W9fMpo9jq2a2UOpO4BCYzjUmA4o6w/O10rBdoAxGOQVgbEjaI/hk
Khw9LCEb6UJXukqBkQCIAtDpCrrajDYhx+nS7FiVFWo4YPtPmyo9/LsNmxEIQmGI
K1oDT21PbsrTcs5tc37mSrbn1Tf8H8ROZI+fc+mf8ZMaMApPZ3MrocSkmTLxe8rf
8wTkHMBwNoORiYkVH56M+p0oyMVJKxpAY9O5mvV54rYKoLW1RDCnqCwwfm0qxQ0e
Ql3k7WrAZmoexGyB+FgipTm4AylihWuRaghgAe4fn8trnPuZSKUR8i/rtObfnMT0
gfe/rHT6ucqBiOUgTOr/2gzLHSI70CEYfqAK3OYxN6Ek5cQfiDxAkVvzGPRZJfS9
hNeWvyTL6qKBrzPcjJpedRg/jW4REF/YCjWc4blPGcnMf46qdyfDdEIQj48AZqqU
51KOZOjUj6/yCrTtn332PU/fDYKjB57hwHy6JVnDLEaXQQh4aiNH/M3NbXPyAQJZ
qZxkPmd61SzLEvOGtcIMH2092bi/ujlhKZkz/0iUb2P+8Ng4N2JT0yHR+T9wx0Wc
fjviENk4su3bGSvR+WqGQbQuc4teCGYMVDQICCg306X/wQweEcdilP6bzPPlHAZs
joRaP/55yOG3N8oOOHsjiqSBhDbnMNq2cttw5MN3xyjLnckF99CyIs6GMP3SF7F3
9r7POF6PEzgaJHDu7sRdi4uoGUeqySt3Q/nUEhQ723O1xDbXjgdrN4k7xyIKufwJ
O9NNFouIHvVw2+8YPypGljW9t3bK3v0VbVanXp9cOgQLQZL0j9H+q0fdZ+AM8jsB
YP84+8CeueM5mAELCjr6cio1fAQBjbTikvAZakNn7jZWjtSwgLpdMFFLav3rnu4n
KqbNs/JwI33zQGGw6/L2/PnJ8IhMTM3/8x6O1sRw+Dnio7NCHXoeQ1/57jekmYSZ
qgfgIJsSlc1fpOFikMy1ZhRoNKRTz0I+y4x6UCSEPnyIeRpxgEUy8MT0zFgPPpjE
ndkyo+JrvVa9aI3Bz82YUvU/Vk2mNrpMbgSuFAh+/J2tyfOjNUPSSUcAQD2cBABF
wVl7nUcBtHoZ4vxioErnORdkiJMC5AWfWMxOqKPL3yT4bsdf2NYLfNFo/vnj5FP7
u4/KaM58r3h8V3mLpLibf4RGOxEdw7KsDCT9tm+NXyB9NCDc9nhQO5xnTBlG9PUb
UImJ7yWl4/U8DTQM1UZPrDn8j880Dlt8Ub0VWiSpacbZDsjDMEXLm8UtplbP7plL
lkkHy/Z5uSH3NUiCROB3ECW5kuJ8q3oYAhWo+h/dnuwJSMFbfen5Z+gFnEnY3dXc
vs/VpeJju2I7vzem/kGdJ6wnxAqweraPvQtWW5CnMz9Frq83e9ON4OG264ZIW2c8
06zeXK6f5u8G6GkofpMY/j/L9io+OgkcxIIGv7O5FusYl3hFXOTiqPtj87pkopci
ZOVLtb5uFCwqSdjRefysgEtZBBw3wSok9+gczFusssYv+rrX6SvYvhBGI0dMyzdW
C3pKzb5ok/6fP7q9PDDf3I5M0Q7BmfqwK3mSyn11Lv/PoH/WHLz9j/9+Y8Lm8KtV
QhHHmJqWySI1Z4TwQnt+ShX99sakNX/mB/CX7aa9bpguWHIJklrC0vlBCqjdJkUY
4cUK4W5IwVFUHAAL9vaqIc6ZT92wMGewsf/i8w5/YqI06a5a/AoXjy+D5333PkVz
JTkPqbNPFDqoKDfHYGgPqxUCZP/U9QSgGSjEu3ryL2Em7TWjjgm52mEwHilwhh9n
m2gHVnPkmkB7M0UFxr+24C0PDp/wwFQR7uve99oKXA5zihEqbk10TOQp1+0nZ1tY
KS2tD56I9CNGrTRV9wHiag==
`protect END_PROTECTED
