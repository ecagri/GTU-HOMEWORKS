`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a9pkOsB/qVjOAWAR9JbZJKTC1xqzGFYZKc2GkCdF0mK0lvrE+9ewtHgcaKZaxAW/
dxTNpDptVo0kM7awr+LL/9maTUKKM5MkgOiPeoQxr6/V2I1hurjBMJoga3D2Yu7y
e7ab4scYK4uCXfxq+foPZ9+lxM3IjLPxzWAdwKhNXjWzHwtqsQFJAHiYtNv+D1gs
eYAyHfMHms0XoL440afAgiu/yMhNEyH6o/x9JKdAz/ZcRg9fsAkbBVHq6AEMU+hT
55RmyQOhYTK8GnD4LxNuRNR7Rdo4e/1zvV1nPjw/UyzVgle224wB9xwFsbbMJB/S
ClbjXxzKs9/PRN9H+GzfczrWY2fpBpFLdbYQQgT+6P3FajAwF9yphFpyCEu+zL/S
JaVgi9PNYqPaJydwpA/n3f6A8brDvRjImhj9p+8u5efDgtJjof2zU4wZYkQpU1HP
m6MsZ7mNKrZYX/0n+un+CMZtgfgMUjlrGxhdQBxvHl9iUQAuIcw7/pxnl1ST+4lJ
1vZGLqf0/+rO5l1L9RmIlqFaYaduCTQnqlfX19hHH/Or98Dh6c4rjGhhvK9MiDal
32YC9Pa4pXVGnsjrNs7GWgjRvVI8neemFIGP7QIzHCjBEiKqm5zxmAWlv3J9wV30
vz45L1JAjp0Xw1RrssVLKCbfQcoJA0SDS9z1bfycoNVpYBe6VUPx/2HFW01hU12f
R4j3vWux0gAbEQJoPNzDglIMvCrW2yLH5pZkmbh1TPjTF0gGmkeLkq+c13gQZqbc
FFeXzy3GbaJB88vuweChjoeO+jfA/qtDgd488aOHVwF/4kqACAHES+T2b8ShTfJ2
7ZvGksm33ji8j/+e9ImotjQkobhL1slbmSVHgprLk3uQHJO6Xt6sLJDrU9SwHCeM
fTp1NexRAMPvv0N6ZIK7XWst4/hw8qx0sJkp9vhZVndqZHgGrMNO51Ej8MUcXsEV
AXNTSczSKu6uh7th36t+9ooPHsDNLpAdcfrTdoHh2IaNsFbbeoJXKni0l+eQ6IrS
8j6iD382hwb9iS9zym12mfD+uKINZUctAK7+Mv7SwZHoW6n3DDIr+JibKMKLKuU6
QVDyRW3hhc6RfAPFoETIZ+Rcj+g1eLtKrTSyykPhDWmNYonazlqu+xLIb+TU5JkR
OhX3NCU/pGVDkCQHN01KyD6zqpgAHsernF3aTX6CQNFBRveKj2WE0ARIpVWlinz6
/y3Q7s5YA07REzh2myW4PInhUZAnRBmqQ/PlVA/rNecrGRyP6Z93UOuOlCuqYnzj
AjKWnvOyPbnQdN2M0/0N8Q/PGQ2YKs4cyxC52GI8Aw7MiyK35mSZlArL92N0YWpo
KKJm6RLLaG7wvrolru4ZzVWOfyoi3bIlJ8bwLedkFU0MtUwx/eVqHGBQ675WcNbE
sswWAAP2ovoW8bEOKyB0qTLPySR8gegnl4buLG/sJJT2eEOSTIi2Cn/Iws3fYLK6
X/hsA1S/maBjsMa7oA8LrrFaWf41vMQHZfn6nb2bGqifIxF03/n2AvtaZKetE5ef
ni+PUZx5RC3XqolK2WRHakvBwYBRMTJgfdROOsu1Wkm1fxE+zoUUnELt/aXuVHYP
thdzbshDL1pY5rR7tuHWSuSFLeSdGwwsP7YH29h10CqQzyxH8p2AG7zcLM6HsSfd
l53RIvV5PK8CoLSH94FxAJGM8cZyZ5ZS+1x7KwZOuhd8VXvLKchrfV26O8ZDtYju
vhjdT27enUix2UcXEca8hVPlO+mt4t63QkurWIFa5sNz5l62/EeR0JAJdAsdaoOB
Qv65lXFsWwJ5Qqm+nZypOqRHrxG9lwzcbhyvvc/1AMsN8BAlRkc87eypC3tit0hc
DdUzKqRg31oDSgf4pBv9jKHR3Ypvr2hhkaJgwTT2Sii/iFZIwv1oWuyQ/C5Y3Koi
PzC0Ay8/aADD3SeDE0Ixdd99RoF5lGwEdJruuT3g2Lt4mLBeoUeoizIX992NRMty
yf2I01jVSAdxh/x7kTgrkBaSdOgNx0N2czH4WVhHP5HIZqK/wVyh/kJxDpogzsQw
NHRa8n4LOFbHIhGQ8F3UApIuwbAYg8ZMdKtl19wzc/hK2NcatjiLbJ/PyOnpNQke
B7IMbggob+ACehPgXvQ0Rl2AX6qT0URmuQtyIiqkuIjqOPfpiMPny4HHIi/EqrdM
dgQi0ojLOUSD4cHQdK2VogtfcUJ0aN5H8xwzfrJHwk5E5ShMHqgi3we+xXh/gBs1
5rpxZkAmo4Yx2DaNiN4KcnfdYDNIDglYRbdwdsbi7bMhWrrSuT3Tpyj6gFt+LLyI
+kM2GpXMkypISCpxFpzw9LkLZlzPeQxOJg5anCjQREzUNePzv13e50/WYkc9T125
MvUugD0YbtvTTcQf8KrJJg3CXx0/zDWDzBMbGtjDxa3EEf7kLSbv1eCUklgQ8fqN
+q1J3mnC+lfNooIlyjKX5hxiDeRyrh5dRlwHsNU1ltjXEkpILDRZskqjpKsRHSW8
QBaR+KsUfu/dF9ABhVRP8pm8AX38L+4frGfbXFWYqfRhGQIAfLzDjG7cFfciRBiH
KCWp33f9Z5wxFajKhXsrlyUYGJiKVrosrlLfaQKyS3rPIDm5oB9/0QQIgPuId1+2
IQggiXq4qRu8vA6pRlLBAJ6euaZ7p/8oTq4ClJe1CgDVXD87SF5JC3bV4vZz1Y58
AeBU/ScG2pqqULh4+sm0GQlfMs/pzq1rOZj0F8C7NpedPD9qWRsVSsO+g/Hquyos
xvUCMsTpwugsKzNFqP6TBzrc1zY1P6Oi4FrgZuSAq7d2N1vrkpF21vkJWWvP0aQh
jDKKdbKUqfTYDK/kncNMOHpx6rjIFkBhiruEr5uCArPVRfV+QB+kZ/FCW7Tam4Yi
PwMN7y5CLMbk5hxUs4VfVHmMOjXCuIdsxZSQEoPjbOMIq1WS56KelGmKAyiplJvQ
yChbLlcPnIpBmq964fYIxeBR89s1Joj8b2K5qVfRFJzJptnsl6Q/+i5vXths7z7P
Fjtn4ILFM8VMmLM2dY/n1yObKUlItMGI7rK8SxXH1Y9IYmHTn6DG12bxZtG/BwRZ
oCOHE1xSwh35oSUyVIC6kkFg7b0EkPCKNNHnY3jDiJgwEhCTrX7503OxgY5ZY8S/
VwOnoz5LZGOnCBn1vUh9WuxlXFtoGq5HnQhZ8FWZTCz8aLjxpQn5mNmlW/w+AWfE
LhFgolHc+n+48sUKbjdHFRYzummEtLl2lHblHdr7u3c/S8D29snnRhm3rGJLp4n9
ylXjx2DNPwh9olu/kt78MiDiXp8YCTrXpGvZ+pw/jGRO08/zCq4Kf9zihaPcyq0h
IzULs83k3RT3TidD1WLClaONkgBsB/cK/bf+a0o1lBATLrQMioa5RsmWVybnFxM5
JqTaGbqnu0voKSyr/mHt1DnPkZY5H46O2M5dmVSAX3OaSDIr9u9bTNGnj/8Yl3EQ
qyv41y2lvtESVAFB+30lzkXhstJBOJycs3r2c7temO9Y9Vmi2yy3JyCj8dg3gdPu
n0NIjpNwW94k9eBE8J09X9qp1I086hj13CmT2KxtJhi7OzSnpPhDwIm3aLc9Ksv3
birOvhMy04kOUIQVfGHPPDN20zehck3Uq9w0NwpCuCArHhxdwQHO/EiB9RUOhpck
J2rxLgOfpzTmTSBKnpdIEibl8XcxR4YyGA89KQ1wXdkAc0AiyXte8QPaIp2R8vdV
vtbtu4P6LIPBlnK75dh2A8Q+fwP8x6FUyh/tcjJRJXV2NjaCYZZ3D7zsqOAQNIdS
TqC+6E0CzV6xCcQM+b6BUQEtj9/pU84Kxvgk1V5okFIqDooBWG4HFJWXiIexP2xE
It8nJ4fZfaShBcV+G1oXPqUItZRAd1lgTciShW+BFv+xjQk0de6ll4+suNSgsf3m
yXB7JR08/nDkWniL/IcwrcBiS9QHTEPLn0ODjtiRcK9dOxBdwjOgvccqmJe+axjT
s2IjS2PCdVQPFS05uuafm70sfiqiiA1+hxgamDLY5ja0+HtulfQLWFQq9TmD29sa
JuxBFlZi6+fWmoLYJu+y2FkSvyIVbgsgjiImraVUfeINqJC3gUaOfjeut6EGJVFZ
6JoSG4241LB/5W6Ej81UDRm9GVym0NNJdpzORmF9/ZZFbB+yoEEm6lL4mNxHgFV0
1vF/C7xmf7d+CqJWwBhLKRIChB9V/UsUvwQQNkI0Dk6gqKh8S+IhWFHdbogN0YvF
FspZ0g2I7DR7bQFrJLqV5WOdbDFyFcoiwrqGh2HUZmnT46a84zLK2FuXiYn6mYo/
Dozk8snfrxBcryNC4S88Y3r2OjkRjsIqADQ9/lgfn85j9UMo4Ah1uMbQOTmJnvXz
J2WsV/q5+NPGJt+rdu9g1iMqzLYT+MJf5deSO5uHaqm2/9U87ghmnjpLupFNqfCN
TZ1Snw0uUC1wafNkEJ4jyoHa0H+/xyjiRsUaEqb/OLWGZTjJf4bghAY83mxI+WKD
nxI7QLmH3+w86QOvFRXND1Lzdziz7UIBBzX42Pam0VsPwTCAtacTzeHypBSE5roI
NoKNZar6IlhPhV0rCIYu37eWwvni6TnkYZcshdR2Ab0I2XTspgDaXQfBV+orcqH6
sZLkA5Hv6wJNCD9/7EibkYMp7unOxhBpopooPLJQaIoI0bKk5tSAV3mP/I16gNfp
BAtLx9SMyOSgQoyLQvaZRU6GfmNdlXxkLi4o9mQQ4P0CaySw9uvSRDx80/ajVbpG
mhyY7Nq4wxb5jXtVp9tdMF+0Vg3KQxjYxHmUbKGUICq38/pxDxZpJSmrXs7T6TPS
NpdIWKJNf0tvH6626qnwezIORCYDMN3jLmz8W4lJfrmmg0tdoU2PBX/UebE84jPI
kKGTfCl2iOURM0Fm+qwwt4rJyuzsZuWZbkc9acUhl0+l+PJRbA9I7ey/MezFu2G4
hZWmAtz5LEFndyttQ3KWWeaNATOrSd7EN6WI4cAjJsLSIlrUEtLWJigzx9mt+c+H
D978YNc/R4vM7KhakLt8B7DMzM3/tD9BLE/CprMB4x6tcygdkxPhh2VBZowSLZ0a
gEDYDhxAnXFgKtCgrVJHaS6CIsCrU7zZw3sFCccVaeQknSuw8NXS1W56bJGwDnd2
f97ysf+PoC1jACWL6TPLmHHAZnFT58uEqufGGDggXyLhWDXBHyToJVMZ6JHcZlV5
sgQQ5z554Gtw3RlfmK/WR2dM43AzeDotMdquy5DfgaMRaKi5XT0ofOhKZBLxwFhH
1XTn+E16pD+ydoYRhCfCSri6QFlDDVPsfvtKao1LrPTiQ7GysQ+i/T2Px21BeMKt
+xkChdC52zlpEST0vVavKs4GVGX5YTibibA6mJdXSKpC6GBXRD0zFCy7ZjaiJ93e
3o7tSxu8uzisaCGwR9rJ7BP9jSK0BtkgEmB3xicQlXsu3m/hWQ2rX+zM1coPNaYv
hP8BzeI76svvLZP6OoIcuid2z3rzxIumKBMtpC8J+KhkeI7Kij7J9LHS+KwXTZT9
EEZPK7yO4VPKa+tK6efci0sSEqlosliFHeN1eNFfV/LZPjEH8bXkbYFtWFVoiC6R
C4Y8tiEnmx7th/Jt6F0Qgl6sqfAo7TtRcAE0TzvhkrSQGuHc8SMKtCo8wRwqsJr6
DkmO5O8O4YWbtyVe9qPPG9pgMAm/9fySYfBe9TPeYrmzW9eNfsP/YQXFovBZSu/5
t6SZRISQUhdycfio8tm/5bHoHPvjIodi0+skU2tGR8oIlwxoyaO2sEdf9wURWgdE
M+cdr+5+MoDeFMcs8eT/HePXFeqwoCEIoBB8MdsH953SL1M6+toFK08R3tFNDoou
ZGJUdapx+L9zeIXrKAJjrtIsja8PpnOBaB0WQAKnyopExrI48wqJq9VE+LGcCUhJ
gmFHv1yDnQnKyrC0G9unT1cbnuK/a3yQexeRyuV473EIX2I78nZbySUabCZyZ7zd
UvlFcuW5VVjJi67XbLWzsheC3E66d5AH/aW8K+V/p2HrSdesurj5M/i8KHbF9Cgs
SxShWn6OeaR9AO9dtzPy8C1EBZ/OG9IVYA6w86/Gj2MiRt3HfIzdWFzl5CEFBpmJ
ywTTMQgj6s0R/48KO6S5j7rFqRQaLvk5zp/QLyf+97uSJV+2z9bVW2+mZvVsN99z
jo734D1Lthrj4LH/HCftE5sL3J+TBVtofl0QiNG+9zl+Dl36KrHISLyMgNMmormF
ryzbNdjl7gSS8yGYVkxXS3BZfvxxc/7nzNCOmTlA/D4alrHljpseK3oeLMbS3FCp
ro5xcDbLIIt8Ajksvn0JJgxJFzAR4ekr7fsF3pJTLbPYdl1iGLam58XKXon3hQC0
5oiE7zWQqSypWcVLS+YOlb5aVLCwKbRIsxNpKnWki5ndX6q8B4zS5C9hPfGJU2wU
iRX8WPOP3QdWbxjSO/S9Z3uUzO8UywPbEWOnaty4HEQlYG09yq/r4QdjwFjGCMv7
bFBF6LuVcVl572x97saWj11aWV9uBq4LbqpGZlwwPJ2b6mdldY/Yh0UnLhgntFgW
n8kc7wI4MpMEjfGEmBa7Z4u9ikv9ncjNnBSUt5hIolmt4W/Lwa+O00w+sFLJiGn5
SZddyCEEAESqc/WTizphe55w99ceWXNlPthU+qPQYX5RjKyG38SDDxOZnNRTSyYE
sfxrhUETIhaS/XWgTpm3TWxnO65JXhrY6szFOpbPcBPUXUaWqAISrhKZDAY4B5rC
xffCh92y9DY4ZB+B1/Zc7P8xp8ZxA8TB7gAK+qVCfEFtH6B3+94eQVPYxKtRUKMw
4sktF1acADDFA1C/QuJTg3s8SnU/qFNCN0l6EL1sLeyC8vtEQxpKwgIR56YXo0+y
SCp6qldcMRgF+6Ayyre89UvvS7yprZDEoB6yzvMLQqZ9i1Fr43zOkiZwMsgy8/k8
VxvLIOmQ10aF4SoTV1uwLbJ7Ly499iMEb+kHfGaKs08E9vFbQJ8pIqfrkjKBiEx3
1M4Ju4TqNC9FjPqPLBNtj5lZdwmh2mqVH254Yp+hlXXooz8LE6ajVrbK+J7nG2mu
hkNTuYthCrdLkAjVoXqx7+4j5+hJLY9BfUOEIbQCGERkAF7QM3gSar4SGM4pq87Z
Ja66od+jNrn3IClw38JbYfmyJJC7w0nmtIOHPpGJ8wXjKqVRuYBjfTdrkPBT3drh
ogTQOBtWpR6jzTL6qJUznBkQGz4xLPlDOajCVRbKo9VPz+6g+xob0nPEo5uqJtSt
9KqzGS2x9ANwJQkUIwON1u6YI85ggVQbES7kjG25rsYZDxGIO8xF9LmZD5PlUjAb
/rY3Ks8sA//uEZB9wv8mE8ViV2KBTRDSz5i7/7Kd0d/1b8VJQs8aa2sUZPEq1Fu0
GesE14t+BALQgj6vK0Iuc16pOsdDZNNC9eGG221yI9x3GrdkhwKxw3tGJygg+XZZ
ZHhSfprhhpmYP4BTlpgsJHTE4GBoHi1d3Ltko6lRxS88/lEvAHCE1khImQjpR7+D
L2UR+ec8a2Y+sVD5JPLt9S+gqMEoRhHDlNdrUMnzN6qN2+2aXWEFCsm0utDA1loC
xb7/S/yvKLzm3v8fp4q2B2HIDUlGoUcN3+3qv/Yh4AHo/YMDEu74pC+scNsutLSf
3RVoOKZiiYs0KfQHqdv4PxIx87XVh0Y/1kvX+kmwvRKqEznjlThF/VvqS7/y5/Bt
aDK0BBhwak+AmPG0F8DAxwWP3W1TSfAJazzcx00YbzC26Vm8g/D7w5mqzqqeNfcM
2K7C6av7/xFu0ZdbVhL4hCIOXRIzDXEGAk5wpgxBLrZy2jJ7nuuRD5qmw7JaT1+D
l4haelsc8Ibc0aHSZZk1uRqklzb2q3rWz2eWuwJvkGAqcSni72FsjX61fsCDcJxP
FkvdWO4BlD9u/jUWqPeOJZYABWD8tBQCSjFUGW19nRqf4dAJSUy1ma/7ZBkq42g6
YtZLgJT0p0sDLq51MHdqaMf0AyEZaIRgY6i873tCciHhDWK6V+JnWx+Sf9Y0Bxo8
YkD4n3Txw2Nc3ltYLrXiLnvVT7eBYkO5T6vfm9qsvsNpUU5zgXasVD1ZEz1+1KdK
v4jdUydLk03yTW3btF839s9q5RoUn3UZEN+pxHAK06/H8CinVMIE1jZVcEpPL9wQ
eXBXzn/4hqhosYPaX60pL/7f6bLaFksb/W7uAveY0axaU7AJ+OO4pJycqp+uE+I4
1E4JAHx11I0GeD1x9X1gRz2I7H5Zji6+yb7wGC4zXchCRXz5at2EwadUW/Snwd6p
CKPNrXXfprlk85piGSXwpUFP00EGv1ENviziAzotei2UF8ILvLFMqYBt73lT2R50
UABgpnsUAJu1gupst2lR9yN3P5XDDKaxYfgr/u2Ixs0H0Q1SSZQHYgHOku9ay8BS
KiM+Bp/pOjfeaVZ3UvuZ/XarhiKIA+pJdKYizNdkrUTIPjHUFHjO+EEholdGE6TK
mFRF8bHtPbLJP+qah1uDCrqbHrLzf2D4LkWZYrpQBJ3MyuVMgERSWNnVlcPZKhb5
Ijw3cRJWzTVnIN5gwNJsWHRghdQN5nY3OuYcyOFuicpjh931YcbmDo4UY0RxrVY/
VDjyyt30QGhS8NuVTr5MzW6f5ztn3U8borbBusQeixNwbPWCMg7c7byTBMVWINdM
3fCHhwPdrP+BOlUpfh4ljI+VqP5Koh8fvz6jLa6jH4kBFG5oUL35YRMVpbetcTfj
hJSR63MYNfZZvcNcjITqLJQXGA4KH3BHDsqHfjUfFDGMIfDxNuSZFv6cqM+rN+K7
1TZSskuAXZ1yzAtdHKDkLeoUygOIovSK1+ufHWqk9wQBSDQxxCTHFSAgL3Wm2sZU
QV1tahkHrCwqbZBwqBO9+/KTfUfcpz3TTWimEqJacX8=
`protect END_PROTECTED
