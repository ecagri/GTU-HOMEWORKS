`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sxwkNiXZ2AERKy4s+VAYiW7KiZXKjIjoGSgp76fYorceCnv/maqL2cKyfgOmRVRO
gRUnz6bna/O5dVNZ0TI1brx+C2pGp42yRX+GnsBhTAyJySzil9joIhRvWRLJHWwu
vHUNa0xT8Lf9ViwNrxPRJ8+sYLhk97SkGqHxdIXQrbHMELYPd2Dli7g5nAF/IezS
YmxqQSxIkjaJnNKkd1PZwBr7qi/AWrBXwKa2o91wTcmQOo+q1HT5nOfVWfVXqEfZ
LRLQK4SrEDbttNxK00snfseQngqqEPrtu7YTG9lS+twcraicoCsE9Ny1UfTDcBKV
srANdZD1KQYxnQLu3eg8ByRLDybQhYEHPJo3K5A5nYE=
`protect END_PROTECTED
