`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l6X+1sh+H2OwLgYieOVBJ/bRIFZ8dGKFiqm5pmB0iUuZe0v9f1rVOimgSMD483KK
ugsckWPOb2ikmVnBQT9K5K+dWbMp0mt4oPbQMk2f7Auvd9g2pd1Dgjuazfh6DvB9
JPcgknTJTzfUZ3Y0aFUtnIadHv143PdNqm3MQec4ae/0YyxnQRDBCGQctBljlxKm
gmeo9aXdK4sAEEkiYMlhN1D3hcEQle3/fCMPoNdN8HkjlrdGiIgRSQ9c/ihfEmi6
imcVCHwQr+CPIfZXSEpcjSGw7AJoQXWd6KhaITFAKhgXdEcULZHvMQXzMpqynr63
F2gXSfTCYn1j43aQJn9odnaAbV8E9bJnDYmZaUWJULQESNfmxLUzCCYzcRb2Rth2
wWWJsRrDPVTk/jPJppAbWkMg26wIu9nZ+Ux3fmwOWEHN0rT0cNr6s2wJT0b+J9xv
J17nWGDB7LwhsGmnq2tXFPyjarmTNnIw3zntpwKh+IOhvln8wp6ODm/ee3Jh5P4q
/YFjSwXiMXT1Hg2zu/Qqb6E/ByTTQqTWVyt6kk22RYMvh34dbA/OvgIx3etZTA+M
m6rmbwXYpLTK0hURf3mQY+1p9EQ73b0V51mNIBUb3HRLEWR1ok9u3IQ+ZWRBEvaK
bnTCj7mvJ5n6TwMDED9IdfTKum92K1eKFAQ5v5vQ/v+iA+dDquyVPkoFLW+98uFO
pZMA/aB6k2OyBqk1rzLNXfM55QzcEkusRV6coWfvrlcKhynpbdjH2Et0uRsRiYp1
qGDrEQ7Xu/VeYujHi5tzoZDiiOYke8Akxx74/qVcznUd+MIq4XKQqQuMB4+qxY8H
r8ufF+9w5Bra1qdfkl/FSfZSE35enAamWVNQ0OlZ3cNrRxDQXxi4l1VYj9SKpBhu
1JyLforUOHMJUnbAoV7aE91mP36EZG+k/tjXXsiGWRJkDcGoeQERHG4GfmIR6p1t
QEyZsS16VMkfs6v5WHZzglxxaXql5WNM0UC6RCRNzSpwziX08fhUh2v0SpjLByoL
`protect END_PROTECTED
