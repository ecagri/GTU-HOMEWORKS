`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tBg9t1ggt893pU2acIEHz58J/E12WtjaFpyPl3bJ0xHXSyHJoa+X/khzW0WRiFRv
HBbHKuUut+glAK1VxPV4mJciTZ+XEHKjvEziXYCgZ0LlgoKgP4iAVjN0hsJ3pCrN
mZUdb7g8H+vFikAv/xEVR7vXm5YOV49esvmU33Im6RSBUAf1IH+FrFF6zkDXHEDk
Z32jLh0ne2aWBdWo6f2VdhNF68JB9xrlmbL4OkUaFwJP3wO521+DnHRKufLcdRjY
V5GHk2QnGh4LYArC6HH95LiEoIMYNgI9+7SnOTxPC0xL+ww7FWNjGEeAa5pIXtzc
rbOCDgOKN9G+BiEGxfEBxSqTj8OCclglJUlDytf4l/EYo3EQZgD5ZWv1U8ujSmFX
KBl+zg+k/DfIXYV963QSpBsx25j1JaRH8chTV7Wb/epbpWT7un8TZWCAcqdZoI5+
JnuoQJoO0e++2O71aVsgUnTRtHJuxafXyo/7cLm2qdZRYIgEVmjRWt7+Rp1/SaO/
ZBR0FSY5V9QsDmvYgkMEvtgxq7vv9RKikT7FRNgknamAnkXSK9HF5Uvc7zHzm0qt
O8ZCnW47S9nDZ0br0oZZyprH/1IZmEWVgRNlUkIv1NB4gJo6K02VnqcrwR6+uFoq
o5CHdT8fpxje1WXE6pQUfqdbXasLZYyAA0cm+LAJzVv0QH420AyaGrhFbFTpootR
Nt5A85hzkag3BKf33f3sw7AmR57aPhPxZwUNdbuzJy5pciBUodc9xWTKojKASe8/
nsE6VcvuKCwC86T/X/ihe5MTE3bw8xW2sBNCH9illwDdua2C4a5MG4o8741Rryfy
29fRFmpwTwnRAHOr4cfv0nK4aaM1JjByupjd52wOxevZkCAb5yFcwyO+68PRqyR9
k6jvt1BTrPuqJr2fNvLCqkasKrHYsMPi/P9k9tLwuBY=
`protect END_PROTECTED
