library verilog;
use verilog.vl_types.all;
entity mips is
    port(
        clock           : in     vl_logic;
        clock2          : in     vl_logic
    );
end mips;
