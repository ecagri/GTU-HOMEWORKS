`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WRLPBAhQJ5DIaLShkEJEHt/9Hi/mVV70ifqPA9Q8n7bdBhxUzkdK8Nfm2jJerW/k
daQ5iIojxjdWwP+vYfmHTp7NdtKMMUnWH298dJIPcqcWdSe4i1OYiKe15fEqqW9u
FfpZh2k1UKC8Xn/DgjeA4CD1x0B0zS7w+zvgrqSXgl/hV2YCEWYOMjrOF+vAWWeS
o40cZwOR+PK3DWb4z2OHHpq9/2hK8l573eb/Ap6HpDNBgzOz8t8Qn8X+YeLeFGqy
seUES0bympypxJN9a6zODgIoeOVpYo178/fGh7kE9Jj/u6mKpSf5nWHPwJsojuI1
eds2gCFsB4LTjNwAjIVbVWiyaWRQJLKTRuHEEeqNRYJHSf0Jeg44rA40ezckO4Ed
yJ220KLTuhfMNO9x//7IyyPfcDPUgw4G1exNgUSCoTKYOGD2XWKf1wpfjrjT7lTP
NnXWIYwwxCzE7+FvAL/4aQH+auarNvD9LeH4C8q6tvxRNMbtJRusEQ4w5RLcJsj3
5uuEyuI/T43pzGh7U9OsIEWZoWn9zpIVRCzcU+ajnuJc4B+eLMh6dOw5YLGhHIwE
XJoy4M/Qk+zosrJaXfZTjO+GJQGOBOEym5Wt2isZeHpWJK29fEPnLBRw3gMItr0q
0hbqReGNft0RZijQlSVGt858+uHbtRa2Gkq3uYJ6U/zNdzXT9CVoo6JDR0fLpHJ0
/wfpR67viHZMY7hhdZtgGFpPyhp/1jYfO1w14xwvbVek3qAnfNIPcPQR5Adv1rN/
iUOLVQYuaYDCeanUw8YnwB1pUCOysqJkKl/p7p6Rg1Dz5KC/FH2KFaKfgdnnTv5k
AuXnUOmMHGJQRFgC3fuydgVddG70rsY774oR0toCWGZKkboBnmEStwx6B2CvQcJq
Fm7era7zwiQ1XcWRUZCp/W9nYJKuHlOsJmyt5EBys7ml0Eh/LYVDNfKVtlphQ1MN
glQJzJqvnMNkUs9R3rSCOwekisL2KwtppE1zPpkElg5lg84TZ2GAvE6ERgVMlrM6
XBfLIRthOwLBD/cIF0lbxN64yuOLlE3FUWWbCvmEZDANsaXlWZOSuNfYyA3wtRrT
OCKOKjKNzqY14ffBGI0Io5drMoDKhMKjwWZGv9bO6Llhb5src6Q+GOxIBI654u15
F6kXfacxcu+C7DBQGxi233GXwGklNDLn+TTgcXtI2uz5RI/AeawC7lSiZCVAgRMM
bJjJ60dKi9vDuoQBhUk6NB5oRPkyTnfgLe264VlU8GV966DKUzbISMv8LL6GGzKn
hfQwUcHX+ISaFEAZz/kuU1NUc1Gk3a/k5yt3myz+uIABXbO6zDPvLiGzAgkMTW2R
08W0kL/LRAksjgh0qb0h7CF7CUNA/3kaIGbzfHmpG6Nyu/xiRxZLvTjzy20UX8kF
q5f6Z0Z05tgx0EwMLrJehg==
`protect END_PROTECTED
