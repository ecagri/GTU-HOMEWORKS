`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bik2HBiOfvbWlaDMOov/4yDhley2CRe/zXTeekoM6lroBjRQ1MIqhJPa4CEopeuo
udi4HpEw4rhP4sn8ip91S0kLmtqAY3sF6DxYmi+sb2BQ+dFTsmfiCKrXoQWTx/u6
QAmp/Eun0AatuXT6T6PhAdTDDVtb32qGY6HmFdrZXJSps5fVix2gsm8i6sj5z+47
LEPKYviUIJWKq6JwIvRzGLLfoRts1XsPJP2K6VdlxFUz8QjwAnF5IcWc+eqAla+y
F99bJO48V6uwTqUzKJQmPnATm+OPe1zlQRFBVbnn5xokQIzvxXn7p9ItUIUPb4AU
0viGXIHAxDZhzqIoPlDfUQzZbE5lw2x+N0VZ88Pcq6OIwnIZn21YkgMhl2S9dmIM
Qt5AOzNP6wk3srq5+0BnLV/rYMY+keylmEa2Ki9T45wcaHvtZusWGw4gx1HurY9r
bSaq3dJmMHn9YYguilnvr0HpZxjni+0hXpuoVw3LzYncs4X8H+f0BUMq5Q8eAD6v
ucrX25/5KHYG/BNZoVZClHL7hWy2nqJ/RsJRqlQYprd23SWFpTSMZjNdjDiovaTK
qbjasjSyBsHsUmaqhvDrN4g3sbkeB7LRgE4ZNUP4VF5i8gY/Zn6xZK2qOCq6izq+
TKxJSAfOf+BK0TmKQQsLgDJjE1S3pyhUnUNNryzP6zna5jeY8VcwRE7X2hnBbuiB
jBEoQ0Busyait41Ghh57NSsS6KiugU7HpHDeqcN0h1ayjg/kjUJAir3z0TdZ1pDI
PxZ5Y0LRdwkDa+z504AqBg==
`protect END_PROTECTED
