`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SAD7sTis73dIhBfx0K+y+lNEmeP54jWxoeNwaV+b3ITHamSdOjgVr7LtIhfCA8lD
bOaprhAlE61+xkFozWxtIxYA/qN9RmECvN4OQ+iVCK0lkDob7AtbCEe8mTRY81ck
dVhe2hDiLiWC+C1c+GrA9cKQS4TWZiSXMTNZZpAvO2jS1U6hJ27e5Fbr1nSn0rmY
rNwWSrNCraxCJz4CEvH6mvhMarMlRd8D5B3FdU1I0nWdlj1dSdp0omskMFlPvrZo
Oz9Rb9wPwACNH0Ck/4fsh5LyAQLI87dhvupPBfsGTlyPFSp3/pvstyWZL+dNly06
RSgISoXgE9nTYwprI7j7Ks10hIHoYGW1uVCbxs7uRKu7fKyr4HhUnc3z9Pe2pxVL
UJIEr8XCKzJWA2SmHlKl1A==
`protect END_PROTECTED
