`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zK0zvshg3n2kuFhdw7c5e/ty9G7bOH44Q+eDC+2wP0ePlt319EmXdNo7pSlfVGc0
fm0nKPfXwDN85mG5DhcrEpwDL4CRx/6MhbjTWvLWIfWAU7gZv8r5mIRVyZT/9URk
yDp63Jh6Ctmj+NTR6QFX+lKsJ533lkQEIjIK7vxPgP7WfQsW/SN+NxaI4AhnsQea
4Snu7GOe9cOwlkwTvGutawLkyN9wkONS7iZV3XbqDR7lQMpBs7iL0ogv2qjgM2Qi
S49SIDjbNyXyg7HG50eTVTSgxTU7CHCNZjxeh7IDMypxKueSt6l+YfyPlMpjpW/i
hxWoNLZJKFctn8qMEfmmEYXyUfl8A4OP/pwSJPI/gFGJdxpt7TcwoR5zR0s6/g2p
cwh/9DxpW+I3N4NKeg6L6+BZAig/MZu25ouh+OgVcon8hSHbQu80ORSo3eo+vkft
OIhHSClEB0SSQiChWCylgp/5h45nWs7v8RzneCP3fSmbXbeP0smr3Rx1uXAkVSwq
cSWiUSyvAompZC6rvcz9r3Hd0yE/HtZ53WHC7Q7xtCVwljsEry0AwvAoNddfiM10
kcQYZox3yi5GsRAdEwZ65Z5vRdZirNTujOmdh1LUqkW6q/A8it8FKpw3nmZstCKX
LzBoyDbXPOgwZ/8I1TCthUmk6ykqQhjyIzRVy4WPIY4s/C+9hlgEtAvp13Za7HqS
i2hBZ9SjZUmCQIFt6l7xPsBsm7xykJgRLzOAWBBZAFC5S8aEbfiJrVN35+IkqoYI
DYb30SZuuK/Y23x6IpR6qSeS+X/VmWJeH4Ana+pJPflybMVEToGD5TVYk8pKaQqI
do+TaD2WjGQgESwyAgo3o41yJgXY5UJVuM0Kg6RQgjxtWVn9VI85QgSIEj1eNuJm
M1qmfQ6AaTwD6bzghFwcnXQiEGs9Qglj7zNUpdF4jZA7jVO/HRrWlQVDtxtv27uB
vEe08iRzVGLQPqWe/Q8ft7QT6I1eUu/pchSQtr4F6nf2tQ6zSN9ROeB0M+vFYPaU
mkTh1BRUT1wjH205V9QNiz4B5EwbZHCrxSvoMYne5M2960oX4jFUZ7eoGKjKaAbI
AXK5AJRJQb3R+4kA35rCKvuR6j+s4s2RUFX61R+4eWNXCP0TzcPElFVK/nDj/KdD
xCpOMM9UPz3SNturQ8kQMSkLcOpicco8a1lk/ATS/hctouE52qpBe9pttGoGxHXk
NfcaYn1ZKPd7M3blkP9s6zb6//cLwVT4PAjRELJT6hMB3Rm0Asbmh8jVTSyA4ILz
t9vsjoHIosOUCH5Rp7PmcTtfJ5ITO8tCuDpK3UeqZfTo3LE7q4kF0PpEkpgQiZhz
YZ/vupM+bXdXsKphBIu52sbnykVNuHM7yAVql9Ps9WxHr7qme6kklvBntnVyK0Vu
RKQ/OpaoPhIiQOUcJRksmzXVgnYCOHpBl+0LmUstcO4Jeo5TjyaykM8vfTw732ww
74h+7x/Nc8LJ8/WDQiVexy4v2tdK++jA2nz2UZD+tt8n1mgdoK7rEpNwVYpe3kkw
NCKuIqrI2m+knCw0oyrWtlxEInBPq5C7m9221N32eVYoHGs/LekiJ5kEtKSRgdVr
`protect END_PROTECTED
