`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PXjXs2gjFi+ONG6htq9Yb+bdRCuXp8daBa9gB/0WtZ0i6I/nzrIdlKi30x2gn7p5
X+7HoJ0dXPQJBPeWvEcWfuVf4Jlk8yBGVFSlifc9LpbzhaiGak9nvhyDWTgAe2ue
zZhlgrkviB6xomP4u2qVc3PuCC6TStrxw2h8vHWf+IoXPg/f3tQZvYoPnMCWGxH7
1no14s3mx1XtshROgYYwKX8F07vhYXLPPPOcKZqY+RqaykUsa7/w+IrlpcB/cauB
knvPSgpJgXK4U0Iw4E+5VnzVf9OiXp+oxhKPOBDcaHRwlSVozEyC0gqgmQg32bQq
UNcEu8cLiew0r8SuxUSwqXVIflKyWn0GJ98K5gWQgQsbCiiw5vMb8//vujTj7VEO
jwhAkd6/6MQrQRm2/dkBr/yKXVH1bfQihuobL5n3tTNpCDEoIpW21ERGaMKiML+r
KJRukr283VRRLLXacK390tXUc02vxsMEeWNlr+5G1gXj8csjkEZlpHg9BIOfIRKq
inTP87f7kcIFx1HYCyDkVxuBTz/bwCxjpWHNDkc6AHptDneMRRIZqWVOEbDL/iOd
dSbxK58BsBiPGfOtOjMCkjNDj8YmNcnzm0LAoiWSZTZV0w2QxAo544ZGaU0eZs5E
BsA4OFQBLYlruZYyu7GaexvZo5y5uqbiD6m9u8YLUbFNcwFc7sot9Ale1Dz/SPFT
hYyXceWbMZaoAY91Db7ionBoO08hKuYub1moGjxeiPwKGOlPFap8LavwoEcFOvlA
MneV1n7XwblNdlnsNNrgOGGSXKr9M0CyMz/DyU6iX09QnGSHZWFLGLBT3vlciUyR
rOVj12ChJuwAzAjSrIlJilMbj2N2ClOCW/nDecSEiWWm4UmjxS+6tXzz/lcWBxdc
vqYArV891wSem0PQ3OfRPtbrIuUXiimRWGCe0r3Yh+4lT7tSqoI7yvbs1eMzwDSO
qo0Rwi9BwYTb+qR1yNRNMy5cxqLqGb+QX0L90ZCaQyZSXvqlGGIY/8g2HOJ03FhZ
BzNQqWXi9mbAlNLjaYBsksL97I8W4NmYi1XCgA65LzlF3ZFzeijYQhi1C5BG9g9Q
glUh9QID2/E/PnxuCEjdlQOrqx1NJtz/iJanomnhxwYMOCXY4nmT3SGYLgKrjtIo
ssrfjUE7KMW7yMA07gjEa78Qv3K1SI25j3ZkFsUwGSgJHsIrzp1L+1eXI3p1UvRW
mE86jHB3Am6i1WUOMHGFEavl7FGbQV4NWfR5ScDoobEeZJkDTA6pl42a1yjYCBeU
`protect END_PROTECTED
