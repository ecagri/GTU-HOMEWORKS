`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/zSx8qsB52ltY1R97hkQxDWwkEyvB9HpqQ+g8anEEfGSR7P2QIoZ4RFvW+OS+bvy
bnEZVBmzKYZzKw5kM6nfv4dIr84QNTTaAu4nmojEmreFat8XkmmYngAOdOfRKwJY
25jFQ/1jlwZPFKL7/+X8cGfs+R/1enm5JA09Vhg4VV4Gb+iXjcILXwi6K8F5Ng9Q
zaCwd8FLYjsq4qg2GNKfIlM/1U+SK2J/pGqZDJA0V0YNRDzo6H53Y7gXs0+c+yRP
bjVPVR6HYWD8LKqm0g/q12vrNEfkHLz38EMGWKd4uXkgRKIEn6GrkcaWf6HkRpuI
ixBklxC0s+Kr5Y2HQ1Z7us2ebiKm9YA2xPP+BQOmQzoBwE796/xhYSBDXG1A7XoX
wI+7JXQWyn2yD0LUdqvzZXWtLUMqIddOBntYz1PqFIZVHE0nLHmPy//fCClWh9Qs
tXCEsyZsCgbUKjgvthGcDwOTocUfs+M5qdHVO0fkRO2ugcQb5Is/tELeYPBFbaWS
OVccC6woGr2u/34i9VwuYy4Ea8+DLTCwaL1NOWTdHu7wty2jH6RH8PDexJmQF72V
Yey+N542ligMhB3QVMpSfhxQQ7li8fPDP++qjd9cox8j/7PJah4E+wB9VsTHMOlB
9WxOs1ZU0If8vuNkR+RnMai9at+z8skjS5jis8+cRV+A9Vc7QSQ0ySn6uDKW3rc7
dgJzlADROVPQddtgO2vul/yLbYqgo3uZJoVQriH+tIULQCJwnicKiYfCQj7506ig
TqEq3nBNTOsu0dw015rGI4vfpyoQMIswn7p7zFy9Aq2voScnqdGXGMQISZv/IbGR
m7FsC0AfHu3hNRaosbscEfLQo9mVBKurH0tDuM2ZwbbUH5TFsQgngyeLoMmNyQ3i
d4ZjiiagICeG/HYZV1X2gZZy6SH33FPhv8FQNpmglo2m1ZR4wE48dmktvIrE7z61
sUCfB3B7DF/RrRRHNklSHUz/yAUe+UiMua3oVKpCQFlt9bMVhHrOjXdeX+V2lpgu
43UCtVZ27J0Ki3PZAhviCiABKX3jYYy5352MBVMlYyfWMaedpeskc7g/f5sITwB+
5zoHsYvfx3OGZ6QUHUhw53gW9coVkcWlra4eaYD3MQnaZzGHU6LciWfVWNyQwR6e
H3IcaDlCJH5FDu8bgqPkpTlkxhHDhBnEauw6KQTvjP5Xw/28cm64vyRAiek22Pzl
/Zsi/qhgRJjkQHC8UlGYGxkiu7xvGFdHOU+/qOiD2B7MpjyUkslE1F1ph+KDJBCq
b8PEt6rwvDIaNSxmODgzJ3mZiRFAMBA0j/amVxE2vY3QM/tsaT993qDCaXzsTYGE
PdJNTj342DAEG766a47aWMzQsLEVSHka1HQ1eCv0RMeYwYIFKvesQAsF+y3NVuxs
8Q+NPyOZR71Hwr6OiTAIim+y/F3CxW2RwkGWEpYSexWIlYfJEmsZYAufCrRtaceV
zgqK82fVEr0DB+HgJMR6013Wpnx4NH09o73xEso+wVKJvuGt7nhPVfWIc6sb8fbc
s/9e6z7P3RjoAwV4jBpHMVAz37vdlRNwUGym/p3gy+X0Eb0ZokBuoRcgFciEgGX3
tH4ds88KDB9wAND0uHM9Uw+XqWU2W393F+vef008bLWZggsyraxFEx2xz6Z60H6n
6gkwQYCBNBxo7NrINukviBqMXdnA4Jebrp+lnUOpmUL0QE7fRC0ERNAWj8HOzDgY
FIxBS/z7HIm2ftA+muo/iaLkMGZBMAepTMK46UZ9K+ghv8ZqgdFHSdSwN6zgp3mn
bNs/DatDnycZS6af9IigHvG8XCOUGX0kdlXmZcMVqnzGNjtFLKgsy5c5C9wDMSRr
002/uDUDupKMR5KMPO/E5fLvy6jD6t5SxmFYlbyHxlAEw6bN1baqdOiRdw8xtroW
F6jEUiT4hsXVECiqDWFWNzzSr1UhabGaQHZOfpxqr27ICyTnrVFavcRWtHq9jTqe
p9xqrOCeehL8J8iG6PajvNwzoF6Rxrsz1BbZeeQx/fvxpIT/X9Zp+jFD0DQ+slaf
TNt/d287n/RYkC+2+ll5lO/dcbKL7WIMvZZ1gTqSdwXCIOsb8JEcIQjg0cYdx7IV
iZaF7EqMiObUn9vx9XVPEzsC2I2aBr2Yq3uHQztU56AEJs7KK/oVjMbgvuPX8wz/
ZF4c3m7eY0Bkn2n9c90N4UMxn4nB7OYjDD7FKHp1oL0v6ED0ytOOO2I1v3CWMSe1
m6Xb4axymdiSrenADfurSPDAcWtnAIKC8OrtIH8Umg6iRxKWjFu8Gd3pQ7XW0gi8
V0SuNe56tDDkuCaWmLVCqOSVzcG1zZBkXpmvXek/MBOfW8/rB5n50L0/NwyK7edp
5CeN4mjFGS19o5Xu2Cs68VtNwgetUVxIYn3Z592tU4+QRNXXsvdW3ynlFnFVo9dn
Z/mxWG+hfFRmJpOeOU9Jwf8KN7p89SvEwqoHkCnzSfxBQEks8Gydfw9NWTdGu4zc
OeAOJRB0Kbh4wuebN9/NWn5kmxFSTlAfIFyxcTkW5Y9nO2rBVjoXleuwqsOgMltw
mtK5vkEBISV1Tm6JNcj+WOy2v0+7XpRXatC83TZs1XEmJLwi/7agiE1TFJFO8OsG
rzRKzIe1P+5WL1wgJnYjdlfu0FBM9SIv0P+GkRsKwNBw+FAU7gDbF2aYDN/00jZL
/QX0+ak2bo/WsAkbTytGgONNp4q7Ce5hv/OC0wB3TRZT6WAwcR7y6+xrMbp1Grcw
zdj5uAQx8Acoto2DhQMHfuAXlIaTFX5V+0k9QVxv2yHUzT8XhHZixGVcUZxt8rHh
0bKCuVOjlrigLKYb9MjiTqUUTUJpkSpuyWho02YFXwOsmamBLSBZmyh6UlWvGxjM
IiOTJwGkgwRICxS5aRGLQ/Y0sQuR9COoe3wbWgBHvT5pIqbpDiQw/2zmoK4j04uu
Ki4jXpAaK375l+aefxT0s14rMqlTkedy6vBYxxuZ5pjmw4Kezl/Sz9T9ETClvAHZ
eM9JFUY1AotjWAepkuh8YzgvGch1S6i1NH2oYzQhJTTja347YlscR5DKMmD0TWUV
WuuuPo1ogtlc+A0gC0WU2T+le/vM/agZrWK7tzWiUVyl/w4He1LMzWEm9J0fWZv8
EJ+RGeystcnK/WrH3vqy7l9wc9anEwURBUxv7Z/ZbBu+F8iw/r0tbUe1RIss3TyP
NuR+0ZsUyaVtRcwIfIXDz6RdyqDuUbhj4HmwaO4/yFxgsQ1gUU9iFwLlwp8lvF1q
P6heRLP/+RrVbyZRTAXI9tjW8P8Jw25oMCfPWlb579VQaebOgNmffPB0RQtlFVp/
Dfkcjj3goEBeLxdNWQgUmh2P9mGNwzAILr2Nsfpp4TNAmiGT3/NxPdyhBJXB4NXB
D95WIFdSUnQySq41z0s7Lxdyur4Jzjwap4BNM+y0LGDKZXfeIku4GZDtPd+5/oGY
fgiokgoT06oYDJnzYVuFxkNbYDBJ1Y+TfyeEVSXj7mhA/b/0Venhm0b2w15kJfgP
VheBBectFvIxQabiKUe9ANles3C/SBb1x+k8fRE6GIR85voKxBWqIsP7Ag2mNcpW
ZzEAHdtVCDjwljEGYh2RTbMHk4gagPnyONf/JPf6mowabN0/A24Mxx183bHfLDj0
Fx+nQ3aTsk4zeWgi5XlmNnYkH35MhHEp7okzZkR2qcYc4Oc4jItx8rtJVXw7PfVZ
fhvJ4Et9mcALfwHKNR7vglpjvhNQyQ8GuAe9yt/TeWy8R108JRlxa0pNDDW/6jwX
q+59IWIHX6TBykTyIKkSWej4tF0+GJ4etd9Q4Kbi0QVSBnoGtB9z1eRslF9ZATV3
plrOHKIAKUlRgrgFt9FrhO4Cubqv8YfXVFlFce05bXz8dlz/zEDJVBHBz48XBxxh
bJP0EwY//Tq1W6qbQ5jXu2PfDotP1g8CSKoxxpNmjP9VDd43RYqd0pGup4VzjBFw
PK3k9J3XvqqmtDmLZxlXvg6/bsHYqQtRuB3lc91YXWSuCL0yU5vnniVSZZe1cSqq
Ybm2Tp7i6QYg8SRKO+U4tFTMbyPQBB60Pbjy4BnCXRML8Wqf3c3xT+oybdai2VZn
n6d94X4vsIUqGLOhFS7R6Igl8ndLZwx1+Zy5wxu3qhZ52EnenkdvthqWtulNUqdQ
57cQMVoKAbU+NNaer/1UtSYCz+96mbQYY2oimrrtz55/8sc5dhqbD5aCAYo+Y2ha
GZ39q+EJPkMgUG9D+EoO9CGscXGDCH7saCCyWJT+vBYxZSwmhjdzBMr+SaOa6NNk
WOh7jZWxi37jgW7+jBBEZqedccYuL/18VnIFb+IJAne+nsD2EwPYD4ST/OGP9gTl
3x8IMpE9ZeFy+p0lY6OVtWJuIFijZNUxTvFfKqanrpC+X+xedIyPU8ezVjGN2n/l
cg8ZkEs0m9JW2YhRwFkchl8HUxCnR/Zn7hhP839NQkJ02XL+8xlr8NMtSvJPWeWw
S032UMQ55nbRgl2uz5G026OQ2N8upmeXa3+XM4G3BCI1URdNAQStGOkY46bH18l2
r5F+6GbETUSVuNntwWgA8MP1gykJ06msffrz2nJ80Hlyw/iPGO5X8zcqrEXijDBo
M5NHXGUesZp/UVtw8JktuQhUcI3WRHZeD+A6Tw64cCcmnPcKMsEV2Tii16cs7L5X
unFoUmtlx22UAZnvZgyyVlggc4rzSn0lVUXokAzy9oRBqd18h0o7ZAkOlmjQEiAf
dMRm30zHJfJVHxdrktUPCGa1HlRhK77yC0T2r2BJLz1llCwFBOKBAVSMZaMMTabC
xt+L/9yekPcNzHrAgfWKkLx15Po69dWSkrTowLe9aKE7E5iZQhbl6DGkrcDoRFUr
uw0+PNdJ8LpvCj+p2LpHzoFehw+HvU1Bx1fcmtjUN0eoMSgA8vYpkG619tC+qfwU
rbe6OZHWqzJmryspC0xkitxteBnJnoOPpxbHdC0iJuZZaPpB8p7n3DkXPWucYJt5
7OuucZMztw9fiuEWpIP8mfBVtkCgPxNoHn1YzopV745S+rVuyt6TgpR0TTxsb1mn
nuGZuJYF66cVa9TIuEjmtXVYlwqU6njv3zawq5n69pwN7b9Us2LkY02N/hsbmneN
TQsPgTqaDBFqYioIUqOFx+UMAuEwjkwqE+wH2lyBR/zQKPnktYicuw+WNe894Qle
gUsOrvJtr/4mZQqmVVS/yhF/yNmgMxUlERSz3xF5kQQ5GuLtk9oqnextEQZk2vKp
/hhCs82lkfaEbHzyuGzNfJGDpqhBNY7gPDhQNu5eO62IMQvpWrx6B7L6cEb9YyjP
8OTujEzb4Z4e+6Nn/fiSLywi/2NA3rB2b4Y+DCxTfnW5eoA5q8ij1GHvPAwYeVVm
MdUXjxElg6Vd04xpJu1uaDvjl94h6mubFSRQm9jn/KFm3Vy0ThMdkUHZEO2y2kJn
vSQkMKq9Okd9+5tCFk6CR0Lj/qJukA0sslYmrQbHsIgWVrKMfgDbyY2K6DIZLuvT
HIdJO5WII4tTh/iygcvZ8Na7Kk2mKhN21ndDnKW0GNuRQu3AeAW7YC/UGo9cLfHB
kgsMwO5F16o4FtXO+1e89QUOcut6+bLHQHpfl+gHPUMCta3owcHfzTGgH93/E41X
AT1sbqHNA0QPWde5o9leWCB66PbCUlvXA4Ug8GwqT8BDqW2aRW1lxN47oxt8xtI7
QcUy69AMUiIMc3pIsgUKoph/uJqFybD03Pjxexub+/HPRby992UC9lolOLIHZLjT
ubB3zDuCilVhUzQQLA7PeDllkohKe+3rAOrcedKf4Iguhi2J/FiCWQX8RFw020Ov
dBbrjHuN9QqTxhmJrcOyRno0jcuRlgIvMhYQzoi+51WMGvgHwLXIKS+v4ep9gYoY
RAEeaOr/fPRkqN1Vcf47HnRMdS5rUWTNznTiUO87FkyOVc2dOj0C6EKc7ZXG0+Gz
W+WOYBzUNEuR8Fefe+RE6Wauc6I+7PIjAmfW9EhtYZKKQoL7kdh6ur5mmXDWZ0mi
t3pE40HWPHPzpYYmpiB/GR6HowWZL9xOFuxqqvFyKvqlJRs+s7as6IdP7EJ+R0uj
u/rbmytAfwnI65smnxmWv5wNFlneElwxiBpBHJDAeWaoHwcKkmXO2BuYATEyMFTO
84creY2zM5JxqrrdDJx77vIzrN1E1c/XygkI37h2ZHPmj6DswBRJto8u6GBNOq6s
186zMpps1wheCjBDN9jp2GbSOPHhTitCR+a5PEXZYye6VJpxH07usDlwH8LQ6uQq
GcWKv8Iy6fG7grpXhtJXohtDQ15qcy2d+ZaB2vcVTU4MALXNVFj5/FtyNd4PGCej
6b5LDvS7K+GSVFOxaHQApk3fwMstsf9lr/EjsRlnD3Kea0297X3RB50+s6NzEeNN
O23zjrR7gwybgKKoPmwznOPYEkK6wzxZk94Et1PuVda4zNAj/XRZWzBwOmBQYpUE
YUiDsCm1N1FkfVOOEqJ2tPnx4sSYHW4a5RNi5IFSSaVFfwefbYfdBtIeHawANxZn
TrU4Q/llnUjSYgLhr+m+S/b6KREPIsGptBy1yWZyopaRvUcOtvjUROBVjNKmefNU
L9nWl6HzKiSvW3HKK+TPXxJ71+pq5nNa6Ta5Hjm1EQMlHdl6yVLiCcGc3uCdwWtm
eS4YWwpxggLL/IjePEaT6lzII+6zL+8UdMNd12v1X5q6gN6JAll31oRLTrsSRy50
pdRfyQkyD8Wa21Jw3ec4p05oiCYfCy8DHG58ZM+9vo5/LybVYfpdQ6fOO+uftrCi
hluKoK1EOFxR4R2ptGvy+P1KoMEB59KugkkOIxibGvSvkhX8QO/EfEiZ768eDkL0
5XUP74cdsBIAtYZj0zcj4l4zptqvQstpger1wnK8Uc0zyI7+pTSp3k+T4lYNJoBR
Pwn6oCugANmeYiAG8wBf7wWBbK1gzHNo0eS7g2g4kvmUMehheEQe+73xFFIgVYFe
rUyFZPeN6RpkRn+PzYzcuQLto7QX682TMCBAJCP5HKGdjM0tvHxxd2ZxqMkOgAiH
bx9/ML9MEOvd5XWFFCSDm2Z2g75fCsyB55o2I+3sP5EHdLUZ4lvZ+zp0KKg3U2a+
4wokI4MhbO05aOD75taEfR1ggbkEwF/JWqRY4fcumWmW/VnUXQ+poOZQv3x60RmQ
yA5QRiytxUMkSMllUJbo0aj9ib6wt4s2W+YTRYrLIEBwlACCqmMSBv+eUp7PwDhC
Qh1Ee9qP1Ir9SrNX1/vkeG/tqooZr0AZjsqMkLXWwReEDMb5ZKcBdJmK/RLd7r1F
pKvn/1oMRDZAfA/a6xzFalT+YoYGSL+gyFghuBmsTm7jSZmTeSxRWSZzxLdy61oG
RGcRN2sxHYzXWPILV4yicYBTL2VdlkRz/pNs30VbH5RcTzLJdRr3g8L5nvkRO03E
s67pWZ2B8RppW5uoVvXS7LLWgKErTd4R6u1j60KNwvnMZi+HyMYF5zOfX/1bQIQw
3umMYCmP2wfAZMKJZ6ypwTcGORZha9PiTbLoL/rkq/RnzLNnrD2s+ChfzxiLWvoM
QF+fP7CLlFsGBfdBp7h0v1ox4dQQRl0hUiBOmGfUcer7fp64FdALwzd5mun9rjMs
hry6v3tAnnkfm/TbaPG2n6E2D7oc528f+J8ItGJI5gNB1UipnrJ0s6oB1ggc+41d
0TKbty251rnAZAgpPQcb0Leag/lMKU72b2vaTHl8PulmxKkSwMSjInNYebThabsp
NBAyI3vRGN9u3lztHl79n+c23d+Vqb7SKwFXduCnQoFHzIBWKPm+lPaEVywFfVnV
TyDR5isLFPvTZJk+diWyjAJB2bi1QULsnuiFoKOlnVVFEKGLMaNcUZpJXVXFUMr8
MTYIivY+v2lpz/YBgUgwQVFbrfqD1UVripSlyWYbnxZi4lRlXutnp7E8iIcAFEmJ
JBN+2JcISs6SDzYtKKrT/pwe0tgg5fbEybRfXeEyX53N3ZGjBMYSlIwJBqEzDr5+
z+8DRl9Nuk3mb4glxwbrH6Eb1YugCKxWvNo/+HG8YH4VKgT4qfwoKeBVJCtKwJhh
IKS6ye7oLTfLj/fokQz9rFVXbD3UB1Ue1O8yJStTFFwG/b3l+H8hkEu1bnHJvSvq
I32R3615AXVMS2qzzWH6TMQ0zVd0GMaND1TaTmasPqADXLBHUkRS1aZt8dv8tyuC
MIlFKBNFRr5N5dnLOKH8EbLvCYGPLqvWVPX7PfwbKhZq15p9WrUJ5Zu2f+oil568
MoM9O78ROigo7zvHYAO56G06TLxlQI/hAALJ6KltZiKwv5+qNDhUPINltOttKjgP
jlJgxO43A/kCl0BBRm/r6fDkUHzLWbNaxjmRobWO0stnBfVRV/LArfVaJeJ1TuMQ
NyNrJyahHiwqhQ+BwqLETL+QSd1HIbPxawbpFIfAETIX4AfrBrM2Eitnry0Kn9Zj
8B1gbnpRskEaFFBboqNO0QgscFh+r2VOcZS2w930AKZb9MDsjUZPTyAXS3UVTpLP
tIDx+spdoHNT1rTq9WfPBKpIb1cii3hIvlMvbKJMxakeuO9NHcGEwKFM3OKh3jEn
+pd8YSPYkpJgc52vQQQmPV4K272e+Kn+P+BF99ZDW4Fn+C5z1qyF52orsycIp/jF
uf0S9AcoKZobNvn0S1x96X87qkqzowdlO9znfqmCvevcuhXgluarLJamehipfT7A
O/iXD6EaT/xGJkWbpnFAxGgOmJdosshyyuXiZlVaTc0dVWQ6xiKwdM4Pe5VCBPet
unhzYRO9VeDURXqVFtdelEM89r4ECvgEUMcU/xOvirwqjqRjSp8YwVhEAKeLHsUF
RV6QQgryKxSNF9p4ORRTKCe6HOfKljQ3Z88f8/Nw6Fn+kN3t1Yx8damOHpoGOnMa
9fozyZSHSJVsu+/5MtySokrLJ00p/NAkFPAgSRq+YQYuRNaiVaRJ2cuEtM+rof30
2iO4pU1nE4KJG/daTJli7xPSeRN7Tan5gMw4MBEzWftHzNoAGCoyG0rjm814on4B
+1gB/mL8hDM6+ouShfekLfy0A4LD+tf9HV6ebZLXpUWTIfaaYuhKON0EXQgPYNhh
WOLRLCsD9SAMp6IDWHZ1mgbWjYil/6SJ2r2MILvjXbU09+l+6FW9Yvs5aCYU3s1P
km9ABSzcfvlB8kUFzZZTOL6K6i13ovH7mDcWUHztSyohez7XfO483+Cu03iT81RV
S/J9Q2V47dWGMH7AalklbvcLPlvRuGDaQdqaHYAfEH8VTBRFqq0ep35hCCL5B2xO
SBRu2Z2fuZ6Vh/se4nutqj1GDTOQ1ogYMQCsIYEeGT7g4JHzzRCD+5jAuJZkTfgG
ATcJ0bG2zEge+rMHPoGHC36cQ+D7KU6A42Ew5udu0LaQidH9zznqNVkPzYyHKKIK
GcN6d5riM/TQ3nS511u1CV1jOMU02doVYsKYgNRgZwSycaI3E8wvjEIUOAHnuUR0
5I93z/iqJErUgcoKita4OYnQ05hYanWMEZMAkxpd+TA6cJwGKna+0ST5ZApgHct3
lHgUEyQT/m9xvIV/qw2xA6za8/xU3QIOz+3vNkDnyLldCglVxW/cV79ihEkv6rNC
gD5Gvfe4w0sNB+y3M3DLmVhumHiL7/LrqbCl8+UcpfvGmQtrlmTOdaIufUlaMhjG
/KmD8ZcDmVQmlgAqeut7I7YrGvFHRtevQ8t+kwlYV0vniOcXavmGBGw1K7KD2an5
zNDfA6m0wTdAqCUPjATNQhaR1hhvf95eUNLgVKY+aHm22p10ik4OJF6m3BR+GAOM
3iBXCHJGp2flGmXzC0kXj6wr6zoykh3ib0wJUXQTx2LOOjoY12Hd1jkwWNLdiglW
r5b3mVf43mhTHNcdQNrxZeyolk48iFk/mUPO2KJKtPxa+WNK+ne7a0YvEZCjSodP
d/MzVNivlzIFr53f4IEmopN0AlaqZNmOZ1PWAmUmIa7QfNFVVFJx1HZ7T15MT4dT
1Awz0w+6t9MxnsulZD/L03sMJVnXjLorhYC1kgOEgIJbWe65/G5tKdafa0LFW1Wq
OkoIrs7tUkhfulNzyKrVH6f3A30uB7AGpXneLT/jHsqptg4qH7OXQZxvWMzPxEDA
0MTQyZxFsDkojjYD2LpF/Mtkl4OrfUapB86MHWFCN5rlIazbEWZMSj6kmrvYC3sk
NlRfEWayV8hFwIynOzQCkM7egWr05De7DK3JJK11Ufu34ZY3SRRKWeI+ywKfvEJa
1mmPRKGaN60cfc+i5bQ9tfPpst+LkkWHkNqKKH29xvaN9AyEnVuCBODrtOff5wMc
chXekN5nZY8UWo2gOChm4S8HrxknWpSIYdQ6wHaCabjA7L1+aWoNF6bfLudJnavO
E0dg02T4WOh2po9GIjCX9V4Wdt7lF2KpTWo88Migq48Hpa5FUFI0dXCZeJXY0Kx+
7+9KEEBIZdOdHzI3lpHdAJHoy5z/J6y0JLK1m0IxewBgalXKs+3Kesz9Lt6S3Ysw
g5raFAaq2I8B5hgVGKzHiTyEmkJ2DChymaKIGA8EE7xDcNPIALTBAB4xsBQH3RFA
vcl3HrYJFM8Nbbu/Ye1P0KdwD22pYbbxKPXSP6o/28JdAMG5Tto+kktwfplPzvkW
zi4LLbue51WbXQ1t/U7c9e5OXsqk6FlvxAuBisUpNQTDupVxSE+XcZmOBNhF9w+X
q72NVazoBsh2FX5dtYq8MJplkDO/MDpkWm5/WvqviMMcIZSTctMKi+RZScQef4HW
DKS+1VafJa53fnZ6+cjoYFMNwmIoBfwwrHhalv7JvjaHNaFhbxG4ey8VbJxuUy0V
CmlG4tmvN6hUFz33+E+rFGPwY+EXIyyXtVt/JPn1miRdzP9yGBrVOV8S4XrFGUWx
IdpIQZez7zV2XrlbL3VpNA0MEqs+qhLeAc68Tr/SiNp1sPNWrktgDciFwecICKXp
QhOeyhwRsZgh1sYtnzNWSRjktAHwmjwsLCVLfossRcN8gUeEnc+h6uHZo8IevqG2
9tEjPQeWSLLSyUshFPsgKhhHHnpkgzx58m1ai9x4NyR1hb/Yipuyb5WM/YbEi8AC
+8txwTOVmoYBwlqc/ag4XhoIoF1sia5qPgzr3+CUkuJjyVQY+AGP75VmbLH+Mtr7
oQSzx65KfqdNOm3AwnGLGQ5vUMgVnK/3vIlxm1TYn+6DFGk3+iXO5WunHX7sRSJf
YX1/31HasNkXlaAjRSVIsxLbY6Sk28SeSbtqWgLiyIAkU0yU8vK8i3PY3eddKaAh
dO6ZyTS2y3FsqS2eaLVHvDjcC6/3gES5/ut7Nu3fpo5iklQ/5HlnbTsiOmhkWWkM
Dv1W/C9PAmKvM/EWghRQ90m/mksVj3+0VULthKA0Ar6L57jQTlmwMAA0AHZVslUy
ok76OXV0PtAxhEQnWVuXLgUJcQ6Z8Rvvt4uKmAe+zlQoAnNfg0GYS0YhViBpLxoS
pBbx3K3xDT7A95GaLY2qK1srBcic9GILBdH2/XS5NJTmm0iRDXPXpr3jgdtATYF/
3Wn1Fk3HH8c/dCTepWbQQqb4F1sjbftTzKrDcjtJvMSoWIx0atrPmtRmMJk6k+d4
tC6oIAXlkd6aKYzQTfkad6RrHkNsNA4b+66mghFm6QfYh0wQ5cGer3hR3wMnenOE
50zsvRvN0773+o1vdzQK/yS4j7cZZqWuovdGS0O/311RQq+L8zX/dwu6KPxXkYF8
3ISvhQaT+IMVJQ7GiOwpvEgqU1crKs3jVdtDgF6WKm5QhhtkYNg5dC6qExIkYnfR
HF8+w85n88Q9rEfIRqseBwBY7340TRy43di9YOwjoIqPVttRcM88ov91bBYAqdsn
WVP2Q9aXSGa0YVflz0Jkm36TQJ+/Cg83OCHMTX0oXG7XTSVThjPYVTtAW0PhBrhI
3+67DqdcC49ZDnsa4bE0JmZne0akO+GQ9S0g+V0GT/Y5V/JYUJ+rA6r0FL4dJQCk
kzwx+j8an9ZD2HQfhTJgyxioLHvDIOWuSsFGXbK1KFGI5UKNczJUxtHgw5ey1VYL
nB71SEMEyujiqna0LnTIqB2gCHoJuTfUXDBstgmMrdpTQhF5GGC8jLB3gPgA4Qaf
sYzI8RkDMTMD2hQTHp0IqaoZyKBM5aPkWnUD6VKHRtor8A6MWuI/EHyCTdZEQvJ8
wKJUViuixyJ+BLt/ehVmAkFFODS2ZzmIkxpsPKSW4kv3JsHtLZtvztg2dcH661DU
1YH4+IzYO0b4DUjokVLKou1SxFt/e+Y3ZQHxgXf0e+lV2IIVH+1bkiEbag9OfI1c
OxFguGWjgIulc+ISOVEPOJOFliyrZTl9kqQxt5eMHUh4LunhXmo/xT3zgPGLC8Oh
5FEQ4PtFgd6vqbu/V0zDrUGTOupD7l97j5T5s6z2J0ks5ABBPH2PS/S4ykj7bFhf
l6qsVD2uxqBr0DYUOCxIf8CrFXfg5U5wH1GdVNW+6H8NAlwcz/oS88jQELAGKbVE
wHT9CyCYI4OBdmj03nYoBjzxMCNkzBnqfrooS+ryFZvOEA78SvmlnT7sp9HuFEiH
d2ERRB39DWWzwlCyoCjyVRx7E7+/r7Vm9u8ob0ReWye9UhbDNAH017AbXVzNow+H
cMBLKHy2usTCoxkMb7PMS6xc8qkr0hMJJBB67VISI9clFA6RS5jjJ2RlXaTEPEH3
K1fhcbImD2WQ6YfquxDf2be1blsAIhotf+Tp4abMew771VXn02XI7fVUIa1vK/cs
gWOShdUqL9tcwx/Skz+e+svudSX2gm0RM5AN8z/sbb4+CBvpTr2yaNlqgTA7zj8F
2iR4X862ybM0gnpNEJV6erY57o2Enmrg6byqG4t7YXDIZ+4A+vjzmZIGFy8Sz6t/
cQuCRQkIiJiXXKk3AIbtKxNDmHnV4PscORN13Gidv5PQ+WOtSd2unmC2gvTAE74d
L3SfAR7+OCNkt8dZT1scXHwvMqTxgXT0/xTCQyBp74OgugG40x4CyIy7Z9efqrQv
HmikQiKuMUcKQ3KUCF5XkJ3n9gxfW0d82X37oGHqkqo1lyGU14X0LPlXo6v4KLn4
C05+yd4qXBkGVUqOtFg1eiWSMhQaIgrqRBhhIWAuoGf5hP5t+Zs7q2mzXIJvfiKE
Dq9cZBo3+JPfbZHHYZ13Jfrd4eQY21eT5i6hE90mIIH4roWT9D0tvWQJqIot/OGy
4vs+OppCz03ZL1H5iRsY2+3RqngZkemgt5xLA1jpcpnub4hU9yrPAmfA0HTf7z1o
jlDyhdC7YRGjw0AGPtTRpqn61qsI96MdfA8tFzRgXuQTNrmjgjttY/64a7L+CyqM
eFbOW2Ayxmz/vTKtYMaduRQw0aECkvKpusz98TspavgyNB4sMLI5ULCrYeUBn/GU
3LL4uM0swXFkSxBKWRsJwGSb4EW0CTINR77jdUmyPDOvjN2Yhqr+VscUo3UJTm79
ZPsHsC8Y5/8yexcg1rPLGlT8YtnjbokQrYCSc8rd6W51Egw802IjtkZQQFQcira9
KkxWJ0TsgDOjvUVe2Segpy2FcM5PxFhhAShjT0AIfE/dEW9l7gpSUO41DUZboiwi
/MIfdzgb2/LxNfKLqEWQgVs9zpxE3crxEww6eun2L60tR/JQ4YCBQ3fHFQ/FuPqf
jfP7aB7YFq7TM+3+o2CdAUabL3GRL9s2N0eCZhNhDW/UCBIfLGR7jeW0SPeRpg/s
mvppdBtmkeTJng9ANcyqr985mVEtrQPwg01HXN3DW+Be/Le7dsR/8RhIBUpQXOti
soQ1/319JM9/6usA2l/a+bnhwf+J788E5I10foQ84FPVtEvdAzO5M48GlcbnSBiG
x4cjoQoip83Dy3wS/CJVh2OpbEJMLVRNRvcTotgaDU16JTbPiDSPLg96X2egoLEH
Eln1MfkU4YtggmpbXIJ8D+fs+Cu43+7Wb84QR1MEnjhDWJbU5bdoY9AUcLtkw3X4
Abb+Rs4RnPW57oM5KzI7YUi632VjDumXI+lgZ4ptXsKRSzJoWSgYukDsmcUr6scr
wBOt3MnE+DhmFZ3c79GZR/it05tdPhtmn8Wmf6FX1wsMTUdUNtvADMFY7JGMafmK
1yAppm5dkmgc6IHgD1ocXtUHlWXm1d5qBtWShnEBPIPnEqtlX0YxNlB2s/M32/JG
NhfWGABZVHT4w5fqA05ITmuiICGQg5S1fHLif1OUO/o7m7Ocw8ovPPW+x6XSRWnK
E4OiIEWJPbdYZrF9c/KHJFr6639z4WUSNaSYT+bosf0nCu5A5V0bhGy11Nn1WwqK
IbA3eVotTjQCcQQyewFXyD3c0rRNy1Scr/0nVpl8u4QQJogBFaGITq+JdCIMWmwj
AtdTtsEKpaiFYA4HEQ92LNs7dKkdBUHIBc7k3KFM4U0Ur9hUokvCqTb6CqJowl+d
uUjFOd5GZrW6EaneRmgdwTCz6Lt289ZktySjb+mfI8xeKmlOGCQDN2bKSx2h2Pwa
YrPSOtT6nB/1fznuZzF7QsOu7HgpngQ3Al9BosJfxFG0EyB1dVb0lzOzuVjPQOKn
C5VxcuNiC4OdPKI5r9LTUe/rV60F8jqiYzwPL5DGQrOetXwjE1Ho0SJCt7ICdueQ
CVGKTN62XY8rxR6vxAo3k+F9re6/5BJ68cPg9hujBv92d8uaUSp9d6no/DUxd1VI
eQaaJv9OlyOvjzhxdrrvN/RGc8mkekbvdCV94SnvM6GkqLeTtnj+BF/C8u81Z7Ew
TobwX0A1OI3wGHb9m1mRfl5dztaEr0SeRdmMJ9m6KVXKRZwBIjJJxAp42bhdiZrf
aTnEgH7iABrwyzMtJ8LT7HNEg6zH9WaGvAXnnBRR5UpjC2qmCj8M8CztcaaqryGf
4PO8DNDgIvMOgpF/Jg6M9CcWc43H1uoOAN1ShPFWqZAey01p8yJBI7W9EarBwf+1
ipzcaSJobl0W6otMTltTUVz9zcGvrgWB5qad4+4SlPwXxvQXTTbrAPuaNnebQGa5
OECmTtYTG2PNx++8YR297O8sk0hADmusRKA0fHjttmX4WocWFube1GekuuKStm2b
7Lw8qCmH/UGEVP37QaZTPararxU/D5/CqCmUKg2P402Ul0ZMRNfPOEcyPIMj6+VA
cLuyYLOw2rfwA0b+7VHVxQDE7jSNwsbxb9LAVo9CBuDoDAIawhUOm8jflTy/8Hu2
sun3cEpURhqgQHcHqpGDhoDPWNuy9hEHUh27nO1f0dca+h7THeSDu5pZoWmEuzg+
U8s9KwPPOQtNKMK7uSsLk/Q6vXih/UmIu2q+gCUONLg+GGi8mirasYCyJKiX+TS5
wkR41kf2byBqDPSypq+wzOqVPi38ljAuKXtiAk0rtzyzZrLKtUOk7prOIH5PZQE6
6MlJB4SCXuwMxW/Eyu1zvI+jLP37cMIO5eQJ+sA3Gf9yjw6XxDQf4r6YpNEojmLh
X1gQ8zvfvmGOw/B+I5aYeRFPbeGnEmqd9XB9NfZVH/ADHNHQV1rzZIHbOFIKi1X1
5UpAYUaIAEJUhxlBYNsaiaJwbQ6+mcbv8cJRzEXaAwoTvJVd3t8O/cB0zQ+RtSkS
Ha9wu4qFbLJAcaeC0L+24pQoz/nLUTD7NBbps35jJYl4/YEOt9SgZcBtP2TpwJly
aAQhs9gIulAKXw+aYV7rO++Zs93reiHLHQ4btF5OQs5yX4vvowhRWfFEM3ZWvG0j
4GPbv4xvnRhIlWLK133E45sfFs1KnDB6O1iXNVOIemq/7eG0opjfbGw0c9+xnUai
DbvqGdTokvCyvex8a5cnv5dIFLA++o5wkrvOBuHbvk94C9uEVYcaIubeO8jOWcYS
ziNVvg92kC8BgnH+L32SjJgOmBOiGDLqWrM+Sszx+Zh6Ao6J1arD4N+omuXKmbak
Z4l4ds8DRHCSpu6ZaECa+GeAu7aYQq6KuYLMsOSrZQdJczZr5i4rE9h1uJE/VO0J
qljV8dMgyBxOgduLUxpxjhHjJAIuHjVLXVRWYkozKLoiz69DCY5yLOS4hPpoP3LI
h8S0BuR+0NyBCVr8G0siYZV01QFgkApeRb8L6gbgkXJhw4FRlG66upm2TqG2Mk1r
kaFrAJl4RWOk/aBJD9CsKkxnjh74+R2i0FD/sub/r6j433fWK5f5HRWJhkClBQFA
PtYEe+fD2aSwbI9NYYqZOvAH+sE9MsRCFlP3Ye8+cXgwPh3j4ZjsZZZFLYNurnP2
BbksvmsxnIZQtcgOqxSfaqQHWEbLqChOkQZGXsETSX0RSggc+0eML2ZTQWO+kIun
+WoLW7CriHKepmSNStb8vdd4VzEyq3L/a/P4obpiPIz5xo7ojMLNvlRfVni2A6Wd
JXgPqb6/d9SmuXXQfKU8PzdnT02zY+kQHtwt4OlUADOyr6ydSH/0ZHI1iOWFfdC5
v7DHwoVT6pRZue8DygyxZEdUBvL6Ly2L41gVr0O+SeZMGJJy2LF/3sd3CKsvtU1c
HQXqgsAbroM/CRUjqUrAoldukVOPW207lo1LzTn2S5R5/VFCXPTBjYPYK1dS+AiQ
TXqYHRaDrLgCV8ON01GK52mmBPkObeOdZKzkHDi8LaeZkUUBb8us7uaqZJj32ir3
ReqQZ3t5A9B1qw/oYkjtrQuXeeWClzf/uNs08P48kaA3P6ilOtWEqW5inERo1347
XlL0At6x4FePMiI/dKhR/QcSTsMSADM9RtxDABNwH3e9RBaYF2eZs4A8DtZQ0jmX
1+RvWpFWfcaFZE6LWbaxQTK1BIlJpr14zSQwLjdkhp3eGmBH5Qekymh5vNxMNToh
KQplRXQv6n3L/O2hDJG3a2rS3MlWkNyX1Aas/dEsfZSvo3Cc1CQD69e8Jr02bdP+
38k+Oa9Hb9AMdj1hZezdcp7fWiu9QsPjpZhEv8YnC8HwMgOCee3rpFp0E5Yk1apo
sYZ/nHNNnrN3fKIiGN3q+N8/kVgYGd1Wu7lXvnN/xYEwhrM6q0R/84MMq+3QqOz4
bO51dhC7dp+tedeBr4MX8zYlI89Adexhbxwihiqxx9yYAJBigkrpB9v2yOTjprGc
F/pTR1K2eOa4IDfQRATRGABdCcoJczUABoth5V+AdgDytZiEd6Hz+ma0eDdFOYXT
tXXXT8Fx+3mcFbjfitQFDAri5TSKlXOklzD2Djr45QJ0z8VpXAM9epNTJ9eRf3Pa
7juLNWvUBgDXfKdG66DVQafpEaTfJK6/Px+4ENuXyNkPWUtiYUJkwJMnTObBgnRT
EOaPI5XDw0R6/HxONLR1ki0Uf/KIyOurPi+6Pm0IinpeFXklZdtG6e6kTOim4Yfe
sQVHsXoRH6gm+QqoUhdsV1sL1DXrBQYpS0iOqNB/NHZ9g9o7sbdfOdy+xvu7TJjk
AwHD2aexgVhahpTYZZhR7RIMhKxW94v0oTsWTLp01RP2dNRfvf90XUAFQSfMKWBQ
7h1Uv1zO87OETuyamTQgqNPUGyUPFcE3Ih37JRRphrFsAd6yYODdc1IkTvKsZlSd
uhIDj/XYPKO8eDgpj6UxUIVKcaRIsIUGz+ZEd6Cg8UVyuJd/04mL5zdxaCDklyKL
rLwinbPdH5qVsmWeVA8F4sfnM1dA3gNhw0eOb41WCGWP4zATQgNmDATUg4Oq0N5R
8LDyyq4PDUOibb4IS7AZ7L4IvV3UBVk9ALqbrMc+mWXwJhGAbhELQnuUQeVuiDiz
Z3VRS8BA5H7KQDbIeoBnf3+ZvdaMCpTvtmzfuYy1bMTs+Uut+ZZ/XnzwEvPBebjF
57+F+8v32IYt925IUIktwPi7CAvNszhWsiKlaSNsWj2ARiM8h6VUTRbL6zPexIJ2
drhbWHzRFwfH2lm2KWDdgAHEby6Dj41mlXA+9zmafAlGOps3ws8Ydj0hbD95lKS8
y/37hBd2DmLIXKbtbeZUllPpx2eS1UZz3KIY3PC3qAbyML0G6w9v10Wjsy2ahlPV
QqpxWMMxA+sXljKU+SO/3SVWAX3NsGPtzWs1fUeiOAdYkajBYsG8RMKlPOFaKZkF
reWh1VQDy2Ji3/o7IgayRBdEgrZlLOJx4deln++4CYsKAkTwCpyyo221HjLgsb1n
l7ZwkOsH1joXNyEVG0DPMdR/WvsW0URJGpgSp51aUX/scGMvBPaZNxTiV2I/HgfB
Yaa0wmv0ip6e4aKSpWhYx33PpCBFl29rtTKu9P4o9lxlECBcVyQbooD7wFn3F0eQ
dt1Kpsqx0tAcbCGHnv0Gjj8p00lcuisf0Gm2jUnCtuC13S08p4riiwRJ+NRoa4np
vt4q6cfNyLJXMOz+7f/Jd4tyk5jSdmu3lzrT0xa+fDN12kbSnQln1IpxjPTbjN3U
JpevyzPPGs98oOfRpwSlQxvkINk2SdqUpdgoQ/KjYZ0h3joS6l/i8bSCmdM/sUZN
kYpkkLibGdxdRg2Ng7XfSymvg77DgGig555nI4xKYC3+3WSA7yEI5SnIKGDklskI
UJZOyuMl5oG+PVd/SvkL2vETRkoAOLXROohv3x8CjshGPR+Vhzo7VanUaGXBg+RX
f1dhqdvobrJzzjHvOgqVcBCwOQI21fJR6AjGePOQqVB2Jtmqyw9n9ZxDORVny3P2
H06RuENCZ0fdnzJd0gP8cpoqqoKbHBm47iAYRN0MyR2/VpHLZhVOo7Dpv8MXXHma
D/QOULR6dyH+c60MFX0qE8sJekqCee/f8CKJfiTfL0awCVjSOUx6ik/ZUSAkbLzb
PrOWD0LUu7th3/eTUsiOnesK3BIBgPtnpwD7bFY8UeQPLo1/jqDRnvQmY5iFwpJH
6rONTst2CdDk2AWkeS1p8UvwbBzHqicW8ZnCgzIgGfgqrvwk9nqPg1/x30uD39k7
8XrIkQSorwmlk936kOBEPTDWKLgpBEGDay4ruxDQXc48SY3nFObay9ZzTnaElYm1
Bu6JCo+TcJCvzprbGfHkRxFFJqxftXekeludm2HgMjyzEi9nuNYCjx/EvXY9xJ7d
EG3FzD7CgPPg10EZWD3nCNp2MnS/SS3/WO76/DdLDbrlwwvyqroWP5ch5N6IWdjp
Zeor8ykhV8mQs7d5a1wY/BXc9hRuexawt3ob5PQaJ2iJdxNifJyluNgq4By4rZGP
eusA4MSA5fZooTrpSLG0mJx7quCcIwd0Ttj8Gfkq+x4QR77VnLWfYbxkIxX3BjNU
2bG8UE4e1Bgo0YyGECklcTj/Y8pP0rxMYVcgM+MkQjfDMREgLkeHEhwCDKE55fvn
vlxBh5zgxRtiQoyuP3KB7qhv/RFhL+eAtuS7Xd4+irGoApVGzfVmQI6pkiOuZlxJ
WSZgKcB5+7C086nYIPPxPuO1H8T/cXxpgxYHeF83/wU/mJ1k090eum8AAvHPNQ4I
yl3dywBQtGZeOlPjJxtejfWGrgRmiIOwUl6fV+FSkJroHE1Qw8nnOFOzjkO4OXQo
9S8AS9MycyYUibVt2jRY9fCg0tomZy84qLw+i1VQrnQT+Pqb+Av0N4xLzEH24h29
Q9WslIoUNZXpasnRy/Mc7RrVFtCQF9ZKDZfs3ukvBN9lq6oYSgBfj+E2kL4Aa30t
xBqQK3BlbnMg9G+jgcDCl0I1IA5gcRnfuYETPOmaQD0WbZ0ClF0xzDGzUwldJtrM
SlLejsYsuSNvCRw962uotsnwcTWKIczAvPZ6mkw/1mRr7RjsI5BHdCoxXdsJb1jV
F0bcq9+Ryw3BvgyxdS3mjUGSqIREyOgFqIgShUkmxEdTYwUGZQ6417aFWOUUPEDr
ifvjR2BSGvmaH3ARWvo93Hbicd4k7GyQirhedUOt30gDMdT9Wa72CEvpdu9oq3ZS
0CeQhPkFcqR60uaurdxDKIV4ETzQJDTkYhYy66cOamdXgTNptJo4B5G0MAEj8Lhy
F9P9Cn9gtLyfSa7FVKaUrn2HWOE4ml3D//8fWnJIy1fYIN0gOOJa5sJ+Wa+BAA5j
vYh63t6J8oJfZDhtCy8z6HUxGMS5boYF97FCbxX7UDnAXPR8hOY4bVzQENaYJu79
B9BOveCuKkDiXaq8tPkD5AoILJfD684nCE6aXa6QdEaa9tRQIZHQX4j+9Roh5G5Q
jiuHnBy4cQL3ktT7UX/nvwBGNjlUltvIGrVEv/7zemzU36j2FDxGBZLpFmdKMJpp
3GrlfkKKjboAOq4Fo/5uqmlDunQdO8gcs93JVigBo11i1Ir2bjDRpdVS56pY3fgm
QRfTN+L09a2fErT+ZGdXTdkxz5q5bdJnRKP8zBmj9eqEHFflTl5/LnuUyfSdPQ7E
YLhSwLbQeitGvCsmEYl3LTOEpOJeLWkoMy08BbHlTm4Ih4gsatYD+PKmDTbY3Btq
O6xjoI6Yv++jow9VM1JNAHXEI9kB7x/yw8b+RQM/R+bOgPoU+ic6mRSo9XgkfMnZ
UMQ0D4BkkceQlTunxA59kx+8dFCbD5K4sD3fn3e1s8eU0R+WugirHmPqVzOe3iHR
Nanzt1jaBR0KRA7OyIrCEIgu4TJemlZMK7mua+QVYu+kNioYR8cQWYMDyMpkZgoE
k2XlMCjZuiIWChk/+Lx0AfkyPJBMc+F1nK5OSvAUV5NDz7H9XteGY882IDiLlsey
dvZOfoXtN6n0UjkhEI+SVOdZM//B2Gs7ZqEXJ5430TJZTRMXGc0FUsf/2QG07Mom
8Zc/6LEdcpwkXoS39goApO8w1n2XxOxB25u6H+1znlMlsrGbUKUdtsa9aFA9KtiI
L3NR9KNsTUL4zaZB0ppsEqBhv+XzNKHGiqIpDGq1+nLqAuIB3gGj/AsNJz0rpAO/
hHWr9CCwDmNSqp8IizP0j7NScuRMDyWF8KlTvYd2xqjt5aBSXPRqgFEsQAoxhB+F
w0fKZGGyAZ14d0CNcqupIufEAOzLfokLP16UIm0A/VmR+2bJUNWowbzMtsliRqhe
e/TwVt27z/61pAzD6SAslLaiB1KqDhebAShGARA5GdsAjMLrS2RJzM7CTjmstRvS
6ikRARkfr3/0dXrLGfLnQdrd19tCwqZOe7n+WNRW+ZPUHcLXHvofP6B4/DbFiPE5
ErkMmSHnPuHoXzMPZO3UcvnR0u0LpXJreqPa5XVsOXuqlqIwERHPKL08hNCj4Rnl
QuyUPjOVoYFS2Yhk1elODk6Tbv7FFfM4a3vxVvjrJAo4nSOrsifPf4tYyw3ffh27
+JeJx8jCPPNWV6ngdq87Ks4VtDl9h3r7kZUlf4ZQzpYX+9le8EGL5I6MdXaDavAy
XPst76LWG9esbnRyVKduDNpm6lXFBxcurruJDXZ2Zn72+f3BZscHT/X2k/F/HYLg
UIqnoCMDZjyeBCZDbUioQGjhAxdhAzFu9hzmRhcOW+sK+uqLBGLUmOPQAfJgMEWR
MJwZPjyooYX1qt2v8DCV0Dl/oYxCir6oHXZmI4EMPe71uKEV7SPa7xjoxx48vxMz
KabkvU8+OL1TiOGD/BCqM4Q/DJOjPVIhk8wYn/+WUH7E0D4GeOqP0+TDHQoIbYKp
ooI7ZjEErtpsWGuIqlsMIYzlAss2lJL69zZ1ozebtrpYPEwGGML3VnTQRU1T432m
RTVo90JXl+9PGK6OCXQEgKRlHIHFxSGdA9LuTd7F3BpJIkoDmc3H/LFZT8BRUuWO
sZhwwdzEgqyiqO1e/ya31/7FBONi5zkUJIjJGc8qRn40xKHA9mZoaHbK+ZWW3tsG
lHboNHPBgI3jCpQ/RaSMa/b78ZRSxD96UBPJlxwMO9oi1id0rGXVrIY2zo87i9EG
sDPpzM9BHF0PIEifC4Ja5508jwfzjE9AJnCBhoQg/draqykhcWQE7Rnv4QTN4e+9
KbhC6wyPmspeHBrQFqrmlPGRk+kdX4nCXjajQA3AnMencOgF8C8Qvifs7p8wIM5G
lyCqpxGHtL20a92wZlNs2h7jvRPl/ou01oa//81MXxmccC/MM0ko3jJUSbaENqww
/flFMZPPETgPCAK/h2v1faz9MO8bKr6JDg0zTREvHecbu8UnqJonCK+xidZwD9zn
/Gh7K3LEGEOB474HPZrD4odHwwK68qnoUcgtRrLpqRbYU/aKsBrGj0oAqD0SDIId
zNPpWKdqrQ+yoN3rl4OyTniHPrHOycXH4oiLxqsTAYVo4D8sgubJbgzI9Kz4y7rl
26qHMP1P0M+e9xtWmWbeUdyGZYaVfW2mbdCYiO59AK5mJToqsuVpHmB0HlPTw7D2
YyQtL12pQq5lRmiZ7KMeS2JzwiEusfUuhdc2ffH/UL+8TuHXp7QRCa/nvIMHGsF6
KmHRUFcqN6kzw1NpaUwrmoMBeBAlaISV7Q+29mfqPM2zk4ve4oHrYwK8DZlAS/h8
S/C98wHNeoq1G/sOWu04ecL3faBterUyHVid9SZscnsC1TsYoCSmLcmuZWIxr51i
LtVcGjyRMliO+Sk3dIj9WJXK1mDNIhznD2aHbG5ERZrrS2UPd/2mmC02A/k/fLHK
3+Th1eCa6YeHaWCBYBVqBCMywq0Db9gv9a6nuelo5m/b1NiakLzYGJYGWKslurYg
i/xNCms21j7BgRNXJhCjxf/88TD2SHC3LqpUG8aPbnJ57cNLyc69jl/1TkTgwX3D
Z5n+yomEAUF+xLVmfe5IQBHjev8fe9FjLfCng/jnk44Wn2z4mw4X+Djhq4Bb32mF
+1z943r+/59u/9uE+qaI70Viamz33uuzaeygj3cQKhKBuKcEY+H1QZHXkVMsUIrS
m2LxXeeEFBg1NmC5EJGdMk2IZNOpjttdrVV87bdyIt5s9e9sfbagu9HWKqLAROTJ
OgXiV9m8Rj1fLbe88Y2cvibPLhBFsYkIIV2CkNM6I8gJTU+lFj8JybxOboNlAAlX
CGnEauSjqP7MtobKXK7QBzi9y2m79eUkuOqhi91EpxmLe3TBOeArRA4hRvElMvR5
JF6F/KFFHIhj5vWkSmiGd+PO/OSHgkfnz4/nL1CaqsQGnd3oS1Qtm5tVriEM/43S
DzTh5rq4WngysaeSzhtUFtbU4KO0hqdgd1QqK2Bnx/ze2f4rZssTVjMVXra2qQbk
iKKoCh1uX3+Hqfys6tBe3M3nz5BVHYQi6jXWj8/cXdvDN4AuqA32oOZEBYgyO7Dk
PA7WvJ/zHISmnSrGpuYJJU76+/OgL5AGCVfEdXNR4OatjgLOBNjGNINDVszHnHqn
XcMCMBpale1nRhunv5VWcFwCdTkLp/bd3Mi4NOMxOMTtaLXbaDNrwqzodL4zfAFL
J/4CXRs2V6t/xfDDuFC/pT4yEC6QnkZjudITbBmQcTWD0YfE52GddBr5DxmkfmW6
xJasqeIpHeP3zUSFYkVoJcCpI9LZ3pHAZl04ddjbPhUtRqxUVVZacJrscHHfh+MK
e/y1fQEKVN/HASPvgnmNTySzN08H8QeF57zcRL5d5HeKaalIZ+BCwWEmx6p8hJXr
3ar5CQ9GErblAE2Qvvfp8GK/CPir4vH2uv1i4/yWjGWUcrXOB60PqF5io50M/Cxk
VdLEXRY94ptAY5SmDRaUSdjVscK5GHf4rfKydgOfRwWN7mMind1emdPxj/NGwuQK
owxbsRCYxgsF3a/yjrkFNZdI+o68pjbMQ1oTh60zkrf0ZIbSBEx4/ZwxDfsjYMHn
WT8BI03WvpUG/O7Uz4U23ynlso+vJs/bsSv2AlxInbTkkSy4nrUHk9jcrYWgoOQn
BYxJSw+ldn9Pq2IQJSBOmGhncss+uhx/GQoSTd7dcjunuX34H61k7JtfPDVJeAI/
CJGwv3OibRNai1h+FUiavddq1BHywkhL2idAU/M41XOUxEKEwzdNYC80gSXey+La
VxYEXmLmkfgjkhJOEC0PsjbebCWina5GKlOVwxQmG5tA3/S9d4mrGBWlOPVuWPwR
rpg1xO8ZQ7wVmoMVNycj7TTa07BmraSOOG1/enMajtMj1iHRUGwppGlJLu0nd/D2
I9EFj+RGTVdinWDMIQeVHw0Z0ezUhrPR9GiTgtBlzrJEWEM12T8GxJ1U2ebkpVQ7
s6k7Km6EOnWzQs96/ZiyuhHK0TU85bKGNkWUnKzztHpDVRqT9HMVGGnt7I+EbnxK
s0MRH2SAtkhQnZbDnkcc/ZX+9rHA8C+7cKTEwsKvRtIBXtfcinwrv0FucOu2425C
/egPYgufetjcioZ8CmUM72Y8WHeDPtdbSMrh5z65wRbct2+9NuuJY0fx3+IpJOnl
Mix35xRuEouO2dVfMNkpybRt0jr6jTzbombdK+dTqX9c4LfieDol2Nqflre/340o
1ZPdM3OBZcBcENkruHrZV/evCjMkqA+qROgGwhbNi04h1ut6yu7nleVAuIJ4Ha4h
cq5GXhrAiUB0U0Euhz5SG9YVDgAZlOIWSy8mGuE+xOq4NiM2O611xB9PMccfJdyZ
QQl2aCrOq0x/gASQcHQ7wFqr53mM7ZUTI4StNg2oglVYdQLFyjqA+LRQpfZ0pZSV
M1gnUH+Tlgq9K8OmL1iY50KMp1O0owusM2Lgv5VmL3e7/9N5qhcHS7pwmJZ1/UDA
hX6K4dX8jwbB4+KzLATz5hpjjatHemqB4GqG21OStf6ar2v24BGAsQHC8j0B34Fp
KALspR6vI8w19PWPZGOMomO4qyKm1uJAuCtx2zYbtqMydvZQKHVU/4DKt/h347xf
UkEo/RIUQc4kMdY/mhtrrXaEVD+Nk9CoO4+lIwuVhkevvjYJ68Ko02qHnyaDr7x3
pI5vhY2IDDNlvUpctLChhNAonxtzkMKzLeAewIIIdMHvZYuMmMA0MrxHjs242ZIi
r94i8t7hsXlN/yP3FVHyff32ysTkVU2m+cTH4dyxdN7P3Lg8BEkgpfZDQlVRX7Ns
xts5UgeZ/994N8iTEf+DrMJAydvjYRReapDck4wrdypfSZ12rfCSkoe3ndDNadWN
6q/vQ1Wfd8g4NwSMbQj73q2xS9QdzRsS+5mR60swOrDOTqH0LK+RIoJwDZ1N8cPL
ASViCc9MPmFSggyOADjYj35v4mOpEjqk5VYN6o6kulB10yb3rrgrdgR7z2N641QO
49qAYC/1u0/xpG01UPf40A2REPmJlyxVUVN7szhe/L6F3oGebEXhj/3H95K6eRCe
n1O82EmAEuOuwgeQN6uhbRicx6u86Ai4oWiGSokMT7Q0YWoZ/xbPXZ5Dfczs2b6h
+yQTWVY3oilBqEurxucp4gxMq0G/P+aB+t14LsUsO5VFZ272AET6cKNSTvZrLcTD
RM5x53fmQUpcPBaooqIimKLsx2zIfqJmV+Pwsu8xco6NqHIy/3xdbih8L/8NGtgv
T1mt17yqFJ77Q1oWKgAa3AJDQ9/wXU2m++tJ1Oc4NTofFYaozf7PakK8gsgx5AO3
JYMEcy2HEXYpBofsmU2RTQ5d668cBN/8R+Y8b0FrRe6UIV0UeQdDRj+e/LBn2J/+
asaqTzgZOBWtXKuVOkElC53HiKzh+90+KbzWkEMYcn7ECGZd67rVjK9Cmctha7bL
bj+a6gw0mpcX1Att5r7zIvrOf3AwRck2ba3pvBsApmnjHXbDqhxIyisvyQ/b3l93
tkGjsh+PgWMAMGpXsoIVY2Ri0MjFyUzRWKRGgqtNUBwg06r36ook/5+W+Tu2UcBE
ZdYEkEQHSsG7wghvP+TpGfTNzGePj5Qpk6BcDpdcs/uHkJlm4gh1OIPS5bKEequV
Ghpo4eRnXt5EVfchTkEX8oOWhceEiu/bE0lrHi/Tb+8cYTRF3Xjsw1qiYx2Huft4
hXr3ieJ6NJ9xKELCjvIZHJv+kC4iR4VyQik5MpPxpzsVnVHVsQhja/069ix19+pd
kLULIySHq69iA0c/Omf16swpQpA+GCFWklZPeAg23AIV79QugJwQ3RvVCKdPdhNv
0mmtPHyYBF6Oc4XcFt4e/5z9MngJV23zzuRtEpAQ6MdfbNKBcgwQguJE28JI7lHM
Sf4ZfXI9Ib/FR3BEdqVceN2U79WaepK1CLfJ7VnNja7JzuVP2+qJIakUo7h8VKyJ
vzfa2V3W4++Who1nWWT8ve/i5nDFBJhpwaOxlA3+ypEqFEF6EEz6jWdGpmRThsIX
UxEFutAhRMoaCvQPFvW40/9SOfQgYdkWWeEkgOHxovTrr2mrMBU0wN4tZoHln6Wj
g0gAMU5ipapYl5BSz5aNsaVVn7JTrWbVdXyWLmZRy/FLq0Jhc/9gOW13hsPy8YA+
8wRrypHPN2sp1IYERdt/rOnVqBuYmAKgQsO5+eABVlVDcHBMfc2x/gIcMOk27+vi
7VP2eR9aJ8QiNs6Hf38qtucKoJONEwOsB817shtX7giJT/v0zTrxOQ3ohvTd0lWY
//Ykfseb64slkFKDdrewUO+2xWaTccn8dcGAxpK+WRqBj0Ju6rt+eBnH+D5rzaap
JgNegBC5zF81AyRjs25cOkpFb8ZqfPWcPovgK89mR7ZW4kSw5stuEBrXZBqAnZG2
kUh3X/kubQ6zQa0Y6Kgc/Q6TCDJ1aAbrev4jd9UHQjQ0UHLKmzVSFnnwPQv9vehl
X81VR+2s3i4oLeH7zFNYgg1yrmH5AAL3Cqus5CYa2zf4yGfMT46d4rXg6MZ5gCIP
XuwBxeityhyrPzMZaFBCP7FOr5sorotaR2d8j/45RU+fX2mPF8t0zQXb8qP2jMAU
xiy4DQnygXRdB8/C6YIAl2h6aNd/EXz25kbYWpwZ9uiES1Eu0N3orpBY+wHbrGK6
ZQL7tSu7VfqAdEnSVF6Elbvn+ORAglOBbFAFoQ1Q+JJ4q7yyvCe03KLk9RHcrdvm
IHOQSngqKQox9Kz3XjCkas4vld8s6tt/BRTWHWESSXEZP3EZ5MmJFFe5XRUYwqpc
aDAtMD+HOGB+YZnHo867SvEKtSYTITlySYK1huw9BwuAWd/DAippj0eqfGQCxWph
XtjFqnGhcib7ozxvorq4faD/DR+U0GAPQcjKP/m1rJ5Pjye2MeDmSf4MGtJLwyPP
1JiCC8XgqLudIRLseacf6Qi5Ifofz9V9iMPZwpiB0TlDFQSe0UUqnpSaGvm2LGLb
f/gfpJt6+rRyKlu2A1SGIyJSq+D5mLRyHo7gGZpBIobt6H4vrA/CApmd43xKHMQs
RCrf0MIeJhG7hF0YQBpthBKdyhOo5UK40g2kxXwFtNVPRPruNwmR5sCUbScPgpOP
HTrtGt+++iZztcJHv0ZE/DXhcIwaKgNxqskqvy3ilyK+wAuqLEZdq0HFGWNEMJJo
9wlToDJww2F1/e/AMONnzRWQ92E3MGtN8s1Qf1bU6A/zaV9NWJjjqImHcsi+KRqc
Du2B//XF0RrDeG2LWmPGudSK/OX9eiHlPzqDfKK6P29agiX8WQkBhsWBgORrJAU9
EhkjlCgI8NU0v9MpyPbvBQjbmKjaX5R6FSjJnbrAwJAAgEMPK+IzS+H9SXyZeM9q
zQyNI7W/CR608HgDDOoV7szmJuni1efEgJ6mfT/GgPaFFTGMjWmZy+IrojvrhU6q
LpWYSimAKuTnfs0mChD9Xd4Vz2e9AXGACbVQztcmcYqEarLzPGcKthry578wbjF4
jRTExtMhOeAI6ZrinhklpkLP2txL0iE5IlZk8BTvsAStc8cxddTATUMdaCvdV3so
Inp7xwkDLYJ2JIHDCZ4jQeZLc0cFL0SysK11C97QgnVhTBgxLWvzj4jAISJlPbtm
giUYZ/zvhEwPQlcYbQCrCZpds2od1Ag8Mb7uXSQeTtrheNhmwYAOsJTmfle7gGYL
c2Ef0RlgE2BZH3yfVGKjtqiUvEHbXmsV9M6XKqJZm4VrEHwFZLPO0ImoiULeJYfG
70VezV8FBCU7ES/7r5o08N9R2+DPdMRQe+wXYlLPkh2xfeyJ6DKHQgRfJWD+Irsd
LRKvnskNLBqIfoB1J5KfXe7zr4VbMAAyo9NesImGS+jE8M3ScKop8oGZ8deY47dw
pH+/qqdRFw0vpTOFZLoreOLUbryht8+hucCKu956DbIaCR930davH770ipO3p/I2
qtSY+3Eksgm3dtf207sStl/OCq3PnLKCXBdFcIvZATKree3RamPdaoD7tuF33on+
QHYnnMsS4gp+4wl8NwbPSah9ERaLRhkCOQ4VU6a9Eonbgr20MLEOhwysnbI6ZGk6
OMaSbfIIG6Pw9qbiiot1lpkYsqftnmMBvrR8U7s86YQEJfe53zHPZH3LyfaZ9Xop
flOOVGCQIAAdzWSgluwqukOp7NqOm4U4rW00YuC1hgfaouW1CnrRhj6zRKIer0Al
BI9wk3ABoAKon5eW4VZ9+nq1MTovfkeqq5jllp5uS9o/kJaw+bH0W9EMHQu9r619
7IftEQ5MVRI4bG69x/Cqp26CmARpiitY3on6Z1kx8+GF1fuMWynm0gXQIIXtSm1e
UAmmf+iI/c+eZFVvd6FgW4ITzTP/y86V0zlALK4T8fT8flzSXgmNQgUQPgQVBZVc
N9gknIcU85iRdblEDV+OTACK/Yq0sPJjGEVZfqPHfYzs2T1AV82S4hNfHBzmZwyp
WGE94aLYwxJBZP/Uf2/m+KztnMplFZsAB9AYZ7y3LbrqW2svq4vEJgog1v1suwD+
2L3QFefNBsqjgpt13G+m/SWgF9Kav2MFkaMLbYDbQnhHA49Np2qpNjP7gS8k5R5J
mcRtoSwP/I6LGyqW2gZrkV9TDx4DVYT4j0d1cnPknmbGheseisTLNTfwGynRo+Yc
zsExs2jy1uXwLGxW3FxYm4dsnyktXHVp3U06IvZYsN7LSQyOdPEJtVzAhW9sb2/x
M+DT1YbvaM0+r8H/dJPHjPHSpGd2xUXCsAQSTiyhvAz7tzJ7idVTlyK7holK8dEB
GNmuaI+TIa0CyYNzhBWQ0/QiTvZt8JyDZdDu3Fo0X/Fu3v8YeZ/qQV2e2P99HOvf
SPGmGdgSO10Zdw4lJdOjbyDxLf6d1/GSsLLgW3p5w2c9BL/N8WpETj5WrpQfocOL
ydTSDCXAVQkiBQuG94U8W3Vn6ZesTcJcua1XvRO035w6trvPxAYD1nIF8mPPoxqE
gLobbn00V1XV2YCkZldwRNEgBL9SkZWKe0La16yV0JnQv+a66DyKqtwSv6voWlUC
pW36luZBbIBMSOJ6ZILHADG9lugyH6STLb6L8AVlb4GJT+ryBTVYdhIpJMAoPG+8
q9lSpyX6Zi8rQ+igWpca4jA7PVSkhCJsJFkoekzMtBx5QeHj/hYlPeUyhMCMR0Ao
K1c7i8U1UtyzezyPdgT96X1nIyaYeNh7Cp2380nTzjdciLpm0q+DTI+JrYhH10pn
iGlEwLXzlzyN0P4lHrthG5k+C80hXDs+Dq1nNyoVm/O2DZtt+eemHpkwYKrYzpYz
pOnG8eUeoUWgacovW7f6j4pZ54loRpuhlTieCPj+4MUUZru2knhRhkBCwSRkaluy
vIKsAGNOYejzB1GDnj6z6Yodf8ABIR7DFbYenRxRoUZlHCtcz7+0RbK/UEzdI/RW
eTwAzPLZ7EX7PClFK06h7riQFN5ZF44m3LYzVkOtdv6m/aOb25jrNhck4b7yHhUe
2x3RLJKjmeZH0lQAmZaC8Lrhjw3KdMiC8823Z2i+yCKt3TI6iVsc1AcTFpx1FS+R
wmqEsa/1Uie0hriUkYUYOTCmCEK8DANcE97pHcZ3A2cgndYiKTAZo1EpQAU22cZ4
cSL8+Rk2kdws+m6fQnsZHuiTePfSc5l7QsPnUSz1YZLRtHOFrHvtlm3NinYtsssu
nsf05Y7oEEVT5SUGj7VCo9IWhsozF7Liv7BsEJCkdmpsDHAWeUP9ZOEuxiDfV1wv
ciqSqf0faK9DshYtdQScaw7gsJ7E5kpxD0YgdDH+FJn4HS8SDxaCPk9tYC6shgoP
jFPxk+KlqkCHg6gN/i84c1UROhbmkSZ9wUqE0U9gigXv3DYpUjqlYMh3AG9HD2ZR
K5dFNjhY92iF4P+tYAOI2l9+xTgXhqq151eUlSGDCzD/ntgf5xXpoVZ6NdRl4B7F
2iGHR6/8XoNgy7wTP99XZfjLN/LqZxi5dAzb/TIgy7CpYSfVvTfjqIowq7rYtfDK
8eaDZTAUq1GOh2OqoMsoC6j4JTCNBwrb0MgOpPW1brGHzJCbDmRvETyAc6pqeOx8
5rpjG1zYESQ6szh1J2co7OKLdyBaTOpHa7MsIM66nrCYETFRSEKTXfPVCM0fmk4u
1UxrsWNEdSe61C7UTSw1jnwRqCcO8Es8qmhZbADDDb4kaPEtSvqUpB9hC+eEaBZ2
fsXwe/2K4qkIky8k0+8ME0VY/HCzPmKouvHvr+iItE+EyTSEzhjgvOzekfjB2a7U
tJYvbcyxga3w0p9Db0L4uCCAzjiHwL2S247FfItnLEv6DGo2I8zrHQcYDsRSc5qA
5WAy/+4OT+d//46sZeoutLs03QdXYXZDaoIaJkKt1g4RcLTtl4A7/3K/9nYlUPbD
M9YyZybdaI0VcFD+Z5nfN5iHe2csTcX9L47rNVmmQNV5RMof2WRZmwPRavZOH9PT
7fW7+y7vG1ylDrmCi5R0n0vb8Sja+M/Fgn9kG/Ji3gdmg+AAHkpABkaEeFQoZVsK
RFygoI4lZ3Pj71YBRbY1o4sIEhYNocizL0E/Gt+psY7XsmO5td8HG9GWT4do32HX
LTpKG6nnuFiBXcpE4yILeQqxlNRRda1GMvCjce/MZtDp7jemqhY9dg0lo70KbtWi
lzEanu14jSr5JI8RnIeAOUvraMROfOaHPZS6oBa4Iko7fGWjS7pC8W3hGnRvBsM+
KrIRkRahOp+uYRybNg88v2DhLBioE+rh7989++H10h/W3CoojVJHUxScTNuxk/oX
rvMgDDtxkdxR1grcFhV0J7lqCRPst3/NRrRhEgCB+oW3FNsFp2Q9hNV3q9xTgtoD
/ycLJTbjN6yd1WCkKFftEf4kzC3enyGzWA5ER/svZR/7yO4ye6DuSWRU4lMzqrsY
pajZBO338F+rv8iOsMYP7RLPewofLkZMa5PWee8jxFAT4lz2ZhjkfOoZAE7TuSxR
CgZpm+Tgscyvt84yuM7JmJp5rYt6Y4aMCqv6LlPcORymvMxsKvIry8NVQla3R5vo
wi3sVc/aE58y79q/LkfiYwE6McBpPW89l1SWd173ch4wAcXB+i0l1t6ozE2kUlUo
XCISXy/Jsh/CafQQN6zFA/tSRk3B8OIOFho4K/a7Wk+3MewMkm1l9Pl2zvDIjKtp
2eeKVpapGr3vyqWBq8JP2Oxq2vmQAlf6E3Sx/notHh4npPK5nz1uCw1okor8wn4C
03x+vxMBcoVCNnWwXTmvHEyIUtYGw9IjHB02F5QkSxaK4T4bJJXLy8neBn0jJ+ea
vLZnvz15uylY40hCzZpHDLqX9jIraxGNKFvI9V7/z6QVVP3vt2BkRoVwADMZG8rh
LfJEIkq79oP8azlmKYHo06bszb8qaP17VcOb/Jz9aA7wrN8rX3xRBc91/t3K8WYq
0f7ncuviOhGX2AYBE8sSxQVr+2r0Y8rSFRjSLMWS0Oshfs4fyOW9xX9QnVUxbIyT
6lMmO17UoATRPxp0z/GkYm5hJHxyBHrD46kBzq7UHEwrs3M5qtVjOhHP0Bpq41sG
gDuiC1OAHguqy5mvlwz8w8qEgXRDCi/2kRfDrevtZzIiE25u25THB57+XwAktJ7d
uLFlDljm41XNpl9DEEMhNtiMUvbjUHZtGqpP7E6yI7A48hPWWmFfCbcn5f9fSIL0
jAQhIG7cbJIwCVGO1rvRC2mb9H63098GDLCC7gHpJV/gUkLYo7jjGRJf21Kq0GeH
7I12NUQC0W0b4FaZkWNDS3IlxbroQ5G3j1/JuvnDU1npw+4XUikvGpyT29H/Sa/5
iXcAOcm6WwN8itiyZJpBG/SwVPIJhVBRNlN78xjjaiy4RCvCRb5A6+ejHSwDGoyx
R0iAib2pIQhNArxmUWUForNEYhDTWDvhPiZu7h+WRnhGgP49diAfMKg+ZrxMkqWw
xuHMr64jtwb4R38z9M5Ba6FJHLlFjojgF5TCIAqj7wiTSneOo3l0rMfotxpkS9v4
NGeNheaY4vvrpVO/oD5ezrpRzCr6cU3th9FTun3WegHlsd8sAi/z+nlIegEy3uGB
1Y7u8+98vRlIfy3udX1jH986WDza9TTaGFFJCQju4jDnrxnYtTQXnsPLuDdcSUnU
4pL18x0kOe0DF3LyYbMIZ4YRDXUpr9cCL/eNMQPbP2eywDlJm21NCU9qttWuQOpj
KaRJ+3FiqZoWLT5wPX2P6vA9tRdwGBaazkEzvjZCbBq4kXWXXZFlOZq7NaRSYX6B
VEedhBHhb7GlaY3YSmQWNl5zBp+HtkNCm1PMbo/PQAUYnpc2BTG89jPuLjQZKcvU
95lwIbAMhJcZ9L2c1Ei8IDUbgBxPvzDZP+ukYhLXgjW505alEvxbOvoWugO9rjof
xpxev53nQhjAtX+ByrbDiRv/5Ls5w8Zh1FbE1xipUzm4unJjJ82qnRXbp2XyhUSq
DnbCcFIHCBs4ex9v/8p6w5nMflBLooaGgDRJ5NoyjqgPVe/Xl5+TgD6Od8qzMAsW
3a2cpuinItm+wOTjiZo9J+qrbvIFl7LhGrHzj/ne9u8cpqFWLC7r4vB3SUskRO98
Ya0taWTJOA4DKRjX+ppGNQaf/sla3kKXvLXSFVrn8JTg8CUrz5b+Il2X8cgSxHGu
HuT+Q+8iY4SOiQLUSjyvK1ZTfcb6Tu3M2s9YapYarz4ydHWFmwSx0CkKjjx7/YOk
gbC2K4c69A3ixP2uWNaNyumOs5auLy7tFZAtoxcAe2L0ronTc+dRdjvVyuKWWcgG
0ugs41eskG7ZzEQmNHyPIIjRgP06AXkkseYZTwCpw5WPry9p7s2Aat/k+oFr9udC
zPqr897BeZtkoPyJ387lCTOXh9rFJAEYYurFB5QBp9EKzZEyxyilTAcEiCwywa/f
Qw490m42ajgUiSxCrmgaM9Gm0r1njtycrHp1NQbByT53SXVmCHpX0dGg3vp5FpP+
rWnXbcLdBQ2DfttRjwY69YCtOzkwMmGw5fFldEWL+e3mxXo2AGXzjeAwi5uZEuNP
0OFCFIZ6Nll1U+imfNMbo990/ti5j8UIpdNlOM3hZUGY+ue8PCHscUlI63dZJH/Q
AbIa4hnaYHofeANgDKn9osOeGHWhociupZ0n90Xy/tWMzbsiKcg8q9c+2AEFrYO5
5IGLNmBOTdSjNFFW4LX/oVxsxQVMB+lRW7GPKXn7Kdjc/MMtjcL6UD1YnCkqpbYW
vQRFPEz5h9P0X4uH6TXOHfJQ/ZgOl4IfSZZx+nYXs6NFJsDmBPgPrb3Fz1bPDIGk
j5x8h5I77Cu+vZVG/2evmnkmB8NMrMKgDkyr6GiFUq2U6/pTYs3uvJHP+auM8ohc
I8+RtPeBy1VKbboe/FdQIOseS7FQ7GSXcZY12Ikz7yjzGnCKmR6xpg9DCItIcrOP
Dld3aVQp+C1IpC2iEdpKGeNCvHLdlZlGEVLDJrnl+kqiAmmlP0LYDYdxKn3TxNMy
chOhg9f1EeGZ5auRUUoLylsuRPbkxGMX+Whz5byOQrHSVoHoWBwXajuVNwg9nUyT
rMKSZbcKXsCkakMXpboY78c9Li8sP+mL+BdWJ6v42WJpLpj3Zf2wRWPd457PQlOn
rHFy6GwuVRpAQa+2IEQEnNUxdO7SNf2RZcL47I0d6gnFhnihlD90XH+AMNl+jcQb
9vd8i2ADYx6rcB0+asHViFYOVQzEr/ediPPDwsxsiXzsewJzVp3PO+kLEZepdSCk
huZQx2IpHPxuFmxosN5B6eFeIuWjmwvbYiuyomXh5en5OiFm0VoQ2nMDnp1ktJcD
Rv0H9XHCLScSPA2c2IYXc/yVsgM0UxZZ+cZbJ/roc34aDM+k7zXxWGXQ1A2a7jni
OTf+nmgvtgQhc/padxypS+6ioFf0GQFSSUqekEQgWCvxIngHWS2tafmo3kwBaLlH
yybgzXlr2QlQeeRi2m38jVk/Vb9yjPbeBPyjQHYxw1M4Kh/iQK1Zd6nu/a0e53qJ
Kg5VDs5SaXfCSuUKO9A6khVCvoEfIbiqBj1Q7RMNmTtiL8iOKoXpUIUzSo1EKdKG
0BowOhTsD0Z5qbS00RdqSgx9CQ0gMIhsQHM5nxIlgrUzVN7b979d0R1rJyCfOVvA
2dLJYcHuOpE0sxAiDoX2bEAemUViME9J+xuJ2xdIca3agxg6hSGunA+tf3ZOeC+y
B7pXNHbdFQO7j5+O9H4znR49U69/yFNAPwDfOHd2NR58X3fTsLvbX66BL8YiKQqL
ySz8XGrjoXCaaKui5GzzWP/o3MdIVMRqrGhH/BouRr3SDzAUvAKrBpAvjK6n1CYi
0Er6+MzBBPdS4ETuKlZ7DIrWUiZVF5HadTHGXr9xUPOc5D1b/ITdgmQlIGcRl0DP
fDhv8PsqKdaamnu4cJ+6IIfaZcK0gGOYpR8FLsSvGYkO04FAkxFl8bcdOSlkw9p9
ocuAW/mF5qkyPsmfZEIksMjr+mEEFE1GLZdT/LQMoFp/sqTPYzebblz6ybVVpLnD
ewVghsg2olxEFDoS97D7vSTdZMPX4xyHCOT9I5jwLNqpuwhgrbWw168APzK7jAZY
XSsJiV7D+65QPehguyarXEAYrDzYoxQiYxHln9otr70IxP9JzrSk6KXs4sVjPkWi
z8+q958hU9PnyUlqzSkMf5dRVzf8TNgjB9aUmx+HBmZjs1irVGOpwPb/9kkcuOOn
yLg4JHX34dwFryrtvjr9DMeKNFarB96RhMufeDkOu6MuFM12IPSuFv4iFDq5frV8
NEDkIRJepOyVScGdiGliSYUvFIUt7O8V1PE0LygH3ZJiEo1xUeQaHOuwJk1pBk47
mC6lHkSo4/OfLl+wpE5DN8fnVyD0u4IVmxnPbo4k+E5bBYjfHb3FwlveZaUEq261
cnx+69Jtj+xXPGw09BAifJ86T9Qbh1/MfZqMb4Rig9UMkV1TSh74aQT3DEweXCvw
nP+MBhiIPZPsLIG2T5SnK5GFnCYDwF6swWAI9Km3TWaKd7KoEGhk97SugwLnj3GO
MVtl0AXCANQGQ7+rw9fUVxtKCHRv+tYpYKqpiWs4NzV3z0DkrHZ+Px0K1MZPyZx3
8gQTcUDj53ivk899iWIk84X/ttucdXUgvausFSmmtk3XzQfePe+r4fBpQjwI4IcP
315qpXj2amxlLHNVKhbp0ZqS6GTraDeFEH9ichn0DOEvkw3Gv/x5cYAGOW8iEX/0
4Gs6sBjSBx8LF+4FyobO4XKPEOjVIQjuTmTVzcf0upMeLlvlWRGMWnh/lwSPyzDg
KgCk16hKPIx7b36oAdlfkoRlj68HVgWe5807kAbceG+YYEIjjI2QSXXQ+IpUxWgo
txjxO70p2ws43ygGSPCaVk2r8kDIHsNJk5F2ZOS5hwtZwYD5eN5vXtlvB44TJ+C6
D48/MASXXXX2ZITEyNkZw3l5I2j/zzlWg9FV0kpve0EohwKczy6BxSlUHNOapuvg
API0MwuTTEQbaZIVXXyoOzdalO8/8+jIxrg7eP9wwPDeEstlyl7uK6shmHcT/cfo
/ck/QC5p5EzrlJ4EUB8PNgaOir7hAe4kUp3CVZvYPqtldKkxty75q40OZVzksWE6
CVwK7MRi+nB2MVjT51IYo9fUpA68VmdrEeIQm3etXKIXtMUycg7U03N5WvpqyWyL
ZhrSha20rLjA34GvOnMYTbXHDnVER0+46ly4A5ffLu/YXlYGJa4FsbGoJKsm2lT8
h3tqMZf4O2DVUxmhZx7Fxlo5HU/8LzKCw63TgEgH+Xw6zC5YIJno34HHdc1T0KrW
ip5yh0fSF60Mehfi/W74oPQ4sMupaLB/y4moWEZ7wzWZZ6Nxa2DDkqjVuHi6W28K
9LA2N+DrlYG89/OorW8ybWW5ipCPvhyuZlfD7DvTKNcA8G5k5FuWJ/8VSwY54C4p
yQWpQ4/z1jy8EHy59FOjp+2NF/NPNsAyRcYkQtFb+Xkq390lNHYYPv9t+jWv1ffu
wCMVH5RiIX1ud/ofq8MolcsKhHbk/j+6hlUNMAi6nwwhDUtiJ1mY4umoLjtLi5gJ
XluObR/Er6x6lO5yt6bOeKgKuwATzbna4Ujp0t9f4tQZ5Z89vOSvrca7lGTPYEga
90SgSNwNHIQ9AnkqqKsCk7dvdwz4J4GpTpa3Q7grBIrv43Rk2cAy1RRjhW+/TibN
IUvGZMaBqobncx2itWpv8Ox2m9h3SlSz/p9iIbxYC2ZYUhIWWqItJ5MeMmrO3y9F
3ms/X/IbkJJ+IdgC4tJEnL8cZy/gk6/6HrruhPEsNUfCf1g2xANL04Fi2w99wSl3
QSMvnduUk8Mfj5WgPzLGCG4trlB9J014VNgzr7+nOn8XMOwWLuPnL5qltD9QY7DI
vXHhmr8t38sZEccIq4+Y24dPGdQNLdge1b3201L1kAlsZvLcXfZpuSYWbWlpww8V
AO443Dq81MV/tkh8RGJKpdTL4sIlHFaBSYALKMbGr2+EDyRHWq0Bpg+x4shlvd9b
/KQIYa594lwzFC8jwC/vSNFi3aYWRsSWKca+/GmChbbLkzfsVSJDcD+lVgxji/qm
7W4IlG6jecqJshTvbWZmCZQlglyTbFAALtYm69hlBRM/pq6H/NuqXiegzDmhQ++B
yzgk8IVia488/BqftmB4oa4a05rGLm9l8gTbirCabxb/YUgu55p7PkLV858fT+Jo
WwR2+j95G8iHdSZ7W3GR/s4rgBKDLO+IwCUBb3laNMIUWUOYc46HvN2ubBtvd6U7
v2Hi3ajFFwYXPocXIX+RRR+W0U6twm8UXbQt0oA7zJlZU1kLZ9wQFdjnuXocg58k
DY1Tk1GKYsWyKLZukEoJ9AuBNY7nfpQAuE29cPLMBoFJYcNfAdY4CEBoXppsWY9h
f3usSEhXe/T97BYdaAmR2gwFQSJbPOGemCHMncAM2e2RIgCcbVf3sqftxDxNnuhy
376e5Ofb/c+Lw27lFI46/8DEsIioYyYJGiukf30d9DiM0puIZSAAWXBoKEqivKfG
gJynLpdboa2uJvJBpDW3xkOLfFQeF1siQAHTwvJCC7WjYPxC26FpBTxrBgqX2cHc
sKW5LZelVwj/R4oWbLTAd1yZocB3rClMIf4n65vz3RthjXwneR2DAj5dqR2L7ZZ3
E83dlSy3twPNALf0U3kLmKF1ruPbqaLwCJ3YGUxCR1XrvEHnOiS3dV30UYtikHaH
OUl/9GDdvKYd2RjCHFxYMOmlB31w4cH6LdiRsJ2Kvrz2JvzdPiqxp49jA4KBZZla
DbQMIxB1CIdK/4nrkEt2r5NtB/A/E8OunVZR2s8e+LpV4pQk0eOa6XkKIthPleoI
uFxe4puxVvzVQgLPive6VNLdEYpd+VO5zQDF+fpBIgz2T/fjirsmhH6K/zG7gW5/
Q7g9MCLJ/id1CJKzGPWjado2lXpScmmEny/o5ylZwZtTUtEU9XLOIyFvAL9XenZZ
tru0zPLIV171/zzD/3ORuhWeC6LVVNbofr7TCimMF0YKVxUMWbVOtHgWvW4Iee6u
RzYba/QXKZzM4/eG48O8w8SKXFohASXlSwGRPUzsRjqqJKVTPH3NJoo8VyMLuu/F
MWxsTu5xTLXnudSskYpW1jW4d4HR8Z+J/PbzCx8Z5G3fx/aiqQjuYaP8qvg9Q7fO
veyTN1EEP9CyFPDcE/Jhs7tpQUhPJBGl1Lq6qrvN1eTGAx4j4GYh6dhTzzUABYqD
4fkjQ1d+zvToMfohXRNuMGzhhSkWEz6gBrmZahs86aS+gVs3/I/gxghrv536NOlk
XQb9O5XfoRazjL2Bq+Jt+2GS01SaVRHGv8LrGwPA/Ui/FOuu2LsoQCb0hcFsWkJH
pNHqmiZf3yTI+FxKeiJTctTzfBZd34CFLxsJ3xlCsZHfTtFCTJAFrkNDxuIFJOiB
keuPhpFvna7rQGbV1xTaCL6p8trXl+Z+2nna7faH/tjC7dTM53PX+UllBiSIBKGQ
9dYJgOaRoCgEEPLHhaMscx2l7UvGKW0hS9be9d1QudLK1uymEOPfwGr0HC+ds0PQ
5YpW2uax6CiPCNTpsyHIHyNzQCo4QvAgUHc0dHc/9T9k3j8pakvYx6dYfqxhAqUn
NF7ou9L9uQCSR+QBopv2aGJc3pQ15ttTg5f0rQRn5Km1WSrMmW6O8f8khkCRDmW6
v/pR5KrvxN3wx8wKEiR73+DFUO1pXJD6tDbtZy09yZoktXImga6MiiEeRB7peztv
XWA8yCdKdvIe0eCTWvu25t9gWD3ASiseFcmOyPmDQFcDs01XmMeHvvaTgqgr2uim
fs2fzkZL/ci6CfzZM1lhEHI/jGeamqZWiMZrdKYQTBPpTYMz0WBShx8qp9TEbA+q
Z0VM5SfNNmOxqF9mYCZBOffO8NlWMFfhxGrXBsUZtDi93Th3vPq3QPd1aLqJnIuc
2uFVezMH6lkxE42RGAH+8sQsOhIUJnBo+pmIvqVeoVP4c99vdQwg6OiSyTzMVi/A
zv1n8EsKe7CVqkXG0geRnDBoj4kKU6S36TSKFOaU095qO3pZNctkAdNkynwf9tfH
Bb6LtYjfzvSe7kU/i1x+Ffynil9NbzGcu3XlSZF/VA3cTLx2Wv/h9/ltCkfBRcCM
Hne8/qcL4UIRTZCC9RDXxfnNd5Oshmx9smlwUts/aAiuydFJbon+YDVAkDiTLhbt
U5j/5zVokZbbgzKV5Es1mjk+nwZtnedRwJrsYvuwJoA3X0Md/unazivp5WiGDfuT
DIiRHrxMiDGLbobQ1+bG9o7PG3zAEiPP5iWBOg2kW05fkz6le2b0f7LsRMOZ7uJL
nlQcdIl4C/KKR5GTuu2tF+NmCdoOPLPTJz7ygGjbH95mTk5nwSDMAga3DIsEMb8o
Z6lLrPFPFMSGUEy1MO4+gSprp+Ez0rOOP3vcPzO7vHzbP8kgs9LLOcWIP0l0XEpw
BrhJGWSd79QMVtsbYSjJCOJTGiWlKXRgwjVPd0qvIpYoVJ9/2vzFFURggVtyFpIL
rqcSqyv11IvqCkWt+nFr7k5DEwGVWwNWzuSs41pbqVA/JNcHHD5tMVRlbOrYe0AY
KxAqF7Rtl4kSV/jmHNmtsWnX05sM7tiGcslvxmeCfQQ+pegDXamLznNSbDmGVYEi
/Zng5FhLGeoErlnoRXYndpXYW1X5qlVTzbmYW1zD/RgiI86bmJuxuDxRUF5U1nf3
OEX1IblAa9biIrfi8SqoVvU1JQlZPcdgTrsnP9O89D1P79yr03iOGHF/QwRI2q75
OdhTcokvEMKbsZNbvFzWPPvtN4BDLXnYNzBTBGQmrnGpoO5hAw/xH+mIjLpVK1WC
XAsPtX3p7RTciGaGWitcm0vbMc14vQSjTAAMTE6HwN2kstDfxOwIm2wNrOhiAvVq
VefsuiPrGynlT8KZ5WRQ2pnkmQz8emC1xngs9Mk/CUE3L1O58zEYQ8mKfdfXGnUe
RhX2QaGjZiUqvlL5b+2SlSGM+tT4VV2MOS6HGiRNZO/Abve7f5OJmuVhbBFXTdQB
GA+EvK0yvypXUQ0MimygHVd0Hplg1d/pSMAhkLjFGtBMJIH9bOaEf1aoevA6ASTQ
EgL/NnXGbuX001FxGj1Sw7zarkKuBrGsp/l5pzBlqXxweKgA3XQtCHEnf/9v6eWG
8jDGCNVGkbfgUWHFwiB59qqgEIeh8pajBWO2IqrdDYmFQsTBnb0QdbLlvINVTXjO
36iJ/XvhSkwzM2ZMomFqEn2d2beplK1HgtiYDZlfRQdzfASn9TMu351hwjqLyAEB
hlKZM0sFmvtxbHIPbsTJCFYgBOkhF8/mzuC0qyJmLHFP+NXcaPFtEOyV9e8ZEv6m
3uzb6YioM88vllvSHXbNq4nGITtFqybZbCZ/xqB0OtrK6yAjYADLDNNOXVFMWLKM
I/HVca+JNOHvMWQQ07+EH3DJhxJY3/MJHHeYblWXACBqFOkE6WWD/6jSRRHME43k
kSb0VkJ94l4/4uZYpOMXyVXbUKpf4WOa1srOs8Y/YFv4I2Evuf/HriYQRhruxUgn
HU1ZG4FalubL+li/I20gUY7e1xgdorHS3zBDoh0x4oRYg6vph6pdmtoFxn5ZRiPE
lUwUp01hy4+ParMwEtPDv/JusQh261nYxesCVeQ5IBFjjDMKX+Nj6m41tkM7/RH+
gip8Ev+nhF/FyFG29mkul6qFUqa8cdd0YsJjPAcstyUfGbsHeOOlj9IdIYHdwlY8
OdRPYKxkv3NVDIhJ6rGaD2hLAwKsacZZAPs8xFSMORtWXQ5lbEt1YO+e2oOAxhSI
J5wgTYIoyDaTq8EgxC6ohKHMktdgvbCeV9K7/0JTtHozh/oMwhVPb7/V31EHNGsu
Eve7hXfNqqr+E5J1RUUiieMlB2yk+imVvVhPJJtQVkfXc1jqsgrObuffnlAPIp4I
p8jrErKe7yNn9IFJMxjH4uhMGV3MxBxBoGlLcIyy3E1jsNmkm9/x5VUNLCHVcjpU
DDpiccNS/ItbgkjwKu2XiMw/RaupIF7MrkHPbS7gwccVH/EfTInOvkhU3KIdWlHw
z/WOo10zVKPp90HbjUMSDUCK5Mvb2kiMxXoZpbB2fnqYb2Uc87NhQrhoPJib9B6R
nomyu9SRk9W29t17QcrT+KDje9yYaFVk2ChFMBKNUo6EehRedueC2K1oGh9hxLN8
mxiblzNV1kLsNP2ax+f+eFunkQUeCNHRZCW9g0alz7WybcMaTHSUtlb+Q7Aia/O6
nwxmHW06kWnoWrOjsZIdaiadumWFs6IAozuIED0U8kANnRhvt0Lbn95yXIQC/zTT
+xbd0I6NXoB7B/w20YH+TYTVMs3uB1Ppfk1kwE+R6XD3dyaLUGtaVL9my0uZAumu
ECa9xDESMIT1Rc3L1pHOMeUfYHtjX7REClc728hf54MqbXAOLXiPE4Ds9nO6zmaw
rBEIjKgP8+1AOH22mwZLgmh2VauWlnGB7Ie1IldvuFVwsZPtShgClSSiIfl3VTb3
slSSnWHOz/bd87pvuOYQJn9NcCrlsViVRrpOrS06yhdVlMu+KwPOdZ8FAI1fJXtv
X/5JThi9gBkjTt4iM04Bj7WiDqdWjl6Lkm1qd8kbq2MTdyMIRJ9K9rzE+8Qk8j+9
pfKeWHvk98JSyMlwq2iE8w3lQz3DUPBVASPJ1znXbJ1kn9fYo4DqQ+eQPjVm+F8E
1RSj3a1CSZqNTjRf3fVGzK00pvrsYCArfM7tvwZ4JD9CstcIULU4/Tns8agkepIU
CcnW6ZAQ+XhGqQTej2fjo3a7CHoDPBGHdYLsyyMz6jo6yxaJU9J+Piu5BgGvhke9
7et1sR7TNXQAiyy01o5UJWLicLOzL9fN/bWK430RSC4IrgnKHF12mYVhxRDbEu3l
ZCQGV7p5SZeptFBGBi3H2B2WRrDTZo8B88n0Oo3jBCMCAtHsX91Q5Cx1WYwe7+gk
0650yXiPon0oJWvtaWwVRbrF4BUSP1lAmTtdWGSWdU5JGv6A9plSe15aKbXEIObq
B6J7tfVbkCSpewxdW03pyw==
`protect END_PROTECTED
