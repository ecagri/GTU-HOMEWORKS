`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JUevk9WBc8APZ32SMnYgutXuS3PQ8nJi4KX3VRLFP9uWZZeQxvU2vA7yuFcpiWFM
smzXaR9BpUtnkQj+WK0CHV3TnXUT26vYTD7UKSUI8TuZ02jYt1eHLlMWPQyR/V/G
UatuKViLoTDeJ+Q715tZJXQ+UE6igs7Cm2psT8mRZV/rd2bTwUJimRvJe5IFrW/u
h2g1DdRw9dIGL7Tk7vJuFf7JRu3zFlUBFXOUiCfm825JSXXL7f/4uuh/kgEMPDZV
jP1Zdr9LAYAHtoP8WegpdG33Lr7BjfPm7EemdGxiGdQgOwMfdJwdOdHXcmzD4IUF
2wfvj7dSETXYV/IDt8vknoa3G733rVuN36UZjR3x2Loi+yBzPGDpulzWuDCWJeaK
G2Zo+bGe6E1hACZd/vChKL+f+P6lWJYjGxzN88ggUovYrNS5i5j1kElPuju5F9/3
5tnSxdZmFXJwTftVMXOmUi6Kv9pmIts2aJx6p0wGBc6KjzictwyldZPa7hHEMC8z
RZXHcZ4HDKBd0Z2OhHyGcPzcHhWowcAkKUeVbh2W/psXWHF429yKWel1EyJpx++Z
yAvJ72LlUlWAvWZGImEDyBy1fwxtt2KhI34YJisC1jf+75VDJ9MjGH0X8UA18LXV
P+i1YowL7HcYxnLQfav10ZT8s2JNcvRFOG6u/boD2gHXVrvNQv8atAJPJbaIxrZc
PGDmDSU/Zc2cZrR3LgM3OfUDCb3RGiG/DY9Jb5xw8rspLw9hrXxOahFjFz1guUJI
pMrShVM9ZKGUdUNAkWv1UONChFGN79JPlLkiNeaVR4oLVFZoMRXG7uIw16djcEqr
CvQkvRtJCUkW9c31osU6MiMIucIsMZsapu/AA3GbpIiMMKaAi3MZuYipasdJjGJO
Rb9vH/5YNA5DX4Mg+2dILDp1NmEW3QnGoU/0rzjs5hfB1kBoNzSzspA0zE2Ue3vI
EXoIdawE/jSTPUwnzP2yjLu2oVr/HimUiM8MOSjkcqy3CXACXwmauj/7Mn55Yszp
kZ0VVKB4nnbhqrqHxnMKGqhL2lpk+IxmvuLFDQIVd/1FjnWKthjm5mS4K6qdJSo3
9b3LHdGWUSXfwSX3sVXiBK1WFfKFGstQea8FoOz6aU23kdTrIjkIS7cXiID/Bh72
qYc2Sv1eRK/zgx7Jxglb+T/yhjr5Fsgh8bwkerSVnJrXsjF6oxyu0dBsVumMKom+
d3UWxc8EUHKwbPLZ7+uagfsTPJAVOre9SaYazNiLfP+UCJkIe4k2XxqmlP2b4cvl
TjqnACG4vyHxwYcn/8kmoY4FKdE3vZtoxUsrBN+KE1SJksDOXF4eB/4juArgPicy
O6O/E/2MDBTUJB64HHcNdMRM6yW3wnte+C/tIvN0RhY4jwA5TpUat5prFkwkcgzk
bS3zDOi3wbuhEiIIQ2c7Rwt5qKJD2c7lE2D9Nlf+ulsVBl4Mx3dUHemQVbmk2FDZ
xSB7YZjSj0W9XIwlXpKkG9Hd/PZSsJRO3CHrDJSe/w9uc4Xoisk+hxV1L3CxbG0d
MMh+2u8+SC9n10G/MLUaZSrtEpiZgLZoWQ+pF73rv4Q7Pa22Y7vskX1RK0gCxllN
fuj4qBWdvp0acJ5tGZh3UyLPrIBz5NC5rHOZ3C0hPpOA/cjAidcza/t6bsDtXPW8
0R3xT+VO0xff9j9IXIyRl2gb6rO9SN7Fyyt6Vt2IDT0zpX1k+lo1XKm2zvw61KbK
Vbc/K3taCwOBsWw1Q0uNTCZ2IYv6b21eHA+Qcu+fITrqCrNvtQdpNz4Wn72I75fU
l554wRcdqp91oDLQhq1t0JQLQMimiQckRAZsZ9rnFDz8TwLD/IvYjAyNFM0CeDwh
acgDjAAXYVZWTsILKgh/AWMwOIEpGeNETQmWVmJUj1RhVMwAnxfCDhSiVxehMN6z
BN9l9sYZbGJyETtwjoaUckTowFL06BFoleYgceXpxTDvQh+xSjZBVCj4rs7zbYmM
oUACibVBZGGRMb/9mPN/RHKqjXGk8SxaPI3xf7e5DX2SF2vnR3thu+J6klVIxrlO
PAAGrqJakkKImoUkP3vRzb9ltSbw3bQj8p/aUE0Dzn4VATjhSMdVgy3xTJ6DzCv5
vO3nIDMGlzF2GyQy5CEvODFMSvfwoNPqpdm/miTMZiqvIF/qTX4w9uMIlhOkVpjC
CZ3ZyBROVSrAzo1kq+B8upLQ/8b6fHFjBE4fnnd3cPm0jraw02z/N88f2n8owElC
wdNXXxS5Vd7waC4WQQKMxJCDFlPsjswPT86s6+FjQo34jFbeB+tEL2bQFICUHSue
lK2GX2Y32zQ5pecYzRBor9kxCEY4sG6m2gHwIdlXmHvyoLhP3DVdMYnkrAdCVQ6Z
C1MbVktXvUBEvQLAuOQUg6mk1oaJz6EKUvzKfa4zkhzt8mR1eU7sK0gkUOQI9nhB
Ktbe/MvDtyBqi8cvKeOeSR5/IFTCzqf0I8RXiaRcRiSaxjLQVFsHlh6iL9+bsTp/
geExEmWalChm75G3vrHjRdOo+Mm5rJATWhyw75HHRkdr3ACdDbbmvcSOpHoS2vEo
EXLRkMtxuRI3S5j9jHy2hSU/HEwBKLeySBqRH5ANmk0G6g3gih0OoPFE04vrmpkh
q0cRPTajsVmooSeDyYXdZpfWQ+sOds+FUUtp0Yk/5uxe1RkGPlKG+hRQkPd9zy9y
Laj8TnYeo5A1Gw/kvqOE8XgP9VK2x17rKQcENHX2QMt6x5jMy3/gy1MfaMilL7sB
1RillwasY09XlrJxiU45yiWKzP/oksMQf0gAwLXIDjycdUwfG7FQMvHDbJUwtInh
zMH1nRrGGs2ikRXVFDt8hqXT9yLzTyiAotaUermSh3nJBgVw3SWMeoZTD5mv0wHu
Xw71konBJ4jJ1xTSSbxHwZ05G5OtKEAG2JyrvVY1md9/sp9thEe6Ifc/JUVctCFn
Hnfkc3icdNk3bbQUkqVPHvkxuvJlKjPLXohjNqj2tntuSAbsRx6GgQwS8VhYQEjO
OW6FVhLD5oRLe9LPGX13u4wRjtjyaktnLd3/QDT87W/hMK0YzfSRWoNvM6tzYglw
XPq6WoCb0ULMkFddJ01lZLonGB0U3yfPmgS/NbhNqGHR4UwHnJ+39cx68q2F0L/W
e/B9k+lYNPur9VlXJ/UsPBxG0SYRv2UOStQfHamY4KAr0Wl6j2m1QS6nwIfe9b6U
CELDDC7RUUcvde8NAEsWEkTHW0CJJC5tu5KVjWQoE21HtcDuOymN/0loMVlh+Tdl
kBe3b0yPaK5Qy4kpZGP4yhB+Qgd7vFfak2JwKfs72DB9GzIxKc6ja8MrtNn2j84Z
TeWyg4qqG1xKNpyn34qV+ITWRWhsRuChzfgWMFdT0vMW2bpqOaS6KRs+DkwPLVp/
HZe62ekXZUZouFY1gQvYPHL0JLs4b4jAk+Rx2JQVeyCiECAch7mpBYBKvaFKwvtI
FH0L3Vud0eS2oICA23aV1/+M3zMgL11Fek51RlYi80JYCyIYD/LTEA/gT01rXCkL
vWyO1oilpuIVGFt3XFmQ1oMS22MmljNkX3A52b1X98QI21M1KS55d0MU8i4DBL2k
onO4HSvD+QAZ3shtiLgMUNW+qoLWEeSZImKlCLG/zkw6uGY5wdDocdx27/sm+KqU
Rg3LEJHvGW1ymSK7zLgWADVQZQQRDoScQsdFRSfkAgrvIQCawOAYepKkuNEcjS77
T+6Kilyw6ZAPj7Qxy3IgM7A7cKChmta8zyihoNFzn5BjisHxjGjefeLcmSmmn11u
gkPd6ElcsnvNLEEfc++uI+KewgburB6tGdgbZxx4M9lxA6+g/xNWiqDUws433v71
+gN3TuJ4qpMa3w0iqzKwNY0F7BYc47/Rqqf2swckdmxipg9AKlAU4/uxVdyGOoYj
DndCiahdDore+bXSv6lPBqnoZSwAZEdtQlTpriqNN/PkBNr0M1Kdfxa45slmx+zc
6CuGjW3zkBtVNg6XDCqMWQmHHOC3JXFb8oPnPHpo0guxltTdwtJWD5RI/Lf93yjA
j9cIazUAhIzGQrJ2UqzwZzoGZ0+rjtyVbqhbx5pJ+VRpAKY95ABxg3zCkSXzD938
e+yDVQxpW+bN/4Ze4GBPv6j5OyjlwmAHFNr/G6Gn1WdZpQ/A6ZUyNwle8NTtBWn3
4cBWSdXPOVzrtpZY2rnKis0ktqX1OuSVbIuVimH8rd23ZsXn4iK+iAmrCB+3qH+T
Qkug/BmM7uJgcRQJI+cMWBjQ7+3GXyJ8miLx44Qe0re9Vhme105bGk4EXIAKtG8a
oEWFfyJUj0dBuRisKhPjJj1PG/+nY8jmJuD/e7aM0LAE1ORJE0eL7WbYbmuYXv20
QmCfSUT4u9T8tyae2gtcfBNmj4iKl8DfKODdFEOT24z/MRzky//Rqp+D6DYeCF7k
8LVRWfJGSUk9z+ZRDA4E3vgLLrk47hFo2KfQkbR+DgR2XjQqPzYnMwTjCgPOrTeS
hJcElPa6x3DiFhemWpPFOLWDMb/I8W68R0aYh3eLRZFYgmPHJkB3sqrZNuC+POwc
pKzYerXNvVp0HPoZhctRvJVgbMa6FisjKcG6u4avpc6weAKW2Zy41ZaQZU2lYFJF
Uqs2JdTmJWxRODOBPM5yvV1bTIzBhgJhGLnZ15DRjBGUVUVGoHVIF1NNrEmzPVMX
zgScQ2Q8MBvaDWOeztd/g2eboTgILv5ExZA/93M6hftNaEVhN8b05qNosjRsBh9v
ie61jbVXYlnj+exazVJaWlXuhSn8MG6dMFf0//u+xSbZ5eiYYg4yaZfW8Qx63wTA
c9j5bXomWYA2gjh4OFOvVk5W8c8A26euBx8ymNugXt3DrWN0SxzZJ3mFsNsPhUrq
owlJWuQe3It01KKxY4EuAyZWUOG+D/wYVr5j/5mELNcOUWHae0IquuHp1MN5LntF
e50I55pN3737sMEYdA03mDa18QVL/HzkrfO+Cb23cGglZG3LFS0PmnIoYE5yqFxM
CISwPTCxgmjcMUq8MhJ1to8+akF9uwB4IGnQWXUn2TJ8V7ZjIfZ0CEpebsjX91DH
M0zZGqyU7rUR0Q0S6AZArxeK+CareTN1BRq8u6AGxYeeLerkcCiTi7JPN5Mq8JXN
a9PDIRpzMTih4+PbN+sD91aCfaTEyMQ4E4E0gmlZjnj6U5DIWlF7vm2uG9oz7wKL
yIEoO3NCUUalCN31n5tcJKlm4Fy8zUNf+hanK24IL59sCFD/AEtK1gDm5Owd3U/6
Keef49JyJlj64CQXJ07XVL4NhLxxQvlSNhb5aUtV640+hoxuSShFlB76M5TPPXIA
LWpBmEYm3n6kcNdkfk4bi3bxft4WD89au3lpGuv+3UGMz+I1dXYQVn7+ElkXAeti
XgXbWrZNPpDZy4iqzUHsKUBNh3op9AlbxwWug73mVrwxZ1X0Vx0WdiCNSM3D5LlS
TOVbukDHHQ14jV2OUNRYVvycAsW1o16u9WNzVLT9R/xObpuPFDNmqiJ0pZ5gHsY6
2PqYAoX5dNE+hV8yeKeO0WxFYRD8gjlavS2++Xrl5PfaZGcjsFGdWoLtk7sw1bPx
OQF1ZfQbZ61ntEll5FC7417qX816ajqw16qrP3Nvk7KuIRHYusWyT+hV9Jd22tsh
unL6iGQfkcSL51SBB70Ek/2Q38JS3qL5rgDPy0n5dhmc2Vxf24Tx4krX6+eEbn35
EDQBTqFkBPGGhWoRIg7BXn3go+wkFCAH4jzXumOD6hCqKsZalXROo3eFpXXXt0je
+5XRpFjxnQTBkbNqr8+gtIukVQ+Fkg0Jv56baHDMLKNF7z6RCih+uvPQXbRi8sg8
yaoJGD34MFfv3UZ8K0RWdxjSPKqc9mfQ2ClHbqaxw8DiNajY09UTi87TJHQIWx4/
wvDC0whw6MoK3qxDZMnz8Y3hUKNAUwRVFnp3zOt/xpMgaHI6PHqNvMQb/PBrfoKC
ehrpznjKP6LPWba5JgydXlLOJ1s7QcaVH03u1ahsH+m3/tgUxl0uQrK+nD6q7TME
R5sSrFZu/OYGnOP7aCaDUbp+4n1n9yBBXRBV9H6xeB/qQgE+NWEaqIZ3WSfy2z+5
QtL2mpo4E2jEixQTNwLfZes59MlwKv+AXNci3zg4U0iDSYc5pKOfoPW3V7ubF1N9
BexYufjvC7cXjEVrt2Mtra+wSd/WjA6hzt3P3tozpkRkUP3OguMXCxy9O9aRLHS4
SsgvtXCaIyyLMT/Pt6mgGDpPF1KzzXfl3J+VSeQXlHiASv31oCBgf8L2VaPe4EbF
RfM/lcnUdo/3Ha5ZyeL1rJcmRbHiq0BtUlILI6MhMa0YnBfa6lWkdfu3O23UAX3n
dDnPpk95684Fhml/zBb/ho38qOHLc2Ync6K0gZfcluZk8c7JXkKcXk5xxznUxInE
p6bSLk+Rls7hTeoD8sH3AbZIUrL11IeLEfo/1pcQ5mWZd64GgI8FjuAOxDCJvqdG
GAuq5rKTAFLEk+aJ8BtIKGJpGuiDnD7HDq9uNn2s3CNwN9n6rKCIHRKx3v3Ej3sm
VLcDM43Yw6DqabnSmgxeDpwkT7v4DzlFnb8vjDPsy45ovo/FAAfuIPCH0AFYf1E0
zPqLeXLw63BO+ZlIGB/6EoRH4tRWcbf+p5pDfqpWWcGBwYRlZsSMLINVq/KZGHDT
5q3EPM0tLVtqKpYehroe23Z4nCnxwg5raOTLY8lrN6sDmbptypHxpRLvu4LfNkpv
qYjVXz9qqfveF6xIkzDZEvr2WcONa/oGbDWu0yEaFTMf1s3WQ9b3a/Qucr7KbeHb
XNMZucZxMIFLCMEYLL/oITEnZzkyA8k8le7OUqGD/XEErWo3JzAiKRCqb6/37peW
q7qVx6LlCSL07JsuWvjEvtnja60L+4M1KDLIEpLkIXV3lqTULQDYyAasxVsSzuPS
BZWeTCPW6W2oyl1NIQVKyNvT3onGU8i1YRqSFztVul6HznKk+aaYh/s9SaBqSzQg
/MJv7S5SdL9QbT9KaxY0J6jr+nAdO+vAPhT4oyRSC+TykP4eMbIccHlUZQOUPz24
Lgwv3Xm5uI/kPOgOIZNE8QGMvtS+dx3KAF6s0y7mmpUz58YJj7WFS5C0jItX/oVc
BcErgq/BVPrDTc65AfwuMjiS7BG0tNQJKVWsoGbsHafb96yjxdOdd+oJgbENIkyb
6DMnVvubg/OPjQbXMzRfSIzV03U1LEfa0Cd9Pm2OHj7G1yN9tj7T+F5SicWWfl04
WJJ645RBi4Q/xRNhMulfbxA2ZqriTMYreF9kdXiMGVZ6fmTnVkh8xXQzS80KVjTb
MnYAQZgPXplQfmp5Km5jEieNV6A+rICiOd4j3B11V2HActLOBsw4Sr+ID0HF/KjM
iNoAmYO3XiSb48OV2EilJaN5anj0lDRPMY5tHM7HDqphA5w4rjYXh6wswOVZgd/j
8ZNFijtj5ee5B+ltIfjkT7tGKi78OeftD4f5bA05n+bFuEGMVP97aKqdJKcHOM59
d4Vhol4kG2X0vxix1DC9CyaRwQ6Y7JV8HCOO5eRS101TQ1RoBwMHVlvrgbJtBqm+
kkSpscLYq1lu5aybJo6ATMWa9gKHXf6hT1CvflzUTwBmc8x+pI5Vw3azXv1HIOTQ
hdAtg+KOVd99N3aqR1tGfBqpnCvdXMAQMS62T1DViRvYBHb0sXpNPypn7/Fp68iG
gWtg2EYnmYu39cBB+bD1OrnxyyMqk3+YlxXpuBQJQ/Kpfq4d1Mf4wvYkapviy2e+
T+WwD/UtvZ7fIAacnqij5hYpfhywLVPJkez5CCi7PHYaAqPAdVDEDqUqqp5zTMLj
tVV4m/F7zWtF6fZlRf2wEmBXx93Qy6K8KqJWirTOziQPH+0k5pQB6+zyVOPWvP42
QoXfXXKvgwbJ7NxoUDO19/obZ6D2iQlcdQLm/X2dC9lMXra6dgcGe0SAI2ghkESI
6VQYCXE/ozCBNiCkwON+NFpA4hPHOjInRn9t+BeWak4NW4/K9pvT9rEzUQh+Vhjh
1tpRD94mj8vE1pOtAXx23kCNHHilX+PrxshYqJDMH+casBA1nqWfjzhpZqy2TF98
jwSRnZFzRZ1c3aCyIiL8GqpqYBDgleGEE/u8rVS2TtbRfxSem6VkZO3YhMOS0NKU
CwNgqcoNDgnVhFjpkYfDemx09ahaPr/nBFM+hnT0ku4ICQp/h35RBs52YAgItCZ3
ElJcGN7usHWYjLbu4FOKQ/kGxmJhxqfcekSbiLhxvfu1/zSGqJH7N3wCn7YpcV29
OAkyasZEHNEFBDmxlxJFG5jDv/oPLqwRZFJmGFXpCGAzvHXneBFznK8dJjMzgdh3
Bn65XIxC4/VCG6/89uLHMb4k9wiIVtDvzFv8KYChXfnLoAaCqoky+zqLv2eWRzNB
qNIXSdNLNHsquIxTKFOh3D9HhJrHMjffTALUxBgjDKBW77gABIgp7O1vl94f81UF
zPZShkeqT388+4jH9y77XUsnU4NCgoGbe9ynkhiiGTKkR6p+iMneP+OUc5divI7m
aWqDaJ340K1/U/4wgde1dbz5at3l8xpCgtFauFjUBqUnZ1whQzbPbs95u2PVTTZb
7NOcDprL4a/ZbvgrnfTyOL0qXYCFAjUeQYWAmOacvbNt4YUYBvDDPxIQOWBKlvpW
d8mOqnwxmPkSe7Ga0Ry9yK3EU2w+eHbmzHz+FZsm5QKqF19PyOlRv3aXIbYoQzwM
DlXqkxkwG4Ma9jbbQh256KVtgtMYfKKjVCZCavtGbm4O9om45TyMFgcyCrfTLKjA
zRjPJs0TBgs4KWndldeflf9vg4IQaBG6XuFUwrocintAQ9JWg6hbwazcEdX8HELc
VFBe22bUzusNLpKKhqrsJjGCwFqBjGbFb2OzwbrfBlDg/XRj4JF5yDCaMyVtdq/1
SeDFm3UVvNigna7SqwuaYy4Ldk0j660FmBnG/qVzSHpbZEgdccDblTD1nam7hTQZ
LmnBwsvOEtVqfSfkMYXBhksYPAMtYp2Kk94JoGms+QW4khCmcitdALkMBNqgeFcO
BTEx96wPzvIzT/8fK1hZAzH4KdC/Ym10SHI3L7O8X9Z1VAdaTxCyF1hpzimzD0Z/
0m/4K7VklCJzRPITf3NBi9zu0VocfyXrvPBZ9u/RqUtu04EhCzZwZ9zH58WpuEdE
1SMLAZBuI2r8tzfJu8cWdtHftEoI0UsFZpapZW1NdTb2FGyBxwy9MghsXq+tb4e2
lZXYftMQp1QTFtzL7mIBCC7xKov6CkR+ZHuz2QIHu5x/BCTlCxMHgjGLMgPZPHh3
zlg/A+oBwecoFEINFRKKm1mczEdE72pj4I5doHqOi9H7BPoyz/2mcJsYvmrAKojv
oBu9Yq0pTi5DrqurFbmVl+C/gDsthX89NzwrNs+aDr2FDojcRWGN8RGJWyvLT078
DMPV+m6qf2j2fuODczzNBvQAoSwOdHV0bpyf9Vj0clE+dOnklX4pcyCWqCllI99s
+4ZMzlH75ie2+3svJ8bcYD0GLQBvqytQanKk3AFwn9IePBm1Tdo8nLpr6xiRh0n7
nvEze8OySfX01Fwf0QvMAa3BLoSijQohNR0yM3L9oS22pmB+n+5conlHPdUDK6i+
J+Vss6JgzZpaCebngmsuoPM+ngabTK6495aJQEcrLS9eioEIVsy3wdk6YGMtvIwn
`protect END_PROTECTED
