`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TeE0ah8/HtGCGvakxg0sSH8bz0y17+eUTQyOzZhVXZ0MZKfBEZe2m4RHfU5CLsW5
0bJ6G27brt0kh0cGho0L7fsxPxOJ0rvGuTlSqFyUYX2Tdo3AJhZ/5YAedm1gvHdQ
syDGcJJSNB6ynzfktIWYgpYFSdUSqmWBAT1YOv8I3fsXT60KIIMzCzw0ZU3y4TT/
Wew+S33icJZSLdaTBx8TGs84yteDsLWHFRQveRGJczy2b6nDIP/RDldd5kzDFCZy
LcNVHYn6xkjZPFeWuoLA8Zk8w7alytzJGu1dipeCjW5xHlZMUNtTs4m0cZg3haBY
ZfYnTw004ZNizY9ZwEeAgk3A5oNiAVNBLftLWKYNXW9t2TGnfFo0sQKQgtM+SZz8
uQGYM5Ep2fiZV98E7kjSwsdYchmnuGACfLi1HfOFG3RgXKCjQtlMpaoA49YfFcnX
mdE4bFjBvxemrGujPbhxE32daNKyhhPMeAdyBbd0/LSKJlVWGJ31ohU1yr6U3sLs
2A5DORnOLEyxWFkcYaMTE8Kq9wyjvUayKf2MlsofhBu6YFGCNt1awVnme+7t7XHR
hluRaUJaW2Mgbdo+RlGL6bQyrKbxyBhYwWT8rVtP4uodVd+yfNB1RtLuEKJvQPl7
P56qW5zcXnx9YXe1KwKKhVHc6LbdUj67gTK+Aa55seOYV2fHhqcPloLp81B9cFdT
YMnkZS2d482aF99bnGvQ0SHPUDeDB0ze2sufDUi2IAAXkSrcOGtEjXDRLt4kORo/
NkIDGHS9HS05kLtTiol0bTcNoeCq8TMZBtJf26Nv7bZNmIxB9jPl3q7PHQwyIbRT
dOrcPGkZykQRMtF8JWwCyeVDXyGB1PG07GF9/crNHxUZCWs+WEMY8TUcWRVtFI6Q
036W2VeZsmdHr66BnyY89EHkpMFQQ4kvTmVVb7aXAw9lOI7PHYFf6ZUVcM54whkp
I+RO+xCinUZDuyMGUvJtGzvxbtBMXMtntW2PYJfrXaBxecdDFpV+QQLL1SP+t4NK
5Kt29bGd9B8kwhK6uB7GDYhv2DpL5wms5U3JlCa1HcWBoKshDIX47JXlBf98oOu6
sXjs1iuzaolvkfICtDdA+a6TUN87qEVxu6IgynyFldq9w22RI1o8NFdVivz25lbO
TbCxtBZRs7445ygzQPgnlzesfM/L3ACyNH4pKnho4vLgrAy6ncQOPBDbLY81LA9J
GvnB3065m2EYyljLOzYZG0d3RngAFvS98HH14AUR7QdOgDxqFP4B2dOW6FKLfHYp
zSwHHrLEzKFYfHPLdD/KAsQs+lrjyBVtSbBxnot5S5U2D54eaql89Aq67khV1VdW
5blMnllAC18rKnRoKVW2lnFrQwDU2INYZtGdHujaczm3z3oFxmlPxNdWlq4lpT5Z
EnTBYHrXyv4bUaJHkBWTBofh8n0I+IUA3LdNM/kugoEJZgUIaxhnlCWh0N8skDNA
sLdHb6WJ5gO91CXwsTV42EnHERGcifvWyptXKjXTBwhhaPm6Pbf0f0cKgC3bY8dJ
l8WEoECBvLT1gVBh+v+ilVbAHWxuRD9YFo28JlOmg4JMvt0cmPY4Nci/6cxfgmxW
sJ5xw6JKKfZxYv/9MonJdhajXB0+jmWjBOHHp6BaL7nOkAX39c/x8zKD2qxElCHu
wK6sW2strmAdUA12vjmyhM3m66Q7Puj5ghvLCBZreCyL1a8Mepa0R76cFQQcrZ01
lwHm37Adptj8v/s/axOxif6Ub1IzgA71Z8cAVPEJTM2eSK0NHnDTDedjKjziz8p1
9kRpLd/5g8MgmZEuCjKa+yd3b0mSKQmU/ulvAlVIhDosbEzweyWS4rJz6rIX1w06
73fMX7vvcwyGe/c12QR1TZJaibuYWcRnoB16gI5XAFDd9FhCCJzBxlA+f4p+ZgE6
pJMWlfYf5i+PP+u8d3/69FzYhjV9NMLXHV2fhmMwsuhVLL+W/PhLSnqkix/ZXQ2H
tHcJI8J+91eq0ZMYuRU/2byLhhhLP2eTlG4JGKsyyDfzcKCNNk9W5y0mQ7Ky1lNE
hIbOA2rOH0vDlx3tGClLSO8le1/tqx0gTrMq73w4iyn7vGZuylK98zSGN2jfh+sJ
2S8PheXD7NiU6AZDQ2p9hFN1Ka7nUZTKVWzjXUSPEuzPeU9ulk/Dt0WxznV8KiJw
WQ/SC60ygNyen9thGIehC8vn+/SgXts0fVMq9c5ogiFXqn5cBHvOJEwxN1XymZTK
R+zA0iYyAxk0f+bsON1wB6WQd7YtKf/vya5Hlq0l8lze1GynyGNsFs5Qv3bk7zjv
oGtShNAWJSJ+G9Rde5Nrl8pjtVRvDb9Zw2onrbGoF/JRKzlkVo8AtJV+QnskJyGW
5MIENPIM2E2TdFC2nyaenMyYFVBPPYlYmS7Sw10ECnQ6qtMjWowbvXVzcwqAhz6v
4EihuEhJl36idXLn5qY45Y7Qb2nB20MqeGFjOZEPHVF/ZoKMBbirxKFkROSNEhGC
MrJeqqsNd7doasdxulrTOsCu4iCDEKAm2nJT/bHJrI4lNAzBycJz4+THnXe3n011
sbWwGqBY2TUG+iZp3cWUoKAudGj4JG0yOCTeS0ssAslgZUE/mGmA/206T2/YYgxN
Lx2ecGUR3dM0CBK47mBQwBsBrgovSfbixaHcBK2/79qncWoWo2xZzncYmnGVd96A
0jN3fYWEIL7Q/t760J6XyMlMnrA42gCz9k6HHoFqka63HXI3GDuG0BP0fxczOC9g
aZqDAjrljyMDZu35C4bLgU1A6QROUrTs/gHswSNc6cCOGYUm7XHFzKAXGqZen7nu
sqNuGHjmuPigGqSy/MtItwx5Cos0ipw15WVlG6+VHvswR2X7i2cqh0jJG9NNsB74
Ts6o/MgnA+/uSCjg/HSFWQZw0Xa1Cuw1o9VMeD3+HYEPcDLsQ+BMcwSQdRYLbPRp
8YzlC/baJKneDW7Keb5xMX6sQiqfztTiQ97oy6t6YGawk616HZ6SfwVAgO45tYyd
3xLLGRqOZSQ1Xky4e6wEEYqt18X/kk3R8zl1uGyIqY+jOj4aIJNzqKOiIYdnPHYj
jKUm0nBnuzVBHkGipe6TUhfpOagvFt+K6y5VO5jw4RgV9J7+4s0Prr7mjLCKVKC6
kwuNec9S9NySfqdtI7TEPe/yIbVTPgYOSjT062Mp2sVEnHeA1+SrTwEX+kUkQWwI
x4mABbhAuUwkAlTOotPIePis0bwkPKaDR+0wLG2UJd1hHurwB4EZ9YiJb20clJCa
83mLXMRsWHbm7jW+uB1vOF0I42TFI4bxMcv+gN/52BWiYpNum3boyPP+9ECEqpne
7ly/bKwT76rWky13xIwg9gHYj6ExScO9QvYYg78UeDsK79pBj5R2Yb0ESkq5hAnV
hFPlmXEdGYB5iPz5lvSALQF1//+tUru81M0L9O6P8gls/5LBv/oE2uiEfFfhClz5
GSlc4S67FufIxb1kq7zAsEByyE5RXm6Z6GZSnmiv++96T/IMQQpCTW9kmCfvO/UA
OW4+jcvpj5+ihQk+uubfxpVyn3crPZc7tHHSXuAR1nwgt8sWDdobt4GmChIU93mT
2PG/dJHcanuBZMTQhdjC7TjyynVyZ2ejNHGpavcQlsHL3d7lvAL6gbvgupIJj9D5
dRDw9thjjvTqGxf95/eiTT4zAll3N28T8DWNaOJixzPSQxxXTqKk88ooLObkN6uW
veIP6LukvwjjNsHM9zMddxLhvj00peAm9yjQ8Yfvcqz84P0csgLP5IwDP7aDxWZ2
IQMyOgIE+uUtL22Ek/0newu3QYr4DGdXAd3T+ARR8fTUTP3gH9XXmj38geFDBRuR
We23U51LUVZsGhBhDdfw7miujPzJrqI2Dhee1tzML0eLg75PD/fgqh+Ss9QjgAH4
3ncyS/K8rYplkPc/kBYM3auy0ZEdvwgMOrsrK18HRMkvsKJumzf8OkdUGBgAhSTU
TP13wvbhHCEyifeie9Zqi8+Xne8FcSHKso/AkH4E7Bc=
`protect END_PROTECTED
