`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JVzyv/YkaH7YQoW4YtFtup5hbNhex0x5d+QmZyQOVATYsoWEmBOn0j4nKjYa2Ar4
xNjTpRirizaXczkbYZBD8JqTNOsb/udxdCTYKuA7HWVqo7yrthlUYcvRs8jWwITl
erXOZz26fQ2rWhyHICutGhNS+A0fkkAjV40AAqKDTcMmcrdUZoXZazEqBd+HcIPf
R1321VqrV5upQkoBmCYrg4yGXPVAm6LkuJO4Mpia+EwcruU5lzg5ysawag6FWcg9
KqW5gzQZRcaC6BEvqGPa0z3bysKDdj4hLJi8M3F5BwDM+62ALKwNOnTqeczTPKRM
SmqV0VpUEvQNPjL8ZQZEVbLgi6/F6zXK+AyQ6xRarcOK0mFCGKrwSA6h93t8Cvtn
Zad+6GZpH7Buzf22Gyse8jl3+532PYW4tBng34F5MFYylfFJQ/RiUkHlmcIAuv8J
1skvc8HBiXOjAczVMqmA8rkiBMwDYJLEWxYcALMi9YnHCC4SSQZhlZX6wdeDJSAx
WhKR/uY0NmfE3wWlvKb/x28w5WS6JdYH1cYJxZ1yjhv1iHAW56Uv7AAL2D0EbJ5o
EjA1AZr4iWGN3IAnAO2f4JVbdh+3z7hLMtjjIRjv64Ow8/J1jG4M6fcjDow62QAh
9uW2htWj5YCxfmGEzYyxtw+IdDMhtFtxjRjwOI86E6J5EGiFH5fZgEGXRvJPkNCc
qBEsfrmsEWbwAHRrmdA22dMyAtkN6LZktRM+EhP9BiWqOgc0B8J6083HXKxnp1/h
DavTvd/9Lb2n2OXBSy5a8Dijbb9PeIwMwSOMEqbcjb+C1dSGChzlp1Zya58EehY/
hnC6oAooSr/yx8oS8/1enix3++FWjMjHLndwhMwCUOJTKYjTOD7lRLPWCHvhOYub
IRtz6ePDbDAw5A5SVJI7iFgpv0G6TmML3e3Ong6G5Gd4MvJrdTV7XIxaJRjC/dZ9
ut8OXy80xJijP5vklK10y9OFljLZakwsXJW9B8w/ImvVtXQD8TbeNyVE1Rfrmq4L
r19HR5U/ucojm9ORf7PSP2+CgS6rhbdEySB0pXnBf/VjJL3wwD0cBGAO5TeuvYxG
VFjytz5aYztwktcxyRWus/Az7gopIgX9bw5APyOheFt/t9vBJBj5csIwst1yx9LL
PdQ9WNTItbw0Ijn2N21W1udxP27ciclJ0FotWQskCWOvAr4au76ynLwLXl1qad9X
nrQuHQwufcKoGIX9vUkLZwweeTCDMeW/TbyYZYy3JS4EI3KmMBiEnazIpTsWAQHf
NartSRFLKBKSOvcqbk1H2KrquczskyWDWULLFp7QYBopbS0xjJoNKj5rwz+/bvea
0vlH7k10tcQgjGd8KyVLqnCm8LrsVvSfNfIN9Pn9J5GHEyIgAh4MbAgC/aRyVZ+m
YDiGf9deV4XXNA0TAs7P9Xz1obROj/mqK1+ttVFjJWgzJDdBgCNHnG7CSS0GppDt
ahKUKfjlDU4BBlYjmeHueRT4sZcNugOcaFXWSavQHwBeGKu54Qz94xiZ8Var/KwK
fE64q1ChzSra0vAwcXjVGwoyuc/qw0h+EOL7dFjjabqSNfMiERQJUqj1RJ7rXCu5
xOHyhJdIB5w0XizRcQn6MrM7m/VC0B6Or1XUNM8mYjxFtzhBqzImR6R/xyM8a91S
r/P2Hu1TtfhpA6WSqAjPlf0pefTRCYtshy9a5jG4ofoVbwMryTNNMAvNotV0RQxP
buT8f+FBG60OHmUijQWirTEH1jfhz1WVs6E9QAuA7GgYKvYqice6uHK2GPZtZtEa
0XCDprjwIrSPebmCg5OQAHW1ZCAKAuIZ6qdUoyMdNQ5sWuAiBPk0bisy+51nGfU4
4i8piG3bEAOtSBQwLSQhvF5/9FGdboZG8PLPcykjI8hUdIElKLaR8KWl0/nsMeI0
iBg53x0aPGKWEG/VZMD1XFdatuKzJVucPYFIgZC76B1JZ9NIL4zoBPYVMiyqYRa8
imRzymnzBfEIjv0A3xGcnHMACf28VL2Sr9zUWVOnf97iBHd3KKXXZVKZ+/Atcsi3
kgGzQ09EdTWp54avaUDy1C86+HKoJVGX0a5SiBXiFO2mCVtG4uCM/7M91bnTQOmT
twrjIIuM6eMvgf6gEfPfoUr3DcQZ1/+RcBt/8UpTyJpR3msOlOKyGyMabsDBf+mg
RDcRvQ2s8hYJCKfWNRdXfK18x7ijcgV5FTddF1GEDJLQ9omQvckTWN0uyWkwU+Hm
P2TiTCiRMBybYl8PHsFFnCZ2YkzneF39UMhN1WooizBndsLuazjj5TmkPmf1XRG0
GhzNYXH2qYLbzxs5G5NkXEmFyKXCQApWUqcpSOAU6klliObOVfpmnkKjZV/fhx9C
NwbQv00w4q2813l5Md+cg92uEo1H5rgUWBqsagd44TQvO2zm20QfKNCMa8dJvqkI
IH2gY1Uxjit2PJZZ7bomCRRwpZ23h1BJM3ksiQzu5k8WQoyueqHV0Cgx2ZLUQGRY
F3WaCAKEfqQb1sz5SwOHyueTKOk1a76WZ+Bv14x3gMUb8Hy7YQ7299zalflwHIDM
0OUKp9fU1yurw0/189M/0e1++FYGCoBKDHXmlUbtb1nN1k7Fb+susL2bwjyoi/gH
xFecqMnacxg8jNqVTGh+ZQLIW7gxjOcBrTbI8yvHWLyjTBP7ZRssYcdd8Dfg33OG
ZNzI6Ag1i+p0ag3QEq4wbmfh6xoKYXTxbd56gMYnWDGKXAJ0B4sDrpdUnUgkAGky
WfG5EJ2lG0cFjrZjWO63cppQhTrRN0gBN/hPVVptcm0wbdZaWvA0ah5/0ACFsO5B
OVj/vXHCC/uXI56QXG9dN0U2bN7tWmFnnYWu2NkU17146xn6mhUUTrlG1rijs5BT
4xzfcdvlWtmnTdDkcgOCKF3LX4emsdJYCMeDINQciWNLJxVl825uv94Pxd+uGxTL
E95nweVr04R7MbnAoMm/MaaBjTBK50LC7Z5w6Gsz1p4RzttJufrLcTcHLLojMc9F
Q4QvAoY7WYn2b/nWVRFZmezZ2WlWJnyGSOlqpkZoJWO4IONklJtBT1c1k2JBNMwV
uOunYk7sZnkY8VtbQFzz178nm+qyzi+YGBq8Dc+ZTghZNzq1Paj9oO7jrrY5FuVa
cxwvdByogk2MHQbFhAdaiQlabieYCWOfkhLuDXovI8qaY+Eh+Gfuej1ELnHl61d/
aUXDGsvKLviFy8xkXA3H1Xv2m6sZR1wlW9LJkA0VYAIucoOz3+aslRxmN0uasoM6
QYstQPTVdC1MZ1mny59EIjqq062sl3WG0TNkxm6ol95vTXUxAkDaTxgjtWkbXWLQ
ok8KM2K+A63Db8wwiWhqTRD0xq4qcxeFgMLo3/rcW5gXrzhvx+8GFpxRi1s5UYCh
6jKEu4wkKNCIdfMYlA0CPviNd0rz82/xfdl3ZDE1ddJj/8IZnawi9WEAlzMwgmaI
hqWcVowHoFcKMR5Fa4eCV5SaO5x2y9GChI4i/BkNjdw=
`protect END_PROTECTED
