`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XUHdufrsfJiLALcfkUaSvhgYd39Htx375Ay7X80JOZZtLvWaWc6+4/WrIQpICrHt
3Hm5T9D87ubRjj1mI1++52Yq/Utgtzh5fJNpmclWopJ5+3jVsOhoUcdJLOFAASfS
OIOr/2+1iKGjHiBVsIcXmxarL2eaLoFjrhefK11XWZGU4aTLzUfVE0TU6EPwjEI/
aWoS1/966fYRLjfN7mNi8644RV1XDtDi8fQzW3sxcfeAXgC7j1nYLh08yydq0Dmn
ycQzH5ot8w4hCelZ9Xa/qgVoeKt2t/KotUDOme25UayT6PvJH6aW3/HmMKJmChV4
1YZKDNai+draaqRpMPgn3AdZJHfXMF1hlvIGd0QPHWqG3V2hVdpj7O8CbiuIgHuE
Kcq5qHjevD8aal8IL0+gE3LCvl6INhSXluDlI4CFhYdsdaW69Hg6XG5U7NvRD7hw
7Aeuy3E+p16nXchxBJF2+Ro2oTgUnj7mFxkVoNdZGMQACK1eUaFRgKl+4Q2XRxXZ
lhD2emsKn4F3/ATahP9CFBwj7bgBs9sPpMEehl1wDtT8971mZRDqDLTBgd61eBIH
aWG0irkNVcFJBRSY5EvBbRtLkh5HeWDR9MqDwLFZfAnpSEHu2xIDlp6xrEuOVcAW
eQdgSaiCspLYOoE/mamH4aDf+UsmnyyJhEZizRq4oDLWTvb5+F59xDCn6f27IBqI
HQQw34wveB18tg5EGpXZW7YcLNElUfxYQNYSiaU1Sfq+X0xkXSKPFQThZGyRY9s3
bhbubbaelS3DZ8eOGjM3w2de8iXLkJFWBXmczknBQEpjn020fQkt9glxpzUkmKJD
Y5LG3zMMszmC7AKD5msktmDzC1zS/icF7Zm4RLh5TirqQLXUhML/Qumnf5uyOcXt
3+4kABDzDgCmeHYUlD1cS0K6+QlP/PkNmSgXCkuRfa0tIu6qXaAJNOIGlp7xfC7z
y9unLwwxvve15f53WTGZGs7mDjqK3tDpT/oF2ClSQA8GTZwHBCl9R/ThPeZJ1CCF
iB/DVTAMmcwXD9e1+avgminhxUjdz30DcJzBXHsEvzaA6sSiHBjtQCVd7sFHwL7/
yl6z4kyVOfazkBTO+Rxmy/wNibqQAyGBRkjA2x6jjVaYppQybtCc4XOtDt5Hc5O/
GiUUDOZIjVSO2FAB/QMfu1IbGGtax0MNZTsNspo8EMYPU2QoVef0LWUzV6P4pp4G
DEUbmE9tgkjk+fabv31oKsnWAIk/Lf1r0InyJTYaCTx6d5dk7luWZIt8+iYiTmu2
6KwG6Q0dE+Ywapat9/Fflm759WK6eX4BegXMN95lRo3wpFJESxRcfggBDgSRRgx2
saSjh92EOm3gCmVeqCfB0Gdi/8tXwm87/JCP2+UUityT17A8TJCUDucUXG7EDbrU
ZejJ+oIE9/oLsA5c0fOk1q7vyZsnOJe1QWa7NLbMwjVS/Sxw+exX5GHgHLpTdrCy
SKXugXZyotK9ZsM5IxD32JcjkaPzNJgzL55XJd3joiFjzB1fB34cDcG3JInsdIsg
oztlUwkhBsyNPSMsrbz+ab1/jQdPBiG8/kMeU8EyXKK0h5k3y5hce/yRtn9fnjLD
UaTWnw2pizmuogTPG5Kl5wC+GVuKi9B9fSpr8aAcbp4SoRv2xyB3YpVHaDhNUnaT
hn06dmxPxX2re/Rx+xK1w5Y7lyNHAzdcP7NOjwmSjrk3AeP5gdFJoz7zA08oAKA2
ZB9k0iB+o77SmfhQSg3MgUW8roofJMVGjoGrJiwXYllVzvvitLCsonSukUB6G0qE
LXhJAJL8WXSjcaDQmGy4X8xhJUOcwSfMivFwGmCH5T0TgzDWjGqFlRd+Hjg6gdrE
8uco3gI/msruChGHDtcgcvexo8zlzESOj3uPPUeRgzMbFzlCY5146RN59R/waWAO
aZeTkYyG5AKVJBC+YoFUkPpk04hEpy3/aqDxm+sXxjbSHAIXsgCNM4u9M/wzZnvJ
QmD8+n39ikP2RX9D6iVlM2KRIH9x4V2fSJrdXMU589QGXixwDLIWKBpPKMThCegO
kfRC3rYyIktHpLeTzW4uL29DspOExH5GKGV7tlozPOarmSNIe4K1XJuEEwHFwj2B
qs3OFTr7WUkP01+JvBhMeQiN0WGNUPT6NbgdrsbsQtVzZLts5ZePkXxeczmA2amu
qe+2oVHt0QcPeBFIVq8Z89RPqX8wWS8bANJWyQ/5WbzLuWm/or/84Zibj/F6SG/0
2xlBGfZnJ4Y+0ZKNmrzqM7LvLx2pxvam8hv3GA7UBZMukFJvLTa25rY0lfES5NVB
cZLGVziN1RFZD8hwf58YzFfah8m3EGfR7Hc5G7aJWk7+tOIrYN/ahRo8ntbC1sh2
hyBbky7lDSzMquWVf+vC+thlZKWbHJUUKgiAe9kJAVGiJJzanc2ruA5SPVh5orif
uswdV8POsVSnET+22ejVLV5pNsWLaEo85tW9l8iJflInrptOfGHz6SUUUXiDI/sw
37T/4OW0F/d3DEcfNAa4szn8enwK3DyMcGHR85INzoJYP4s2/EzgVOphxtfS9jXC
FQbfrWYQtjaQbCOYVGbpPbURbgHfvEflk9ryQHDp2u/dmbImEIYGAMxT1Hf487jK
H2mYlwU4ZObcXbdn2f4uYJKxt2C9uFXCDDCVF2e8toU/LAnw6fVgd9aZDWscZEOV
JJcQNjXTgtb1Gk15WCnXaWpHCfsAs2E3M0q3g9y3U8Ntoe2J6FUNoRiAjXD33eUx
kMS4usRXYbSvlL42og8hq2aXwhgPBkx1z3LnJB9syW8huoOWuBqN0U+g5Tl7c4f9
Hhngu0FHtrYOf6AEU1N4FJK/U4/h2QVyNGTafppobR/8O0TDsocsF//fuLRiL3Ij
SBTDXSPmRYKjoWaCfpwn0wPz2xukPPplh6PQNss1JcOCWuRMaOy/EHiqhk6vIPm+
sFNTAYhWy8QyztDrlINi4xWx0MJiAHiGdPiOyA4cFcfBsr09wIKbJJOZgWGw3wuG
24w+Vb0EDR5j4nXn5ufdyth97e+BLTadk8npIki/BqCz4KxHyy9mUu+1Lni0907n
tYZFxs+omw11t1Mgah0j3VA8pu8Sur4w6ejqVWTDzCZaEREnw5dUfybaD+cZCkNb
JkDigQDlx7JImCidHC3L3p5TCa4bpD1QMQGsTEAaYxVZwoO35L+qMVA18l+OunBP
PePQSjo+cqpAifwyclrTaXDQjn3dm6tvB5iu0IwXg0B7AzwD00cgnzVKjBejBc97
GXrgi/NHBGa+vTJYvi2RlfwR5Jsz8UQQMRC40PJ6HcWkjqsSj3+4n7AZaoERbEip
2gdt7izjcAR7vnmP5xrvdSxRNCl0F9njkMHPGoBesJ4Pcqz/BlgoqqxB+lAPJSGR
snRBKVj/anllK+G7Hl9x8XoqJbVukg/hAcQMR9tMG7CTzAyh5u/DTD1iUvaYZZzg
IBVz0yS+Ehkp8AHvwFLUx5/scu1rn4e5Li/ywlVaM8M15qYiqsoDdSfhLqC9NpFf
PY0LLVig0E1ZbQbN3R4Mbp8wdR8dYHjVGasqN8iqSjRcb3drKg+qnUERh0y6rSM3
dKzZvUbKDNXvbnfyNHIEJmQTVGcnFcuHHJkmIl6hnsqpD5MhPIDGCtYfRxQ5kvsv
FpZg2+PfSmNlYCw3xZMwTrRN5Yuwt9pBDS4FQ74hZ9olEkCtLXf7LqiLt2mi8yBG
ZFgks3FTJoEm6ty4uu3qS9O5V80zXveYY9/5ihhbyrf4Flca5ZOdl3soPYJqlPzA
3GVt4mpWb+C9nX8EKvr3V+5jDdD8exJsDPwqCtrnm4/KOj32+5aiPMpL+hutLA+z
ByUK3tsEIfX84ifoKxbtkcXlXn+DbjUtJFPaJSyTiyD93HiFDjERcalXuqfECN6g
ybgn561WS9J1MK9gCG8/rY9UFPFgHj+u/tB2D5R+WxOehH5dQh4RwFOsPpKewJ/C
eg6f8qBB7J/rNe9ZHfVmwnUaMTZgpL4WQYQHeCtDINWY7UaChd1sj3uXQOSe567W
+O4wPCjnhJnddKaQtxPkwXAP8iLqkc5mR17JAh8iwBrjqtbZMoE1pymjvzStknu1
iHfSXngjSr5DxnulXAJ8mmOv9oWY1y5IuZwYusCFv9nGNHkw3tgQC7wpdMVepFKZ
H/herCWLQOFmKNqGmSUNQ79JRWkD1nE7se743BkINzfGpUqiOtXeMjbWmE9cbLPz
BasIeaGe7cjHR3hgSz0zEgf5esOCOU5t2DH6E8sfd3dYnbrmY5TwrjM01cngG5I3
naiCiL822k5e6DUAFNETqECKAD8tH2glUF3NQru2lkkcLVDQ8hfu3X7fd4/7lF5Q
eK8YnQsn/lj4bM/XOqggMPN4IvmylbIavEwgt5n7oJcryaUwao6qjMndvxpDvyl8
tIZ76CiNJi29afYxj8tbdhRjClXYWxy4DhpkaXsktVqIfwrg5GabnqVXfHsCIe4L
oGV0CvNSn5L/XstKn2CEnKyDSA0qIfiDuhyWMrGwnKo7BX2YWwpIVFc/cdvKLsGW
tH+ehI7KQoYgdVg8XDOokQ+9Ukq+JqwwTnBQXckayxFbvrye0cY7WPawhm6yPunD
EZLLw4hIwucl3D5gUJIn3NVjMvNlzIGVmvA23CWf7DStTXk0ZLu32QLUuEEAggbu
ucU2yiEtB4h8WDOoUqkBYI8svojQijBbHEdNfya+UrC9uL3AGlLU60k6haMGHTr/
Hz9eUABEN6D6HXdB2WoeaEtqikMtfGQGrP8fKBlAZAzjsSDpI2Kr0Tl2Pkqlnq/M
iAQZrfw8azS48Mg/4gZpwZPk1l3kbtJwpGCUOzenxNPNRDOcFj0vfA4sNwUY1B2D
YI2Ctp7f4oCVOatmXIKRIeyYImyT3nFrFtWdnqiE4gqmKWlGsoc3DIlZdFZ0Cn96
OiSx7SBIR4dTOU3Edo3mPw/X+JZC+WbBQxark66xgHKVtqGWUjHX/DhxFuOIXORG
uE0feNMgMWUGEBqcUCdb/HbvSx6qv3wjopTvVFwMZiKA8By5/wo/pqZN2PraqS10
5RtEfPmulLk498ZpIOINza61HD4eQ4dE5lF36VWmAebuwc11pHHjjT8eSMQiMJ4D
Xd0rfZ2VmdRfGT3Setf7AMaAHdWIypJFYn3IGd+AluJQJYFMho19sBXVMbMJIWRG
kHwAjpRpz7sWt11wk3TTPNQweDL2NFFg3hYVG0nI6IgCep8yhV5iA5r3yqzqEAr0
rEKM4WISRt6lamizf9wQDMjklJtj4Oeh7YeCyLK5gaYEREB15a+lHY/v2+t8Lxuk
z790Db8EtNv9w/hLTGoQrfC4uoCb/lyQ3wRnAuGGkMahR+LAaFxWT9VI8zCDu17O
3lVYgc5STfkpTqE/YuEFHSXtwsC6cDKhrmmcAL8c9P8mM64q7b8ZOn/EGuQ7FYCl
SagkrM2ahwbBe/mHMizZDARnXY/4xOy9J8Ejb+A9u5xZhBAI+hhgbpVU/rdU9PdI
tSvlHBk+BwoPDeNNrJWx5Iv4XUMrEQyeEDg8o+URNENJb6R0Hm7pYDIVFiX3eAnF
0AIQluuAxe8pOKGcELSOpKy0BHNABhg9iBGISEyKBVzckLfNXpcOFAAybPinza85
qSu2mb4rV+Ef+7Ql7PbEju5nwcB4UGyyhOTvNchtiAnrgAvbjSH+YlKEVfTn4QNg
m5IaUZC/NeaOlKjk1ll4oqUMSzMtIFZFkBR6SBn9ju/aXJH3GhLFInRreNAfm0Fp
SMB1I2zBbGe/Q8eN5gN7bAzkGkHu7uqOwpeC86dDxKsnNMSUedjrq+9T/M+q/O9L
MUKU6ZW6LZVh0pwAPrkWH39Pt/BdXzW0DPebYEZ2kkwS95yBcoyVpkBecdQLSHVz
6oRvxUcvDfG7IIfsXWeDLEm4rIpJT75tNFMxsmDSZG5KYbmD4kwwgYPsr5ixqgUB
EH2zEn4CMn33UYX8/+uir+ym95lseXnsKn08DDS6WFmB1jlboM2CAB2k1Pe6nboa
/ikQgP1aZdmNnHBCzhrUqQI1lYAcfLw/6hrPzH01B6WCImLmJ4f/3D09nLIWeMvb
lBmUXkK/m7JXO8ZayCmg+tNAsuIjyS7vO8LeaTjXuThgJpfjypBPuwcGJiR/5pSZ
5ThPp2QEVuCD6UpSF2KU+Kp0CVODJXrXogOx8UPcOnJ4d8g4c2kazPxyM0TEx9uO
98WjmISmQcdImkYZq4B810/Dah9v4TJDt+Erv3EXQuz+Oy+HRD8LjIXM9/5jTMbQ
RqgHIMuMLAhYywN5f9HxENMll3Gx7kfYsdeLdyQMlCnOAhj0MleaxT3UePLemW+P
EzGyWP2/IaHwbu9j8t2GudKyUIoGux8/dB4gm3aiuxNHYRSBd9O06M8FEfru34GQ
Rr8E2hi1f/w/f/f5HbLWkWvW8lIiQORW4XR8sq5V4zdiVWz7SizB2Dgr1Hyx8G47
9Eb4I77GeBeyMJfjxT46YgSpgr9nb9Tp10jCi+t/rBGQw2KAYnBD2d/QRiC7lkI6
fRCyhWx/M5B8TUFRlkldiltOZGwjDWfp0HDYKJShYVUuLUrEX4iXdsgAfV+CqPML
Pye51dumhB0jlLmtVpNbXujZIObdB58vsJkrenTidasWeu42ybWU9kvN+DGu7wAZ
aFEq4txPTt4mOlrnG85sR2xmVLOed0wWDPp1yfZFKlgRSIeqhi5ZrouX0fMwDA6u
sq2Yjxd4wJxQt/KjymwgTDHkTbpsoN4zkWAl0CLa2/9R5PeQkVUdwaXFnsVxcLo6
cPY3YSgPANSk2CJBG5NKudLyw9y8Olrrq/X7Kz1P0qYu99Vn6a+WnlQNkrLns6bS
gmKJztGw/NovLC00m1HSVM2W2ntmci9HIP0HZbhXyTue9R9kE32IfwqdBYdqGXB9
NNDmvhIYvMCf+lwvNsNu199jhucUJ5t3VqcH52k//F3cHlDKQEPB9pdZ0ujToxnx
ZRECjmazRjDkvZ1IiTJZKpcbXO1y7cVjAXwIuUtu4i9FNBan1t4pPDDaqTiEjlod
Tqmhhobz98b2DbbmfOG79bkJV6WWUlG4M5GL1ri71slIuTIUPSbFPGJGbVPXyNLq
Hk8tSV+o57O/pl/FQBond52mpaapER5wOZy6lYNHvnEaLPOpDTViuLZSSGySL1Sm
imohXChgNBZNLVPnZRI8ulcae0qDLLGWg1mVryY5QPgwqgIDmksk672T5xuBhV+5
NcO1q/rfcZzNmsR6b5mAr3d+7aqMGTvYAOgpGdpkqwSPfzL9KoTSCkOzs0aHOJve
Bikxoc5aAFTqT6UwgEXuMGONbz0dKUiID4lQLpXMsTUfL4caCZOKVXnh5D87/Jhg
jYy+Scultzbfm1EAZBxZ1MP+o8lXR08ebHZnlG1ZXH1O9Rxh3I2xix/O7TmLtQlV
ilCYN8j6rZTjc9lJvKmmVB4Uk2IFb6QSDclj7bCOdKIB3yKXABF/pEc3l0Rz9xcr
hsMP+SfublWnAJzyHQ1ecsoOvEefKmFtKD9cEzMffPuanN7vFJyQP44lLECnACWI
AiUxa6kTMhgKdA/VEvUNa/q86+9QwFztp9ae4CwwTC7xuUW1vVXq3zW4brxTXUF/
ZwovvTPbHfVEbIeEvb2cRxgyn6FAyJ1luI1UlQY8ZBhqDE1IwrOeg9qvedK8THv8
piQfWwl487TZK9u/Rcnqp1RkxBk7Dvz74+H8jAFAuxe7Ba1UyaqGc7syWLLLXBQc
sTrmmOhx5hzIf+RWhkXQGTk99iT/Mn/DYTeO58ftTbX8VZs/yq+seSPGkkcuTePM
qfS0Wv7vX5RTsaLiagueDXYiBzaPFu2plapmANN8Ux3o5+UxilWv+s4dGys/cVH3
EbdUa0rUUpGj42sGc5STsd3mWUVnEX+nOcBicR5tHbIiiAfi12KdZlmoWOkCXxYF
6K02hNrvNoRhrZYkL0oqU1v0OhdLQvZ1fzgPK4KpDfvCGAe/rXc/7UXwOPm9s5da
WJ5as8ykGaubAK/x7dhPICU3pcTOa7skQj+TKSwjh6uurQzcsZblRUByp/DdhEGV
0IiTvQaq1xKIGQYRopFdomESQ2iDMexyZyG/gaYrL/90ynC3fmoQhO5QUi+UEOsW
a++kC9oqrT049/JymkS3LIgmBNAkOimorJ+sBqtuZj2z8hcztDcT+NOHt4MSCGAL
3agSNKfauRgJsNMcnG3xlGZrHFUVOWwHVdE7XXAFIwu5Puqj7KjrscbssAVkUjyE
uQUOWp5xXyAn8/o8UuaFoNWA6PwZJRWZ5tvryI1jghwCwFjPfM5PogGLshxy0QGj
L0UTy9aGzRttF/Szy9wVjw95DlZ8HEUJuhTqpl09oBAw3FOOkukfpB8hGuhg6XhC
11Mw2bs8BMNdqnPO+8EJ291Kuu0pPg1zMOiTCA/m2qE/u5Z3suKkiEcY4rBVmLhn
pn4UPiu/Qwaiq+ZeZSGc4/JQ5jlUFsy2qesrC16f1rNlZ8WCS623+uh1VLT6Ws+n
mbrX9M5sNji7NZITiv/0vap/VmxA7FHQkTFtWPGVYJ3GcBQN7iX8vwyFnRKvZmAY
WZsTxFYBWZma6NFsUDkWjBNT9kxCS3cHwld5ZAnPSWjiJ+10pBob44FKEZoPicuS
ddWoiZFMW0XsnlDvtzqN9UteoWqZaHC8P+YaVR8v2E6ZYcB/9Cyl6SzFYwtRq47z
czVJbOtilZKRC/2PF0wYexqFoGAHRKdKmNBfghjBjmm5ejWTHraPkZ1mj9J9oM2J
wvI3PZhDg4sjt6vBn1pyBd2a6A9bbwGSF27tP6u8buq+W1lrCUJfV2ZSAhRlO8Bj
1utxoPSiMzbfxAge1MPq2bfex1QmxmoXGUP+KN5EVzJRqFzpVHxm89B7p4KBBKDp
H3DZsevTC1CfXcWt7o2/MnF0diQSKnpL8CnrMz91l+URVFAlGy2rnrXvSK70H7Oh
dakMF8k5Y5QMMgcpNPsSEOQWHpuEW5qTgAVtDWD/+SrHCumQ0jruw7SdKQojQDYo
T3yZDlCi4bc5jG/dOB4irvt2k5DkxrDSEXrd84iPe5yidFgb109zqrltotzeN19b
K/IkzomfMarRH47kWXAVH/4sXzNXVIEZ7h8iIjXc++v6ngelq65a6GhGDPQJhvB8
SdewdkUxLj9JlWa9SAETPss5ceI1P8HGwgXk0R73TwiQiq2k7wbp+EQtCuscEvmU
3UM436nnkw8kfEKy2fjW4CtqQ3HKKhzyn3su6BxmnCXlAHA2KlTWm3HXx9LIsayT
O6ORYNB0RPz9Qn3FM5b+K/RDqR47/r8ukotcgv+kC8wxdbBpr2IgitlqTtxcwopU
0ZloJ6IIeuBMZD1KG3m96Vts95fw7kSanU6EcPPzYBkQIM7FBzgI1sNnetOmwnF4
/UGpDAUS6NSWsBBcofGww4WdERj4bvAlTaBZZhejdNzrBgo0frx7+PPbxNVKON5g
5RSn5Iu1Q29c+4okQNBh03c7Aigsnpo7Cmxe5YkNkJxjHQFtO1Nca+dJlRwzvqAc
n0t1Z8xHQmLE7m1Ylv+LX6oShsVzGE9Dy69CuUPdt0A2wZJaT0msHsJIWADZMWS1
Nace8fJDB/rIic9w1xZPgG1xJ7UY2XB6tbat3klayInAKE/a+13M4b+djPEM9YOE
MYlS7UNqEffsNbyKUU5dSV8UVIsoXtbiOdfwkRs9TuraqRYNibZLHLKvSr0iA2fc
wm+OtnfqzyLXOws600HwzerY3MQaF9jROjRU7mJ+DcoBE7K36/apZ1aMN77b5PZz
sNCHnw5shQWllkqZZG2dbFhzBaSIyP//n/srtmCqbwEWyoCMpfEV2Q84IsIt5tXe
BPbg7zaVAUapNo86P6OHEASYJjakr7coZ3lW6rUAMzfVIa/N5B35BlceA/KAGWoy
4mkNeRxCuPv0rXajkgPVz71/rfE/0T3FbhcIWv3o/mudPwWR2eG/3oFofvM9VWw7
ksWcCgEWIHisP3D55dBJw9IihPeJjsbr+BVCFGVIGcIadAjrZXlD03zOAcw32Yjx
hsB/ZbaHCJApq0XQr6fi402tbCROrekEYIn30Iau/Fyxnss3f5QXTt5xIRg3ES4R
7aMgNzf4XeC50xNAdpKcC3CU+D9KkpjqPNXH5k1rovDHHz+IEhpOKeP/DVT4J2sa
2AiHua6VcfNnHn4sdxANGS2H5IVrE2IlT2y71IF6N8QUyemP+Dr++fb9GlUGEW9K
mBzqjlSCDXPS+wYFFLsApGJ2jgpiUNR6y58ZMh8Y/OWgiMPufsm9SaPC3gbFojXg
FIZwdE9iPNSLbMi72gHqs/v47Db7gtsHWagdyT64qq230hmQnBKkFzC85gCp9QBi
qy3KioQU7Lg1Ba8YFbp+f+6Od7PyYwevyGb/S+Ep/2H2ywc1iVpFOIRymil5fimw
eAtnuVN1/NToMaPyRvXHYRZUKWzuJKm+KX73GGNBpq+bqgeGDb8o/QAxipMIww0+
uTsP+HU3qTdpa6TqnCCD0CcmNNY/VOCGD3ZXoGh3dLIo/qVcVhH7wggBI9zt78ZA
uGvMMaHpwCXoeHLrBJPFjbW2PJWpDmaZWwd/ZejtSb4HLz9uIrmMZCDVkgMg0ar2
noFAgJ6ecCVVT1+/1vVvIrW6cHUdYFExX50vjRSFmmB90umpG20kmPPYmX9GGjpy
t0+SmW8UNLsD+GiRXTysiZ6F0fuC2Y8DvW+mm0JBsbB6ZQL9TDEJW1Jb/8ZmW3pV
Yjfpqf6qFMJkg+SdSzuTQYyP2xv8CloDsvnvqZoJO8HPSC9nDbgj2D2ddmLwM+eI
wXUZyhgwAuilYo+IuSyJIWOuKXVXeodhAzXTv8OJ4h/v3RuRUDDVJh/Im4zDRx26
zrEF1HK4t1iVWFswFRraGjyZkinENU3EkTvi2rvXfS3OgUWmnIjS9AO0CZOpeUjv
VLTSibWdNpdYb1L9X0dXpEc9oBV0n0xYI70ysxiGBYwEzjaMFHnFDcC26WEx8BQi
WGIzJHv4np+UKznkjvSbk9mQHmx4/mbMIeMSzE+tjbzojKa8h2fQ++sOwjVNqx9h
lubDkTP+lM22+Uait0TUCCNBlVINJKIBogO45z6GpDZp6zVaTHat6ysejFfAgjON
GjV5pvsBkBBxIBrfW0saZ80+clHdbpn3TfY55NQOxpIWZ8sf2MwQ4sk9mn7XP7lb
jAUIq0vm5Vh7k0PZHhBn6vAxuZDFh5kPP3ypJluyqYdLLc9ZdpNDnlCUfaFOQ8hD
FROkjVl1+TxJLg3ihoiyiOw9LYRNubzu28PxE6TuWbbkML+W/01KxELtbS4PUsJm
ZT3FVkQNd1rUQaLTSDvSshSDlechNT5oMo9XoQ/1IaW66TkHGZs3HqM4RpnJJjTt
JKWWmfH5bXAwllVBwGfzfSJ5As7UJiYqdWoXTtdLJF/SZTl+j1K8s1WxAyhMJ1Ox
S1KuHWql/cM44cym3lH/MQsyOeb+aL6fRsyi6tmwkYnMXByeMkuQqwcxKfjUOSnK
VUbl0ih4vTr1eGSmFexr3V0N17WsAiBTetaJxBLJjeTQ2rtIgrUIjxLLWdCnwIsC
8fPqraWLNTvnD6wsTpSKjJNoclNjEeaV9cE0roC0iXs3XvBkosWEkxYRWO/45f0L
/3hgcfWXNq8UJ56AGhdGia5exC6o4iMbhuY0mR+B2mGka1X8nzOgzCSbhSaYFyRO
xOMHP4dLzQumqEwRIzZKOBnM9sJffx89GTmS78ZvMwnthAykwQ4aH+twTLxWGWYy
UhxBQyeCDY4eVLvZqt8o6zstpedga+x87nVu2mM+pb2zNfpUzrV64okUq+hPjvOt
YChiEujSHPKXqLvCmkRksEed9bwzXBuG0OQmpuDKsEOmxe0FtCxKLWs6UxAFl3yY
GceNze3Ob/sW1oXz1INraZCxsAl+JXzqji1kcgH2sFS825EzkFCXTiVh8vN5uazD
ocoh4bgAwKLTEmxZ3d6r1CFZWSjAsJL05lVCMANKTWkKh/1O+VwdOjNuYXSpIs9h
h5FAZNuri4B8QiaJl3lDXNCg6E7pgX+CoBd7W5Y6GyQ2BlQaTCQKhRX92TRSPaP/
vyJPN4DsVQzKxMOLO/am0X9ysecz1cY/e6Z+Sekry5kY1E/j2zePUXUQfJ6Hlqt0
ojmRITpozU5aUxZ4kv9Ld0V6kX9G0UCwxO/kPvIt/16ySP43Artvzw39vd5qW7O8
w5OQx/WN3siy4JzOL/06+BqS3AORMW7jgCydFivV/85143CgjJz+UrbQY80/hlH8
cJjRxrS88PCWxGwV5NAQbSD6Hag4v/2nIuConz2ZTRqs309myxIUrjziaIhBE743
PZI13CvadC1FPtH1qTlqUmwyE9/luSsKWCB95gb61lIeAfMJDBBL2uQlm3lrvpbr
ILe9PAsxz6mxLChC5PZ9j7hEgtET0Mv4Megb0k9aZso0WPE1J1eoy1Ae1a3ERmX/
fMsQrk2Xo246ZuQykL6qivv0GXPQK7nxcXBe6HEbO5sov+4vrvsDPlLM86RRihU8
0vdzjXRbHf40lUdbYvWqPrz7Byc+30nvH0rT07fcCH8DRapMpPucMib7SNaxOfub
gPu9FXA66sr6lI7ivdS1hbPoaO6r1iQSPla/Ba/1H8X/MpyCI2vaLCsRlFYu+mG2
x8UUsnOfpcg3QRFPQJF0ELl02qHJQHLPaNWX5m6/taVan5dsy+jWJSM+rFgDO0G9
JRfNxftGQVPD09iln48Yjd3HSlJ8alsbvhIo3FO1mlH8WioJZEux4XpjXM7OEtMN
9Ra4fkmIHkhk/7teEABktl6lSGjBdSzc3aA/pVMXTwlNByXf7uBXvCVnNKKT3+4M
3mC9U67QpUQyr65vTC/1uxFPmGio2bFvo/7h8nWhtPbBWvs4Qt97Fl2CkdwgydJn
81+SMGQedxDnoplbSZAOl7KqvdsdocnMzIbFNmMcs39RnSxr/ODD9GLkOwCgrmgY
xfmHimw/O8ZI/QwurM+dZUzPE80rF4HWF8PvOtuQjeGAd1Ts3H/o673kKlsgjZYO
IN6ntlgOdtHYKHHbVlkxg0uIDh/nVPm+PwJbU/XFFA8VBBvuH7t7cK11HpJBif/K
an6rRepiKRZasszATM+96JecjkersjjNH8s6e1cFpu1oF0RbFYoSCjwu4tSpHX4d
LvfCu3/xSZgEDlo6wFmRRVw5VIVVpWxJtuTv3+5NsmGvIj9ZzkN8pqyU+9hWDthb
OIJK0mA6xbiWG5vwkG3Sot4WybZaStApXbIurnncwVz+/woCCRcC08ST3r9j6rER
PA98zMJMW3E+w0Ai5R/WGk2XZAdibenauGZR8k7NO8EQGcr7DQRSLLyMGGgqJuWx
C82NRmwAat0WCue89kxb6A5VZQnhH3J+fEEe1Uz7lVTIb5cNIT/0FNvXM3Wr//+X
aciwRTjQriglFfujvWrC5uArfklje38TpPP/d8ApS/R7HBRpqP8OTuq4bhf/Rd4T
ZS+gXv0fGBtnnY1DQLcnz3qsfMlp9VaKNvrvp2hpC3uPk1ZWqpkvYFH5pc1kb80y
9N+/W+3HNZwqDYzo28PCmRNObYdpK/EPlxTbMIlQG0cEV0uFNkTb/HCDFoKRt7/6
sa+V7ujECnFxGzM4KTWV/Oc613loJRRARb9FX8Rc428JQpI4hPvYK0R/8uSHxZ6N
i3bVAbx0EczpKOwRTXecW5m8ipyYIf6JDxccs6DrKR2DxSqZBAIIMR0ulIwQhQYp
4P064xsmYZuI3mU3YotkvJRgKZN7+wqmi+LplAby4LRbEiC64HZkydUAp5fZwlHV
VyfYZKr5OVBEs/Lpokl/eYs9jYFH/FrhnNYwgtKTmkv8YmZQyctNAsjkfuhKCDGN
634qc+a/eeF1AFO3aGuQdjW4sHxOB0/GO9MTtXmp9oO7aGmCGRHeO3qdVkZ1ChDm
F3St/FC3I3tuxa1kJ6sl+Pp8S4+mW7CWjn0R4r5oo/nZD6nIKJRflluf49MnJAG7
jtyMCauaeJrz246KCh38BwrR2CaNb33UBfWeRZwKE8HgGA4FXssvTnu1pkjwAA0v
ugBQMAE2rRjp5V0Wm5VGRrku83WbckqxCoq8s8jiEYpFZqOmXYHqY/MvuXydLDei
V2mcjvtjb0KKZMQIMOi7jJ4G/WvYrx12UDkeA8L7TwZoZLthqpVMUHBJU+x7RT8h
iC6qKAoj62FhZIPGtH6W1NbtLj9dRBC7xORS2B1wKOEiewNy0kSkGKPgoZukLmsJ
4JNFw7aLMoYJ8LWrlYQZfoIHDYd4Hf7Ei42yVzaJOa8IEymF1jfeqnuhCEpEq1kf
FisSRhk9xPvdz0tAELdALbdkPP8gXHgFm1Feec7+hDuFpExjZLDg/fUilBL2Nsfb
xmC5785pjgMx1dMUQFCYI3pqKmoZHg/eo1u8F6c+qDuYcGgH1CpHA1M9HallA2Zx
sa355nzRKe0SZ4vhr5JzzOfM4+lCmKChTeC1DvTFPY+raEPLCdQGrLNQxU6Ra02n
jY/svKiFnKMnwi3EUH7XxjN5hMiNvhIlGCVxZtaWPIE67TWHjtQYjxDkJEQ6tFII
udvFkgOcKhkxYxxHahgs2uZcJD/LHraIwqn/BPMfuIJe84W012VjoKkysSHE6yfp
BKSLqq45FeCJt7o9azc+ilKPgU/7dUZ+/0PxWM3zUMXsxWssRSKLstvXohLzTnbu
ieT+Kh3wPmwVv3V5mCaGQOIRRFhJbm5RBWUFVN6OrKadQHw0wPuRy6hg25XVsJCn
qkTN1lD2yR9CVA9jL/KMCjMnd0EEV1ViHYbTyGy2YCGKkcZUhlaxD8zkwHIGEMXj
8fnuOguIidWKeSIlwnHbkfglViz9sWgU51INk8Lx9xa53VD9ontksTkSE4ztPEvM
eyBBvtzsEjm3bp5nH3xtz1M4Cf+nuLvKm7SytpGdVz2nktpI/y+ENExqQIYfcAaZ
bOa+Yvc8eNHq5qiPrpfLPcztZxM/FOpw9w5gjPBKhsmHHfFScuOEJTZKcnhiAMNt
afl4RsWLM0QFP3uJL4Wj6edwQ/xzvsP/lxdokK6QTHP+sX2RidhKGoG++dt0T0XW
GqLHjZs0EH5y+6oQGHastrsFremFAk5tXrzf7vdqrsqOBCv6jS8ea2TzK9KaYXTo
N8uuVKszoorXrgX5G2f52eCR/IrQi4WwT+2PM6vMREOEJpEq+34/kq+8CReXYUz/
wBvN2cFU6LDpdvI3FRZgBSBz3ZtMqGNt74Dc5Jte1iAgblSshK1dFxrjNY7rSsgw
n+FSUOmYigr4ioRsD/EnxJxhb9RaxrGSx1J+Fhb/R2Zx21vVPag1LoEVcyPTfYe+
DZ6hAWQXasUbI+wunIbCmwipAIf0bjIgVmPlL36AwQxzFL2BWc7Fx/cNeS/xZ2VK
1r9+oMVIRboiHP3suOZNfXFc7XZRVnwOz52gSXV3HK1q7cltjTFyLRR7QKHa3LDW
yZUSQPV5wREM0DAtRmGnle/RQjO1JRCRPgzfAQKGyxtZazmoY4xmwU+KHb8R9x6z
YDeyWtZoQbnqew9Y/lJ3vOGhJNwVIlYIe2XZ8xpv4KLtewJ9Tr6dq1NP4m5yw/f6
eXtd1BL//RRe/QJrT0b7JXJv+/KE1qs1wKk4VfX49YiAwf8vSmoT4w0qV4HZYza7
yuJGXG0r2T0lSFDcsS5+kowUlSce03kYkpVmrwm6AoIKUdpW6SLOQ50u9k7IgRa2
Ybjxtwu2AXr0E2N9ntgkOkkhCyv7Jy//o9SeBBkkUvlXM/p5ABqmK6jjfx2Y01It
lFzdd/9hBtQx7NAMV1pynS1483jsxUea5nzNhQeTXmeZ5dah9TrQ3pZ1AjBDoKfY
5RTDvonXNgmrUpgH8SNyGCtsroFVrL9X7W6hPaUwF1fQRpIWqIDqZQqLoahUCrRV
DIVBm5iYqeNeOglNCM/8La//AyYXVcQLOnxEion6EugKpZywyqZQ0ofTF6rw5R/w
A/kD4oDxT965B63aj5pwEi6UMKF+yrBqFy0uLD7dsmeH7VqKCr0BsN1516o91FGo
IvU91j5/UoeX/QZx/QJ6l7GTqk9RcGUoFDSE5rwkMo7qCyGdTu7a49VKoub1l7pl
ApXqNlgJ8P8UiWgJizyYzH5EYTtEvhR6hOe57+vKR0EEslJIZS6t4GbmnEXJPa2I
1Ud+xZlA1dYXA9mYoxWLK3eGkr1ID08dCDlMoJXk+8hEDwC4iYgBI9uwmhO5PmA5
oHq+Y3UOksUjfMmf58Q3Sah7qe1RAoVMZk1qJQfNKG81BfjaYMo39K+zBdGg9y+C
+3dPVuzTIREUbXdOjEdUMFoHrLLQKGTGJzQ2BnZ7oetK4d8964kW56r1cr6b3ljK
Iw8zVxgnXEIeGcByxJxDDO9rCniiFSnYekoqEArod/TSxLVwo9fa1c9P2y87T/Rm
KqRVwG78p1sMvL+/Y9lSLgAFDeF+Xncu8PV7bYTB7Y+1fOfwAGPJ0GGOz148JRh7
3RbW8U1opYlErMJRQvAUDCAAhbHLsl8zAck1yW6kEGyyF1jbcYlEeiKqHgRcHgo+
Lyog7eEaqJuqTpQG4zh6pRyeYFbDVpE/j7FoCoxDgTBE+TJoJeDGsyL63QG0FpAh
mlz0hEd8TK40ZANiPk/SOWLj7nO2gpbPiWpxXG50VaQmYdBpGpHhucvEn8qhAQvZ
uxb793M980aCmbzXTm+n5t1Ht3s4mKnfpB/GexDswmd+P0b8gbZdCS9vV1yPIFvi
0ouuy0HkF+CMuxGvRIHBJA5azcsPKPekzRxl5NwLbBaiBk+KsH1486LfiPIpbXhD
YYdugFxtM6ksdWFgAx23YguaVX1x7NmtmKWWef+dh8bjT13na3rEuv8DU9HRKKBs
1PE9Y1B2BgXSvx9x+hvEc2dhz9mwjDZbVIXQsPn70C2UbeZK3X+sqiFKMXWO0NYs
NRfOXMrsz0PFyFdiC/g0xP4tF74FAb0tOUbjPbqEtlhywadM/Lub0Gzila3swzOn
evT3lM6nfl1nHYfzTboE+AwE8/DLQ/JM+nF/cZy2v3Km4dXHFX3a3Phd5pWMxKbU
hMqRXzYECoc5PhBxsTU2fubseXNRTexphUjWwyH1xHM1oniwR16AYrGHWBYJ1uIX
fqP3fD/jWOro0ffX9xckQcHsyOTRn4HY5mnnQIHc/SgDwEd38+M/48GMfrmEMNck
+LdIpj1Bn2KyoHoRPtSfVHNHPN0lBItd7Q70V0mYKUmSrB2Y85JcyptU0UG13FMB
iiwaKgEK49QiGOq8gtk4AzDwrUAU0aK8V4ALcIgwirEQX47pSmt25XrXCZTVLcr1
3eVCOIlEfZ16JXW58Ge1lRgS8f2U0Qskc8bYaRrldcSmxMwFje6V/B4n0XYP8tGe
1UrrVTICXNoSp6tbbQTNwdnCvC432wiFFhHs2Il7cT/dloSWS3QbSehermbikUPe
d+8vlzDxcoN101vlopIn0+d1qS3LDRVGqy4fcF4XPnoxxafemfxMBw0Ll875z58U
qtUza7oLpMxOaxvJSpnMZRvI0Ppc+DUrj6JFoyfuSiPV5S/q1bohwHDAMPyCy2+4
KtKde2ZpiiuZFSRMBVe3O0dhtZE3jxAkNF5boadGu8Gycn1LTq8Jo7DVueGImyjQ
b7tUIezn7kKu2mjMQHYUsWgKmZgOzH+/YGkfEyOKM2w0QqLjKVLzbfNw51kf3Dml
Vwe5oZlX9tJ4G1jOkxJWyPjrU63Pv5PzgItvGw7hY5swwEuplWM6DIfHHl9Sg6xP
u78G97YjcIfhiGeL0Am/GkE8yXDbeuIVhSb22xLSmWCJP3rK8DV1n1af9kCXf3iN
jtBdclU1XAA1gnpboVZU78lo3+1RzHmF6lyEgstaV/CRSg+JlsN5rloJnyu/M7xn
8mHwaV4Kl0tA9y9Ot9lir4kB6XyAfNTBgpaFyATzOiw1CLcoFhR7vHc/L60QUzWi
dhXlVy0/HLRcGwQhWYr7Q91lak5q/RxlXrSc8bHUWJYKHj00jnpwbZeXd/40isvU
2YfIzEE5dWaqkqIH+i9WC+RXU+Aqg7w1uA++kvQgoWfQd2pXF3bfylNkQXwwyvEy
beaRnzIMyWNTtT+kq2FlRJl6iZK+1yfuHjsMNbwWUFpjzsVcTE3na0C2tzp0RNPb
CP4OErqa8mxlVm20A7PIjoZUnerFFwb6vbnROnvD5VugaeVxjeSO4QuTjuzG4aAn
pXXmXP2HA7oHffrmoxB2p9xir5L4asOWoHne9XOsvPmxj43tIhzVxLicI9q1KWWk
p1jdTGdfCsgGSiPXEFVNH3mcWrTLclGuw3stpg9dCmLn625D9RrWJYzCnLsJ5MLV
aqW1w7LbIRj6VONNH6vYkNeA/t4Usg3GM/dTGK5mO3IwBkPkIsTpckBA0+HanymS
VcPSFz5qnin56/hRC6UHDhiddQMysrE/9jQCs5JVVp5RovLRWIMRnCX05Wj4hcg7
qSCXglALqGwWXFn+15W3AtVTNIAmldZu6zmtAj1I34CKTbmQUVaN8HBwAY77atve
54lHSsoj47WYNjTd3oXLARWNaSII3RkPNBLRVqC4ORN7v94UVyHIwmhv1Va+TnuY
pyNk8aY0bKoVbQbEGjrhkBoYzLNOFu1PLES5KF+3lbp7BFZH4awR6C87PjkdYOWU
sXkaZlyIHuJFoyLNH9zlCwBeekiZNOwhujCDDOuj6Q1X5/NkeZ6P0FjcISp2t9Z4
6MefrbrDcAEXG4hUF5MmATYsJBmtAb9zQuWSu8w5ywtPlsQz1y8t4NhZypygkkAO
Umy03LeV1kI/NzVXrMk+k+30XR+6jb+WJAW0FmfVAK2YVKlEK+Z2ExHMpI0PRSBy
5OQe9qrAVGQk+Au9XpLIvl7CcRC6TX2vUpqzqilGrMb8ZgyTYLskOZ5yv18gwMwo
ygELaT1emx1rB3ICQbnGXKy3WIlDFkWj6EmK5crXjbx1t3cnWQVtATuQ2QTA6K87
FSPvY/vKFC47nJj+vnIAJfnUbFxO+OwArPmIkWAtZqw6K13rh/J70M5paGwBYiFE
oRJZIbwGSCNmpUJYAgJq4xTzP4OTwb+kxPC6bpwqC5a9Ysw6XB7fBnLcCxga6dSg
xkp8SAK8N0JVv4Jxq+Ebk8qwM6jmxCN/4z9iDRNYYg9Rcre45xn+/20nit51g23i
Wea16QG1JiqgOgGPso/ztu2+oPIUJKUZGcbxIZwZDmnMQA3FXxIvavsbhO1DFFHS
oag+Q9e+oeoIua0moMm0+EsfRycB0NLsoU/eFblFZ9r5ElHjy7kP1tandmywBNsN
YDmmknUMB5fhNCGc4oUV75CPmx/z8QWQ7h0mGWEE+VcHea+lsSxhL12zloKgoe8Z
zgvbGuXLlX95PQW9AJrPaZFjNiYwuO+Mwl9Qp5Lr+v/YtHiw8Bg3SAcgTdUmfUtK
2V+T7uM0+HXB8fhczTQukOyIpxwu5s5O8ljG/J8ss/VU78KbB7Gr/H3EscqXdtmU
ktO71lr7JZcRvqNr/6OYw0k8mSnd4eQq53b7yZdKANLgP/dOkNZ7lqqi44rKaau+
m1NEOPvc60SfSvzUWOsWMUVvVIweN3Se5SUiV+cqkd4ncUwp0y9pBSNkrIGsA4dI
9pDVIzf18Pj4NeAaZ/2p2P2WwsszlSpfk8vPupLchyxm9c4jNh/w8J2xKUphN545
q1UBCb/2ugenH3f4q3vtjv2u1wrwO2mMptb7ZJKlOaJq4hhA5oL2iMlTTlFCk5th
sbLqft4pbuMmAQM0JEJ8U9vCRI/tJJw2DhpzeZBgPx4HhCiN/S2XM91TVAgEVsxD
XNK8I7aQJim9bg8QqK8cFitVJlULksnmauDF2AdLavQGHFktqaMsmB73FPTce+/R
vhytM2d1B35buROKjHN5KT4KHSA7YuE9jtxEbZIRsqRbtGj7lnOpvJL9eDTPKrQb
KXANyPA3JGOOK2eMH8H87b7RDD6zCOV1jRd5Xu78oxGmUD4UohsCdWIarWoYfqLA
P+1QCcwbWWn1xY1afL0yamf3T+z0MALGGz5VafU7ClrG7pbya/CuwcWCn+FefSJl
u6EgSt8LtX4QYREyPWn1qw9zGum8staegisGCtg8OWrRjzRcwhl9GyP0HoKzgvIU
FgzMH/G++2QrgmqTfX8pyI8qc7sOTDVZeQeUJv5z17HItC0yw4lAaHH7B8OBqck4
zZw0DRb5xNjmHw5fczJL0e8gZsZrvuOgqUT1gWGPlN6jHJb5uC2VX+rynSi2q5fW
j/kmHnJHLjznzR53qoJ7e0FJPJI/NSj9/uRrhVjOjBkWuywE8Frp/OF+kKubnCGi
ggz/xA9Y+D1JcepCEILYd+2iz+v5kUleQJMs7AGuT1hibB1w4eGEbqImqZz3UaRL
zSUd2J/gDIjbDNgi9e7AvnXcHI5uCCHx26aqAaDa5REw3teaY0SPCzgUbAa5PWVu
wn9Ze371nnCGa9x+s0n2stC5dNgVCJ07ik36RaQUTvXpNXhBSHwy07AXJ+xjk+Cp
r7uIi9qTe2Pq3i78T/IyS65Fto5jtZiQilt3zHuLiHx/suXA05OdXKYZBKGnbEm3
zWaClSfJi+LXSsV4VyuxARviZQ+OPw7ifpf29TaUW64AX7Qpj5Q7nUXCwk7tEpTQ
HTlnjSWpPw5YgicLB3ehl2xYxaKd9hErBHaQAUHNzY6AtL5MiAxbd8ZHp3Vh5P5z
wipq0NV2bgvVW5dbfAp0irVbjQhgYZfI4TePGfUkszbuOrq1LCkE/oQiZKgiiNM7
l+ooTIFsfMDqUxjwRXZR3bgfySwknhZX3WMCeBoEMEc2dq484ISQwGJmW15HSmEW
a9aCz7LW2Su5uznnzmPd19lzCW+zdg0hrKMe3CpzIRQxhbAGaOmKyWK9+NcE9ODK
4ldGDYc5f8TH7ksV2VskGdRiMAq1reGupVpS5plzbodAdezqAToMShY3hyUoGiu2
os9VFhklS3u0sAFxkXy5o/jQH9V8JKV19/Z5YHbYzI7Z7YgmBzGjizUdYUsDZW0a
1uD6AkxYiFaPh7+qaj1pU1r6CaIzQOhWehYO3BTa/PNcgk3iWlObU3DbOtkfvLzA
Sdy53SWrRzTIEOQ3FRvbqrGguYrA4fF/G7QOAl7FCvlIQEJUb1UrTAwV+p95mgeJ
lH1Ah43pCPbxBnC1k5bJoeEYTspeDc/QgBC9IaeIn8+b6klpik79REGwvPH9ltiK
UttlCoVxFB0S4I895SY+T5ze3YTPS0j56/EDSFfgDwtfmNZpCBKe6wCTwj9fVi8x
fVw+xRfaqNYU1fToDTWmubsMSH778MZ5Fk2mbNv2r1YoBWBIMNC42tDMW8M8h7rc
jA02fqtPiK02aEeDkf572YoRlb77eAt8T6+zALTubD9k+ku+YFdhKTHtwvHQYjp8
fJG24NjiZoHL9YyytI/hZMJ5AyVFJWH6MQYENzNCyto3aMiRgoGKeOsacyAcjcap
+CA+XQ8Sm9/JEnnbOqjoIS2zP40TBbXJxIyYt4ZlKTn043XAXzMWYZZtbTahuCzI
XwjwtnKDLVjDmZ+k4AFbihFW22TuqOQ1/sFHGFwcqubaUHcCBmGLBV15GN9N+Lxa
QbaqFymXRg6AMwpLeGJpUVu8O3eEHyEJ6UOcDENM3HKSweIbBJC04FHqrNKdJzQb
dG7NG1zC4fOrOlveCiphQrVsoLPFxD0sEUuXI5JwbQA1ITTN+bNAgH/9TbGm9hSm
FqCcLgnhQyUSkLnHYBI9DiApovLuurPv3FbOTiTx9aL33K9yndNSEnRXWGf/cKpO
oM8bza2DCi2I2JmNr+oQlHgP+enZ5nyXQ1LDsa7/yiMGPm+xsKRKc5daAbzj5He0
EKNExY6SJk8TFKKKkRlBcf0V+opS+RC9RBhRbu35H5XPPd/+cgWE4nObRb5LY4Ym
y0KcsHnnLG+KRqeytZvHTHvduVTkDlLjJlaMTL52C7zelg9mwqhkZwZmlgTED44l
Wgxy1kSePBGlbQ2KCr/Eg5VjCANnibMRZVruOrgiweXQOeGWMCuLNhb8xgpO9kyu
LMPNyGvoDrTxM/qavIgipWefa94+H2cvWjhdnTcRMmmmuGMVLCeRTIwXhTkBmhet
YnGl4Hn7ORo38SBj/rzcE0P8ex9FNUUKzS7gA22bTeLgWG9osrxU5JLc3KbYh5c9
2m5mQEJewE1ZWrFsE/Xr4VQTCG8ZKAacd0evxBmCBuzCaPeTkXJ83Oj7lZ+mkixN
cJNDZsprni5zIhB1vhDm5TVyd1U0sIK0+0O5m1MNTNQmboGBu/AscnpxTzRf1ObG
2OLv99c1XwdxxwPaZueXTuabSWhBwXoXTvctoOVssYLq0JI3vRhI+8RYTQAeJWHv
5j8QyhgFDiiUXS/2gf1Il1yCuerkDGRqcjZmGVOnn7FEM02nU/X3lVMw4iUjabQv
dqpDppcSzGYNGZoSsmZo2Omo7K1NgMXJbpnT7sXX6djiQYjXN/UDTLwLAfyQ9UXA
MFdfNknu2cp/D/xoXbvXHRjORYOQpmhT6icdEsFxz4hs7R1yl52wy3BNvcZMX9t6
hS4TEeC2l6E2hl21tNAlfwl561dAmdYrE/ei2G3oLXTjKEoZ8UQA0v0nMxoo7GmD
kh/uXKOmwTvTxWw1hOcSJLyZe45ipZWNZzDSq+Pe+MfrKFQQRZirhQjSthXtwFxW
iK7WRy9FZYyXF01f90UUgevoDLF594WFMpCtWfPVPGxYyrGbkOGd8m1RvwDgCsT2
fzucWEqs250uzQBKhuqBMiYGqbNqnEqIoA1NV1ATZFhbaK9gYPLC7KatFGas3Xg0
CCNYy/V4qPjTfx+KxM64OzdHrI4MPRrBfMhDBoEtIICoAeMCtVyl0WR0k4OumFDt
h8zMfUlBE173mXi40cOwYA80oDVm1HyA9GmX1J+KuZZWUdT25gIdRdGFYNDBCWtk
fbIszA9iZETlcCAg7aahw7Bcl6mNdBvYQgqzKZ4iW+ql9cJP1x7vJk1bYSZeNUah
7LNz64Y0TkPlknBNwQwE4EE/wVat4STBJKlN5aRCqpNsnyTTTOu2dfoczCawbfcm
+o/plk0/jxrOYs0C04scT3E6ruQk7zLUw8cZ1ZOmqmElhuT8ZtrcIa7AHgwdCi/c
DoEfborzeuKXEi3HfqFzb3QLatP8XWur5N72qtfCJXpMyG5qN/CkyoACkivGEDrt
DJF5lr09KNnR5ET98d9t6p4grxwR/Gl4CiGsgWqjjmUwGb4cmttS8FNzLownZK0R
Pw53ndowPkAnzpdMACkinE3hYwhAXtE3G3OJlCfYI956bsq2qtMM4UrAcKJXkipX
F8BqXOMyv8OfrOLjcZGsubyZjfNJvgiKyxgwcHLWMUFvVZBB5Y6E66HCct3gkavj
K2sj+ejJPLvzOnmvz9SINIj7CoKu5dO3W4wGAl2lVpKpGpxy+LendcomK+tEnhV3
Cq/JhO6bH3OXAPd9KfCYC/2W1sREQcE5Bv73Uu2GrYbqZGE6SVldnyTgdenXpBQV
p0DtGJDoc0Jmz6cf+g/zn+kvtuSf5YMvLmmIlOmUAKUMrsiU364hAXeavP+uKiNr
IGBRRgVpSp83QJFasc6stytijpnH3HGkpcZf5GWpBgDLysDXkl2wsUsSeLUvuVfI
rMGBlq+yDxPq0I+sWGfXGn1DK163PoPQqIGpYELZDmBjSR/OHHc9snyAQebSvUof
xW8JMmFQ9Ei1CQd8SRGZGpnxKOnXvNbgVlrxNsZz6KKruYbwm3GnyqNrTFOfWNWS
8z4/ohyTCXSEz6zD+P9UyaeSkOdcDa6++4EB4h0RdnntQHdEARRdqKZhHc1N7lbp
uLQP2I3Rm1GTk+zgIrvyiNy7nyqs0SV+I01QJSupsgKL4VhqaXfA4WPnj24gYphp
6hLyvVaCTL7J8RiT/klYGTke+VXE2PBRRHh8NXpdY/lGDp/ijq5Jwkz3ahoudkgo
qQ4hT6Gb6F6Yf75oXIMDFC+blDw/DHAm2jjBx2Yte1+yVdb+mN7n2sDKOsdZDach
FiYd0Hl6XDV9bRaPMAuoR+7fDEI+BJFIL5LKbycxdGidXxDwMliumZMMnKfnW9uq
ynE2K5GaOz/+eb11bQR4QaY+oUmpdDYB0+WE/xqE+wZDXaSMqEICo/LUuYMG0Rrp
g1pf3Wv9pKiZOSXmSmjxOl8b2IEbqtWbVH75VovB99fjLk4frMxsc4iZBouZEQGK
MgGwdq2dAtSrfrhCpROUb2PtSgwfNDMNZaG0a17c8uVl07zMtoG5guBIAu0a7TDR
njxoGqMvHvtUcf3SyRekhZgLXuO9GjR6/l8IV8TaWWzeLEiHdOg9c5FtXDA2v4QW
epSrrrXWEI1F5xHG6Wy+cYAWKmDevuTtS6y+Q88u3szLqee2d/kO8I893fs7t0LN
dGBdg8VuDZrjbz473DlHLPw85IBrdXhyRyKBbueae3nqWLJeUoDxFVdgvrGqiBsD
Qi+n1M+gMNBbKpCGxy9i4BlcUtZ6he9d2N0g9MRYXbJ/NVUzUXW927CpSIKsa8n/
1kGFfCXgzfuWVLxKDrfO7Axlxx/i68inpHa1/3GXcXRmtkcUAFgFoZGTTsOen160
AFwONvcGt1flpfzaW6868I6SM0qEFcFmvBUnzuTgjD+FQeagDtKYi+FW+7zUqdSD
ZzDBrr4zVXXcw8f+WaKp6JOFNd4vmARVXhrAganc1SbTDYgF0nyWdvdgI5hypRry
6IUy82DSJkvSEANmPy2eOBOh2LD0jjkj2y1pE2GKFUHWqxKMi9t7/8rfiX2Ca1cc
bDnDr7jXPeyFbTXx4pdlEF+l2ZvauvTUFJX7/5RyvFHszPJ6nGvR9gN1GSh491pM
6vXqQRAaUXyKEBRa2VzdKlZVeOCT5x4wSY/a/yAAei0AgaxXVN5o8riC5QiLbdhQ
aNhptjTu3vPQTSOHemRyR+Sl0rTOhmCRL4375rO6Xg5kI4A/Yi7wkBpHwGHVGuyv
kA5Wy1OgzwxFg26AQDZYJysPhXWmws6Bh7w6HIWXO36ABMe+6Z4gVqpg81GTdnHt
md53B4KP7dUUUxSi3KknfBxwEYhETKCHYruUvPFhDpLO7nfUmZPAcoJlxsQAzyaD
4DLcmMpYZ3TSdztw//O3VNuLcwQwvUT2Z2R7cazViUAUszkgBkJwu7Ov68nqFjga
tmlIKtGdFwxLsQRvGveEckQxG07rAe7WOylqc+lU9YyxdvzHUEHN/GvyxHIhFvY+
gGti9VDhi+5gWsdsuw6gO9CoCCHU6cDtpY9FuFIMgv8okMzDhKljCY9E0FQyu9dc
L3ktgBMCiTxhjuut8f683r+x0H1onGSfVmvTjeSsxRoAKulsXEluctHgM+IeQ/nu
pCB9l52iHUnmpFTcddscGynaJWXM6oj6skywo4mXm+H1NuZaxPFY6La4tzAZVNwZ
6i9Rmn7X0yp9mRUebwCOt7rZqJDAfq648TFwzTGFlFnX08NtKdU9X0ioofOeu7k1
vVXT41vJQhaz9AbDCaOqywCLivfGdhd1KfHJ8DivbRybaMO4+cv43sn0NAELroBC
cuLrPbYk23sf959n9WamcHpf88FTomImfudGT8+UmYWgmEkDDCwxPnBln+KIaGUK
kUTZ18iGu5EPUhlJCeiGzj2gcbwlQGM89CScyJ0OeHfeorbJBZ6b+qEgpgXTBLtN
whcnah5wSiB7yeIeSq+g8pdMgzFE48TNxF0fkdQxvvGF7J94T0P/vAUzK0xeYGR+
hqWHRTLAKgHpzWGLpB/6v0QahABVK2n7sfHg/ophswa8LZRLYi77V0hft8ChIJes
K4HcbNg9QrMi9QLVDC37u/UhhG7+JDUy/Y7Ay4iXgWO5dX6RD3in4kAUjhq0Blru
4mPWcjxxWswxAgGx8/+Z86Q89DHn+nKPh3NNKaQE9Fj+Q74Wh1W6+eVfvs2I8CEx
ipxBLoEH/oUpy97TebGmxTbHHdjhPtMius+eSuYe6QTg5De2c1jWhdS5WOgXQjt8
qs8TTz7b7RmwN2ZOneqd8AlAxmqioK7AysERVbNUZ51cbIra6OJzavIQnBX1KFr4
q1CQA6mGwtgcl5CnxvU+xJW/Je0k833nH5eJPlij/TdTDdBcPNTBaQrprMSEUPEf
9Uk9oI3o668s6hcJJEEXJYSzx+6bhoxb/LBUvbYVdbmjT4mqsRjjT1Id+mUx7lYS
lUYE/GvyMNQKloOPTAarqBgxWiairAMj55Qclm5q5HUuXeWKTkKDia0aHC+AmJyQ
VYweIn837G7lCFAT2I+jf0QJKt7Qh1iUPgjWcb+WsA5fdXVQG6E4Urm4Lo9H+oFK
TWyQDrgQG+9lXmf9VIb3MP2WxGjKyquU/LyVR+CbyFzeziaEVecfNmxKRdbDfIeB
E2zPQ+Ur9UEFJnpdIoXk7fNs3t68aqy5NkusWmpTNjRl7WGzj0fURJLbJcE5o7hS
Exy2wJ+N17DARp+dVJVyrR8dQ9DjvEDSEAitrMGE5fRHFDELxv66VLh04MCoITrw
d8lYgbNQiNfZuEcZY7vorMIxY4jJTkKzxEdC+Uu2KmaUNX3HuPOonbVsuPAeEC92
Pk01XfNJLF/ybIeObDisUOEHO8FQjBQacduqiIwv9nr+aHC8kxwLtBwpJcbVnvD1
cC6mIbWULgB78ZG4PlQ/v7nrDm6Qr/RqXQGaEdtXO5L4iU3ILI1B7c50UkJOOxaE
V+Akhb5K2jM5eeSYbkOXqMpb+G41dsYSvvtx/paAHX9BLmsP0HGJXw9/UjvQHaVI
sDEewMYlHWwjRQANtREYgcNP8TEXqdVGdGEv69a5BTYGd6XCR2KN6c4kmGrXKfjP
VwJ15WeffKLsl2HSl+q1JKVoXaUky4RWNqFH2RZeWACvPou5zzvb3cxC6OX1NtQi
SjPRHgWC5HehPVb6xJWTPINGQCRmYbnOOi8TiXySztgxAKXWv55qVQoMfwdowlDp
NfZbqHGQXX8phDA2oTs2XQKgqSlUn6WOR4A8HEElsBEvr1VIKml5XHWDhW8mD4Ha
m/9jSl+AzGM5RJVUAU8nXz7RJFdgsWdE+J6EPRDroV1GW3hyerYP4ND1RsutVP9C
SuGfAU6ZreZUACAKD6wkcnC1huWxjbQk2390yJJqa5cp5k1cBtu1J2lm7UAQwXsM
1UIEeKEQvXVzj3BiOhJ49htOCDuYaULI/t3P/KsdaFAGjn+/q4wM7dKWn7WLHmnJ
dFGKGEPndW8pEyQbq7USCyKGfnSpayuVdKKOjFRshu8MuYV2B7W8riecQjJXdJzQ
ujctOgZ4Yctvu9vHmXh/E/UtiFa1e7jxEB/62yXEOcOf95UU/D66580z+vd3zQc4
7b79m3x2qG/TW8hpc5rwAfSLcFJs1w24oAKPjmdBjfepFbW9YdHPqtzEvE/KcVUw
6fy6paFQ4/q96CUwkKCRtu6Qmh9VMGfg40OR/fZ+qMZI9r692JfALFVEoooFQkaz
ZRy8Kzp+FBggzHZXyUqDFHnvhDjeyH0pJhvptwGcXqqyBloPIeBRpcgsYIfnk9v0
YB0kZ/OV8TnKUoEfydCh4B8fz2o3B63VyCXPV7dYJHJGMTLAKFOhrrGmryyKsP/n
ENAS67R2vUowJFnRcAaDpu6ZPdnA1Zb2TEYsKguyIJ7HSGLoZYnvgsokrEE236bz
Zm9Npt4zpmcDumJAUyRXwNh2tN+fi4+zurjPMZUM49iBoEBJy3e8AauaNML6QC3M
kCHAHtaw4sD3S53m6VMtv2mE8boKINTFZ7eIniOa7P0eCnvzqHr/hM7g/inHiP4c
lvPrqfm6lR4WsR9+SZwRcK6GloGzgvu8yw3HBM2fDs83Ht4gXl5wrVYaTWlACACu
SQ19UUYpHwvm0gsu0dxry4NlIc+71MyY5/TIgQEGWDwfyTxCGBk0GmUYY9VFWYO+
rJdmcAFhQ7ZkKCmhREWmmoRZIC1bhd/M5lbYkyR5T3zXWFzwibnsk6JeC6FrrERA
KP+rG33/BDnU+ScZrBifQGfJt71Gh4REOcSTkBqYIQfrF0GPSxIZZGtBR4cpSFPS
nJGa16u8yce7X/c1WTdmYAGIPuK3iDCjrVSwJcD2gNH3u7TrPsEHBgUQxPuKO2m9
eB9/ju/oyrFsRtTfOVQXxmKbTP1XGud+l6w7oK85cBpo//82TedR0Np1HYk8QJIV
fK7vvy2/Oj4IAbXjvyUTiuym9R3I81LWcDBX1UcM3movuuGLPTc7Es0rGSQU57WW
zcvaWQm+CT7fFhVga01RWiGk3zSqLryr6iNVDJAeDfPvPstjbb7uFx6QvbaIppbt
RwDGiptvxmZkzYgIBvvFqWxvjgoTMK0CehDkjCaEU/dQ+S4Z1bxNcYam+tLbveq1
fjmCVbUnoJJOMGLkhX/pGtZEjnie+5e7AlodEgbTBsDeFhrWenp7NvuXY7sxE1BB
FMEdKwWm0Q9qwlBWxI9/dmyIsLqZF47PV/Peo0rzGmwHtAP2OmtOIz/zhQyGsPRx
FfSD/Jqn4gYHWVnoa2pqG2jqMlBitmD6f/Xb+LSpUV6GpQt6UidRRqOReJhRksPJ
AcGs0Nx7U5fI5UgFDSyuT6U5MkcawBjA2BhZxucyQkZ0IECVo2NTLKQB6f4zM8Lu
w2wV4yktzP7PrvO1bVlt125NybZbnyEjrL7n46mNH7mRZEk5tt9uetRTRqNUKB0W
qQTsUC+19dW6zHYxo9LNQ3d4WWoOor7cQBE7C35tpQ3uSpfiAadn2ubCfPwg9Dkw
Alqsrie9wKLnvHkTm3noFU3fY3T+tC6k9kyiY5cPKhO1SNPnK9btUE6z6wtl3pIe
5O7d6NVQ9yI2XR3H12STjoyHlluK4ecCkCSMcNvYdimqZkycO9rwE9LcCij1Am1b
nryMYOSM36OHTW6GVJ/w05AcIORMKrY0NUa3DOCyQNDMHm9Q07CC2/Y27a7gXUgm
YUoEMguKVREEtYnSjcCw7mc16aPP6TJ7nbrwrWM0hEvH5+YH5ozg9otkkzlLMFXV
2ngFP/XFQCCGOKeTQRLSivUDqVMUTiLErb7SbzlRIEk/kRuhEuYiMqrlmjujO8rw
/bhX6KnZsg2DRo7ohvCtETXW7tBHo9/TGAjSmWYIIDYqAvIVVg5ViTd84LRvRajw
1FtkJnoTZ6vrDUp+Iiy0Y+3Zye1IB//InVbIbuUWBtIoaNakLfM8zRT8oAZOgm3y
v6wmlEzDvL3+5hhTqCNlYGbkAnKiamUt81zlnhji/20SwqGZoHGCgoC4au7hUH4y
mpZEWeZ6x7cZZxICf0v+d4oKDE0JhAAsE0p52DmrB2Pt4EaPTlfvUP60sycN800q
wkSzBKiISOJrXICdHWiNtFVcCWGP1E40ucOcddbsNO/DKPKxBSIifwWO125Ao5AQ
SL7o64U/ffbSSuBeVJqvo7g1uvQB4SZw/jA8SzpzYtLKXGeaZXP6yCavw1LGY1LG
NWgoHvqsFH1qF7cvhUXaz/79ULOlgUsF3kkTrTJkG5Yxgkmyz4SDjqf+Bvp19yHm
JMpwH4xYjSI+4TrnT13n+ee5tDrLt/l0n1pxzzuKyIQNVwH2fsjzPXS1hge5GBY8
cMWOubqqg2zPBhYAs8lSljSOvoFXq47GOu4dt9vpELgMCzEcdlSURjbWX2xqjEn2
9rwbetQsnFCYAGtqFiEAlGQcDXzbpHr73RwkF3W7jZgIMJr9H6jPPHShtHoa9ytT
0UVlCDD9Bo5CKZFAX3PD61IIjVuUodBh1Z4b63Ewh/KM1+RFdw1tPSdkaxSnqE8d
M10qQU30ZZ7f2DrUXOn4MVmv8UO83DnXNH+FuOHXaWb9/3xtpl4/AKPkgM544gI7
BgCeeb1sSa34JzE9FfT8sN0XK6QpeYsvmhJ2vZPwRvoA8GURUV8vYVsk2ekw+JBx
lTpq5b3yn55DS0a7RaZbIxbNi/v8h4S+1dUf7DTLxg1MvEnIcqKtrQjh7HtSS2A0
PnEqlzjG7iMlC04253BBPRdpvnaq++gBDiuSMMPfLuu7v/SA0FR/+/nDcM9EY2hY
v6kDOypF+gKq8nfvJrA5wb8u0R980F2FOuywqg/zlIP612juYIbTxKagi8S2/zn9
luwc2XWGeDehQXGolyeHcnkGBAn4UlFm4997cQj6ZPuz12qY5pv1uzW+f3f4hpJe
Yi1gCcX8yvJi47fP+j5scwk69y5gu2dZ2D4z+4ZiLZv+6WgjINu1MlCLxJeUPGwJ
qCbdGMWdF0axuDOJWzx4J29LjpzgZNVE090vfrMNjHISH8oRiHG01tSfK+IonxiZ
5CYZVkQY5ipFGaZQ/H4aZz8yrcQ9LPg0Guc4iStDWdRQ49L75VJoDGHRO0Kz2Nd1
xVA4qkfvkj0HXPkU6JcfpahneIJkDhDK0Kx+2OaYcENuHw1GZtxBzHnQ3RWLPMnj
Abbo4LlkWrOIMexQm9DxFB0Nx34HsSUB66NEm/Y8q739De230+my2nhqrpAE9STw
WhHfKPkKJfPuV4i7zh/Hx6GabwvyDJqIMhz5Rw5q7h7nxvAqOBP9j2sEeQQNqJ7S
udnA6I/eKfKbOAl8Xd4Qr0fkp50sHOuA9tnekGVGamCtOqPyWs+KUXw5mBh1u5Ju
hAQXYMY/gMgznIpkgLHuCnqMYMMomRqtTAeTqhQ1vBTFEUfFU5dyFIBoSK0oTOB5
MEV+cfvaP9wTMrwopsV0sjpjTc4nImm0E6/L23+K4RCBGbKddxoDy2c/LZN6lYmW
YoZOBZ0oRj0tkyCzpWWEKNKNPzEYsNkeB9QF9ejp5W2LmrDv5lC74Ua1EZlj7/Ij
99UqwrmaXcsM2Dw3HPwiBzTvbiIEZd9DPgvwwa4N1KYqjWSEIG/LhtJ+/0LXJICR
oFyfwq7vz2KBso6BcTm74PWrBpEF5zR9GhMgo9LyTxEzob0Xj3mmeYfKCyvgSZ6N
4qZRa8FsmL1ZnVLzAhmowOZ22sdCQg8n7HxanV3joyn09MJpUgeNgfnR+SclzmDR
vQYin6Ph/UxvFOax+STf6J0H5rlKUhHM2FouufrRrbu+aNW1HgS51jE66NHqodLq
Yjzu6AUOXd5lE0yKYkvTzrftmW2LqoiS3zBDd9yhHmkz0OOvDKS9v0dBgxePT6zk
H2YKtMDPHak/5ay+JIUXpvuUwRc641UY9/B1nPVU4xZs1AjoQK+dK0Mo02gUsByp
xtoMpEl1S0ngP77WbXqjgK4/+zZrNAbmZ/9jtcQVm47MXt8t1/Ly0JRfrMm2mYUk
dpKVNhdkzY3BPpcsZX8gjWQHEzEvXz3eWThOpFqz6yXrpdRdjmMz5STyBwarDnkU
SWIueSRq1t5FDk4ZYtgOpr/342JbCBE+G/cIyaMKQagh9abaGyPyHVbx6HbBKHDw
O/qgcRhZwgSrQKShVe8lgf2YmRkb2YSvA6jZ0GIOm9Vg9Tb7bxLmlcXvSmUTlisV
QTabjKMOYP9pPpbhS7DSFpAYbJigIn4YI++OuhKQSw0k+fqimNNrYAQkPia7g7ZP
+f14SPp1w2YlgIljoWfyzrtLiYwGcnGnuBrPS9juP4qgXnCu3W3o+qL6BtIYeVEZ
9QWd/AT4Kt6l1N0ZxN3cZrlY0wrMzKoyrd7nVboxmUnFgE+Mm68t7TCFAaWA1Qan
naXHL0t6OSm5jBIKpirmvonPw5h+m6zCjSE7qaEZcvcjK7NFWDAPdQKOlkaEzLf0
YoEs6wqc+MW9pdAW+lBKkT641nInNh3tbe9s34FF48+BSDU0UQMxPdCcXOdqYmyq
ATZ59SXbdrWpO40MvK1oUo/PTC0tOlqFwNHoKpDH+zavDkvUQ53d2niwBKtapuYO
ztST0VIhkXavD7nCWi1ZZ3Wr9pF26UBp1iJedNCapY8cT94U1F8xtNPprjqF60YB
oBdkhEKZ/5Gta8EraauO4U5R5LHOI44FPI5jLd8ZOJuDh34p50iogqR84fa6D0jz
StQ0k2Gm5ie80KJRvYhE2YDiCpUQv5rpih7av4rzekkEb9DPMEWesZWkGGnf4HeT
rnmGJ09WZr3FShYa955adH34w0YrkncjaghJPVmI0TvZrruM9dBo8aJuAByeMS9P
vJxlmyEpSbqpIPLC4VIBGSdQgvB+gI4mbybG71zQF1Ctr+CRWAGckXjOgjiDiL8d
WU5Kn+3IPzNfRCq+epOQS/PlXD3qCAA6XfBVblYyAN7JyKVn+1Kwq84VAYkyZSDt
DtCG+3faCKPBskjkLLLVsvzoygRzvcfbJsTAmBakIUtuG0nLYJMeR2Q3J/3vwwN9
4R9pNFBGqR5eesNpGW3NKuUdOOJLkUSpoLGvdKx2GkRHq6875+jbMLZr3pR+Ta+Y
f7nHq/x009XbDvGJayaEv6J0jUwNDwavuONbpSXUv1rIrF4lEikVp5rgzqKApJMd
8qkJMUt0RnwJToZwwRPbTWDVU5henugLRMxmL7rSzmyKibOPOvqMuQQqYNjlLOCl
odYpi+qjQVnr2FSOn62vsf6jcrLVNp9NpWKA6h0aWHSXRehZQH0MfWl09V+B7cTu
NuRN96EPU4CpMK+xK7lBO3axPsy8+Dn4mJzNmw97h8gNBWn3ug9uXt7S3430ha2j
OA6885CArACf24Q/yDz/ZvZNOyb46BDImEwsZyruFX8p70vPAVz3TwswP8B1hUIf
yPV7F7y9FIdVZJnxXak3zuwsWzqs5essgElS39+iW2sxNDAlIHeKYCBkuOdtv39+
o9/SnLbOClnVam7bV4kw2g+g7lFxstazm/GN/YeTkMXDPNZLUWtVPUtKpQm2u8MO
RDKudtEvMko1uuuk343xUsX/jxaMkAasSamKsbBT9ZTAicFcZZN7aVizAWLRxq+M
unix5XLnpojEkYB7BqF7dUq2B/mpxiPra6BuzczYnIDYAx99+poAVCC1qECUG4Ep
Llkt6rNIZsi+oInwS24k76KVLxI8kv/KVJZnKUXwIkQertI6qOPoW0jjApUklqSk
/x2gIV7QbRV6Qq058Ftr6D4n3Pm8nW72Y2oUdjaOnArgQz+5T1DCinKi2RwiPwcK
KLm5gh6iPZyR66jn9ltQHGoPqyLq7Tuc4Y6a8mclBsbGPGN366PvJdqI7D2xYOca
Bh9QYJ5YPzm0OKnkbp7QYha3tfNhr6h1j3EH9O77sTNk3j4XbUMCHvg8X7EDTF1B
rE6zEcvdeyqCI0htkmoN7/2Izlporf/KYoWNqn8th1Jb07eOhalxvQnJa5ORyqrt
jk0g3KN91zYRp67pHJmDsRuhjVN9ARoiQfAUSfUpSes+5G2GN2CGyuIsNu5KHWuD
yYT9EYG9UJqLHoGQnxhdBNDrT1CKCDXGaT7cmjtoP0mwZORTMLrEw9pGRc75MCa/
8LHoFkv+6BRaloQUkJMT9vGiHaxPnKZA/asK3e6ZBLEbzh1N63cax2NShyJQIZyY
FUxcFVm6OzSNeN+k0/g+06mzZ3u/dEdQJFrNHIoqILYeAD/yhNp9HaXQ3xIWDfYF
COA5zC8Ue5h2IdV74BCb5m5Y2bF1VhHfq/Bda2P9OEeQ++5gxmbZipNOnLXNBYVV
trbp9QP+R1xFYeNZ1wZ61b3z8oEmNIC9dZiQWQqgeSjU77eqKknj0CNwww1zZpFP
ax7LQqaJ29LOYO7VAyWiXMAG+XGfMNAoQha6cxyS2aeaRvhg+tuKwNsq5SJRtynF
UeF4czyl9mw0B5P/i/zejyOQyzzOIla42UvkCA4eu73m7ePI0jsNQzQcYS7izPGA
8q7XdsZW6elsZz5uPIohfZBxYHuXWt3IkVrikuxcm+c503a7BfiM60sj6BNDgJ4A
tWfY0bD5xgxxLBpqScTA1swGUsOoZk6mP/8t+auLRq4HEY4JQc2voVzOLUQxl3zQ
QgH69hntuLBq5UAhl6IowYxKWXlY4L/eAi4U/ZxGRLpxj99tA+lE8xH3hp8IGxF8
cQAxqDIKvmhu1c79NltcsjUDaqtb8HG1HQEqcpcJb8Wevko8gsgA0gbA6YBnFoHk
lwQSFzGgaK3UW1ANFKEwucZymxvsT/Aa4oeDM0YAKPXDpuElVqhV7hvQZlVHWmZ8
aLBIz/4rpk9D/xYAR38ti117nQVf2HoZ6pAyFjB/6mSuuatS3QDvsMABBjwlZ9pm
SBf5NBs8DmuzQ4xrBd0fcUOb30uzrkY4t/m/LCC6NkrkFOH66s6pxOaXo+j9YRfS
p1VSLnW8Uwt+i3dbrj6Hpo8BV90vO0uEG+14db/u14nXEdoSf6Mjfr6rBG90adau
kqcnLaYYyt4/QpHUTiA+3FRr+ev+h140JkOSuSAJOJWZM7IjN4jGsTPVWDs9FK3k
vXTujLZ5H71JRdQg1Z2ptpFK2XaIplmNDLdd7V7MjdMwZG7kbSHlpXbV0j63xVNZ
5WA/KIgz5qY4b0Bd+HxZx0Zcf+ep9PHyyFCmeXqss7a0AN+J1fZLaExdahnKB//v
F75dyHnm6VE2YZskwfzVYhAx9lHWvSqYy1FX9Axgvmurd53thws7rRrHWqowewSr
VIFEE71GmWfXTJf4tR++k5B0n7uReCcWCqI6FB8W2dBDP0EcrH1cs9qNSMqKfmTp
DaMYNMJ5bpx8Qv1ihNJsEo54akNEBEKFZyai/jTa/0TDKOvXOjIZ+pCClZ1LsxS0
bvwculwtl9eZTg4dPNaROODB0S6x/ecQMLVyEICc7ei+hzgJ1hGXmbkDOrZGkoBW
pfq2gtLmwU20CoBYuddRFvz9Wa0JZppnxYKYGchIOCJHC2zXpgqfEEk3YO7DLThx
KNnNzio8SmupSPoL8egtTulQtqDnfDIy4I0d1wtKgk8cjS/qEOH6IZiPSB4J7FYp
mJHt/D/P1aSTRAaQv3T6+mpF5kDWuXBzV9VLni9xEixEVaUNhFVoKMwmFSg61ok3
8qKyqoVZ/g3zO8fmHhBCUA0l24WMF3E95Hagjs9jURGlTvTJEcAZmGlXBdtUaE/0
I3qRfKsXcoNGPCkI00SO88YcYHEIK/uUuK+jWnx2h9Me4FhPl4EAqmYH4p5m+PtV
CJy59s2Zr64TB9mDN6+Pjr18wO54FvQ9RQYCJmwyYx5tyN/w7fcscnbbwvjfRZud
jrl09ezFhBesgBEk55RmiMRA68CSIO1LNSrQL3+YzEssAf6OOMPsbF6y/J/al69X
xWLxPsIx2EcV65ugJqYAskiy6pbEYsb5tbpfCKyOadL1gylVMI4Rr4/clvO6t0AW
0kKNuGCb/YNmbgWRFO8rexmrXzmJX4ZAAFdxUTWm2eTTIpKFQaJFNGUuC3sIM/7y
LpvK+MvyaNsoYpxF7Omx8i4OiWnF1Z5eN/Ils3XJgzbe+f73L9TAoO0OSGnYzpj+
phqWvjuT32tKJm1r05Pb7xCWMYK+nlUH3xV2tipSxce0C1NLEQb455CSWsZj15Pu
ywR4IcMoqAAPdEE2oGgKX/6HXcm6cGr13q4qNLrkQo3+zC2e53J1KNj/Ye8c6zDJ
b3cPqHayYXplBx6qIAOnBmpcbvU1XhlQKhLJn7mrV9pH3JMATKA0kq54LfjVMbEe
j6+bdziAItGfr5GJyBcwRpBSQHNZeHUarCErYRMPGnLs40DbChw0YWJ5j16jtDSX
7uEghqVz1fZNSuwqxcmekww3SHEpPUqxLI/+O4e9Q0rLHBoQlWQDzOegNtH1Xom1
MRdb7sUJH6+74VKCyfEtK0sEmnW3y8Wprm6TWJWyhUfVEjG4+Dr5BK5UqlRbBXMj
+oANd4oUDDfdw0YAZWNfNOPL+RA/ZyS/ndvEN28VyL0BWmv88QgjEBfGaKwkL6El
lZ8uOSC3g6lKHKu8oYiXUyMXmZQn8YEUhnyDvqGOOod55Qe5JRig9uZ/v3d6Gf7x
CXRgVmsLEEzHim0SShpHt6ia/JI64qfcUWeXZNhQbPQCY6G9zn8tt+9ZAoTyb4B6
UOVwkRcYu9VuYqUiBlyye+PKoxinjBCiVK0a/I8KqJn/KdiwTluKff+uPirU2N5d
w/mlQJ0pi93Mijx1uyDTQjOZfj5x39oOBG+I7l6AWqepSh/vpjN0TnMD8QgRabj7
tMT2aGI1i4hSU+ap/XA2926EcMSTFsSpwgpzWzEOf1C1X66aMM7AJDQf/+rwEoBj
HwZuW2pPilsdpwyXPeXG7jwGdiR3IrTOkPmmj+CZum8SUJI22BMNah2ahkTbFHCH
9gK6vobCZEl+ZE95xl0J6NfliGYPkqKhtndMXK0MBmvuLSerOzAYZ+8UJQ8iDRpi
K5y/rJDEeurGhndffyDoUe7HZ44Z5UZ6gl687D7w63oUwMiMY+E3WikbOcExsxLM
yqao/M9fhCJHdtvpOQ0dHmuj5xiNQ4eiD4dbmq4O88Ysph/RYk8Yl6sA9A4yS8Vu
FZGXEARvUFya32Ffa0C7JFoH96SI7Q2EeA6csktQHAGxUJCIinA7WOi2oRDXSNvN
McN/IcubqJ2LoDu4cpmylD/NCyyDR8D0iYTn2OOPgA43XAKPhMC9bBlidh1E46hk
0gBU9AJLk8nXiodm6PfSb+YxnM+gS1NZ3JyWd/sAseGKTGlUp3hpFgXChsr67MVT
ncPKsEpofrEeliyOlOz0mQho/G5UBCZvqaep475ddEWw9FtmXhufFt+7s/jnofpI
3OaA/8cssbDCRIeAL/9fZUrbT/VPVyPyJELkkx6YP2ziOeB53aQYSmhZvN++hI4e
CrHdGSBsVa3F+wGnt2qoFDnQWE7pxkLeqN9NBBbxgJIzB9T/NSZkzdcZDHrVKmNg
AnU7iRiKMNd7tLHmeNpQHJZ9BO4Gl4hm7/G/xQPts/5BX0hGwMAi0sNB+19OyZNF
F9bPDIVr32TuAmDkSHDkjiwOCpaGPMSSlkUH9yEiSyfwrsPJMQZ5h83wo5J6OIDf
RprcPXOW9HVOfOb3YyzTGHYu7kvaIbuj1cj9eWCH7oWW0cr/4ByXOpPUX1fUr6MG
HlOz1wm0tspv0OhShzk98djsk2LvlzrMcaqTks4d84NBWT4H2cPkzJ7LBGFtMWbx
4kgJ/3Kv+peFZ77PZ5eHexHBVw81VQbzDcft+t28VVYgK6b6HLXIRTP50Zd1wYrL
MdguyV4P5+TJplupMKH+OGfBUKvmPL7Clnjdl+2oLL8+kw27jRaxuTfE+8w06lwi
b7chcNueAmVLEvZjrvG4pN4h6/U3J3Z+2AS0/KMUXLAnzphK0yIa3C2avryLzFee
XwPGn0wEnLmreef0VpngdIwZG5ALnOCOpqWafiWANjEnv5MHQQZxNrh8stxrfMwb
Z0z8YHtuJK8yiknkJW/ezv9vQV7mUL5h4Ms+aHNYWVBd1zMSjEOTcS6zDogulJi+
ub20Z2DTaCXAlPhImGiL54KapslObhC+P7aXBX/QEkGCk5E/BCyoDLb+pqvKejSH
A+pT5xT1RTO9z66686au2dTl8JrFvpy51nAMV89Dy3WGQgFUdY9sTDKybeLVC6Os
DLtvKhmFMaDRRWMGYsjv0gGGukqzieKx072OtoXkShZpqJX1jC2d1jQVJDWDIi8r
ecbXQhynSLIt854taD5t++FN1eCs0oH/+sFYqkFfsu8N5FORPhLOCsMlvIJgU3mZ
9TutaZRHlTrMkV9q+++dgZMtJxtckaMqCP3pdvLVTwtL2XmiDIHcjbo6ICPlzjJj
7xLKr4Du2ZEF0l/3x6cXy9Y3Xe+yKOiyCka8JWtuqWdq8o3bEYw48ZAF9oIh5V6h
au58OceD9gyjIeDwXn9zx0ylxR0PkPQIL6LOwASas4wWDnv4UZmVSnXJGhBuXGlv
IWRzFprIDMqEdJSk+hI2igDY9e6+GfgV1NY0wFgUuhft8w/Mxf/sKFgrjlv1qXCF
ZbaR3a+YiF2Bg/PHMf5Bu1hizShIrISOWE5bPdAYCeGptextj+uhC9HvN6E+iu8j
v+dcmaLQJvj2c0nRjoRkb7cVFylThC1qdQFWI41OEbx6aNcz/MQFzdu59bbUpHE+
ZX0gmhP99IKGZbhPHmuqIy/DdIVEWgfMaEwTlLcGREPPtnp0cERgXlvD05liQ1qv
1zFCJAEIdJ2OESL4xqN284iOMJm9FFVQCwk5ySNexn1sQlbVl+E7Ofv9hoz+NTIG
dTdhjH9Ij9+mcpDzgv9x5Ml76jDuu+XJQsXT2hg9ic9JVknb0C2N6lpyz70Ovv26
/m+wQM/CUR6H+p3sQDIpt0UUACHUf/IFd5nMdgjxmYvzQ3355U5cFiaLUreCKova
t0xN8qrWJfJ9MD+X9YVyLebYkLIahONsR5U0teQ1yY6X7qk3UJI3nGMCRECD51r3
7s89baz04Fb8J9Y08G1nhRTS1Z0tOQpKGH4eOujCSyJh2xHzpv3aVOM+Pa01jW3w
/QoJL10SV5QTsIeNN6xXRqGS0xgd1v3us52YxraC9L6wzvsSsbdV5cbLOhzIPoTf
GF0kEc2nOcLIN3TX+emtPyHFwI5bjVthFHFc5qpcF8FpMl+W8V1eIxJgJdkuh2w1
jY5JJZ+7foLAcKcVNi48/lKVJqnI7L1bgeFigDkOZoHB2uiZxtaUoqHt22uz1kp5
JjDW+eI7xV/atXL8/9BlMRV7dzI1u+sa6aGUIVfi8nDqSKArofA+ONleCjFoZLid
8n+CD27Ei9N6QZ0M+Z1/fd4T87+yCma3DilFPcYudRHNdvS6ckF33rpwtZSGwv5E
wK3gtL1Q/wzszPCSF0uQa9eNufdxv39fvd3+pId7x/X8+qZQk/Jq0jFPI1+Xui3Y
16jGBwgzMWHzjuHQWbcys8JlTYClyCZo9xEsrdEBuNKCiJgZ8QhjYBm476NBr7AB
/oSgGtj+ZPdP39J5GDiWQpOGTVHdyX+mCtOpVk3N419tvRVm+zVp+DYyeSZmRLCo
/tetYh/okhC2CLjcODA1fsKshpu/QYQRB4nTYI78mBCgGN4rf2MzE8RNgHImmKfP
epUKf2uiOuacWIT4aIeiJycv0vXXQ1kE8gCgHlYGSDzdrmBAFX0YwWsxyAVR7y9c
ThY12o2a8vYJ7I4F4ieQziphCdDOhc79gaVF9cGdv2AvGDr9v0LjVS7XWNI1RWDd
WdNav+chA7KPg5H+uZ4wVRtnhmc/9cWkUcHCAXCcUacgdU5ebrwXMLcgLY2N5XPw
kS9QhmCE+FEt0NIRVPZT9LjAiZUk611fGTAgcth+e+OENLJ1+pfccnrpY9D4jezj
dksY1UaYnxE9EjtOl7TS9rTlbCHI1UpoKfT6lzORR8uIiZR6fxlkqGFrZLHpFkfq
RogiiELGGhlXQvus8RskhSp0ET06ZpVT1sUMsGXC3ckJJeUXgc2jiB02gqyoAMzy
W/QsHH//XQy/8fkBiZb75aaOUeBVjirsDzO/L0HsY4g47eehN53sbHVS69XX4uBK
3RWf0zi0AqQaAkz+Hkt7pGIABIZfQgskWo3TLHVRleWpgaLg4rFfpPA4Tp5xHDWL
L0qwlJOke+545tE/MvFZRlWw007sfqdngs0WDwcDq9MjDu/SlpVfqWF7eWaxJ9hH
knyjgo51AKdi6cAkcG3wa86MEBFIdjvBbITdcf384swo2pK5mWRvqU4ycWR7KQLA
9indiqYZzla+ciuHtLRGBUeIwrpACKik6biAYWviBFza5PSwb6734owHKATeK86U
cEaAQyiSx0VyWuTz3Ay3i7/7ASGUyODyFT6P6wU2ty7FFZr/m0Wro3RUR9pUupWs
9nzubDsAx6SPuu+i1LU8wfYLob/vfiUWzjSwDDJYtxNsaD68/pbgnXXMs35vDDK5
AQCCfrZjAWzkA1e+yCtf7ibQTAhc498hmb0dqc1+89wGTpK+HtGRDLAfo4OIbQFG
U16+63aqasuKthucUwJW2J1872OqXVfPI8ub2VNdhgJ8W0Em5BGur+NGomVhItl6
yUERLRhLVOKzOP+Z/GxN+gdjijiQx5iy11/d45BTn2zBTOnOW/GD6JImICYOZDva
d4OliHS28m4sA+alVLHAgMm3onp7AKLZiontiEVNFYXhJrGLQU3z8G8pYx9TaGws
y4WL0dFlWy4XbTeeQoZvKZSPyQGpwPYfw3hMQ9HMGYhTD6AgIEwe57azYwL7O/8P
6CILf1Z4AZgYO9g/uVcVex9gKBt/e8gJoVD9o+O4NtZKdFaV+fIyb0rOFKLzDWFY
g4qHNzY6hG+t1dusPe69VYgeJfLgWFRJRGcfI1HU7d5S0eU8ILjp09LUFsJhOVjt
aaS0qCcf3x0Qf6C16KLt7WQoSjFozqa8X6Vj9zQi8HLV+Q/dFcPNypfcH1iZk7Od
DqwT58YWSS/JvdHMTi0j7w46oNb1acJuMr6JG+o8GrloL/MPqavoxGbbZJJ8VwoU
rlnaFjXrE3q502jGsWH8VU2/XGVUcjp3qyG5I+ZCjv38fTU7Y4RpELw3y3k+134a
97D7h7eU711H+9kU18LPV7HjIDvkGkXtBcfK5zzI34rj0a3tJ2cN9gSBNmHyHcAV
at6NOyjHvTd3IPqJzJvLzHdwTyGNMVHr51fcaSszNEHeQiHh5w9x5vfOy+uupNkH
Uqmm9jm2NgH0rJMX7LYryHY9eZxatdVn0qJT4FgM+zkIv4ZZNXGTuUwbq8PQ0w/8
MZ/MBgMtZAs3VtyTFcqZw/Sk8Qq3Xfnlw2A0TLESW7tU0GhC6m2499r3FOizetVd
kg1mRx7vqFpOzfnhEOQ4CDtkehqg3FjoOIyusuzXUoiKFDbycJF3wcCRpArGLkU5
kgSjNanHhMfofLBLlxWpmKWZCcT1fFWJbKov96p0823J2bKmrNA37QeyPnKbJ6KS
ct1oIdWiZKjeBhna0JinH6RTOuaRb5+BrU6qHD7q0ONyEUVNuuFj/vldGsxUHfhL
GFeoDt7UQRRFm+Pb/81AH8gl/i6DBdLARAZj38sT4NzU1rFuG1akYY4JE89Il4rr
8+e+Tsqma4sx1szmZTV1QWVo6QDs9JKQLTywX17+Z8vgv2O6O5bKaAZSBs9qogFw
n6ySVDkjA5797Fe0jXdIlPFZsrQv5g/R/WUgGrI+4Qj9Se65uMahMxe0ThA/kphC
YpS0aPXxN4BD7PIJxZzeI+xZsA4G2SBp1w1eO0G4KGrI4SonWxu7txsLzmiiPeUq
N9xoA67feF7ysCzqczan8GZLAPgzhNGAyn+LCcDs1NySE4KDOAraUyOibnKvg6pU
n5jWxcM7xTGma0DDoh+4Pvt6Mj58mzvAD5IcdvtKCMUeWuzn9f3gnv8UwZInwROy
DzSxYQ9JZT/1QhhoHE9BHaeldS574wX/s/65VIPBx/KoCuX/hrPlbwzYqk0c6Pcf
S33yMo+oyKGCb68sqtuBGJfLX9Q0e2gCkM2OjmuoAOFVUDez0CRBf8sR74Homimf
tHVMDK1SkmROWCafUA912iybzj+HMHb7Bpxq3n7tJQwCRQiWjBZRhwkI1V0XquR7
3AnJduIZyDeVnZyxsK0GcTmpqRKtqmFTz9+eQ3p5tCPwILSlW4v56gDH0hrHQVdP
HzMA5dRREqs4vFF7Mv1tpGxhvP0Ve1XbtHhr9r8hYMWnp6H0EppTbdryoLPG1pKL
x2OuvWvTz8F9BJ/FMy8JtrTU8l/XiA6vU2jqJLV+sRcmc8MfEOIXw1WrrAPJaiTj
KSWN+IZxUN/nCxXjIJjQ/0S5DMy3UCEZXjZZEykwb+/e0Zz3O6GZVe1VOx41VcQB
D9mQ2i+FwmZxUt+Re4V+yY95L+w4uWeLzU1uGB8i/ibWGFJLTcots6KWEv21rT4x
Rf1FDmJuj0mCwZDEBmjDJ0tKNEdEShKIgwLTBtnoMVda4M/M/Qo+41ssN/0CUssm
N4Qkzq3S3pxNLegC6cD8CmEjb1arZiOYl+B1b+lYSViZjY+rqLYLWLfXvdyw50s1
DW/BE3AsiRGMv/OiJBWqh5wGm72bymWkwEzyfJMh3xtKiGj7PjLRhqBSW7u25C3E
ad1L9tF+DOPelmKVy3ttkiI7o8KTU+zCk3+GBF8fyfxBWLWnq45yHKe5rBY9ncfG
Z9dyV2luB8lwZYFg1tq2KoeNZJBfwKtcBOgtkzWY+h0IjP89vBr4plbSA1KBwmp2
ZyQQyv2bpp+MfMSoqQgp0YoBKMYh0cfJ482in4513mI/sAvL/dZhiouNwX8ZDM7F
PA3pHoRbTUEM6YfeOU4eNwJO1nAhqWia/UE84LiV7mNGzrLjNSGfkGeP9wO5HV9B
UBwm9rr3fCRjhGW5QcSwtnaB2K3kUmIJAp9QOmw1X6owIDUY7UK68jr2JUWQQlH7
aqNkNoV+7/Zwy83X8V64DVFeTyUjOHQNlsPJxBetuXb5xJ4aHGLB+WrIunSfKUJV
zQEuK2vu70xD9JvPSvUrB+1STND5dBG581UaF2wyvcKVguBcCmNyHT6h5ms+l914
L36+VaFlhmHQM37bp01E4zyCmqC7cvZo5Ycs76ZpC3tXYppOAEF+50X0h/awTs/A
4/PK/z4ZBALepCaP+VyEdM+IoyoFEJX1Q3euUzGt39XlQZOBMeMilQCNSZ+cyJgm
BaQBIX8jun1A0Mn6fcQXGYYywe2m0vP3c4LIWxbFMx5n5st/22GtITCtto/GvYQs
t5AjVA8aprCdfxgkgF7fWPMP5iHoN43mSJ8YxWVJMYnncB7ruZZTETkwIpGRry85
uvLZORekIiebTscnTkugmz6c9B9fsqj3X+jRMQUXiXzMkUUw8+jxOG6t4W+ZH28M
CsIm+GxoLRC1u9IwlSXrl5To3mNeD8bOkM5v1O/j8PIyek5bRlVAnuky7WeyrarL
0WS3Us9QGAGUfO8JCLyxcJJAUsfV/EndPnV242HCY2RGEF6y95UejhzV+e90Dkr2
j5GQcIGuJHPx32lcGWo9yamRrq2xcNRIOnUK1uEy31EjbmNrHxmAzH5t3aHORwal
s6eBfTfjx6EdyxkvqnON8iFTkBfWOj6Tv2OFuP/l9nDpnYbXyJhwdTJPZj8+G/Te
O2Sw6IzvYeScY+fOKE1Hj74yiu6RMuahkU5Nut82cTNuDMpkRuarim9ZHvUIzaEb
Rok0pj+6Jb+/YMbqrjpW/aSi9Z9wYDCck4ZUsGITKQOh9wBiJgCzfqdYm00L/V2P
xmShj4/RxI28TWRbWVP50SgDfZA0uaixQXb8G+FrHRijNxjafiKHBkhmdN38I7d0
Ev9YSMAglJPQNKtRbUZunzN3s0wRv1wIa4mHoyWRjJKrVj2yKGy0sJ3eh7wB3Eop
3BwojYvMNR/0Wkc06p2OgWadJevoR7Zk+IkzbieyUpmlbxElLFlTKR9QnubtzoVT
qd5rtjwSLaQyWbM3q0KX1Si17OZvcu06emrCgiGvYEqoBVAgkih/4az008MDJ5dY
+ik84rAV7mvVBMvDdlJBiCTesg/DqcG4NGTA4GgRXZDGyfV6y/QhkPpT6brcr0aH
YkrTjU6Yefb9kHB09PgTIMH2gBmgBe5T/wBwK8yuCWF1Ly4zJUmckPu0U1y9Hsf+
e+pnQjZmpRJwrj1eWm9vj4JvZ7J05wVimUdWuksYqxphiUyPTH7QPWs/ekD7W3iF
hV/OHaNrTf40E/93PmOirh/rBBBw+yb0Yocf235UvYtwh6BQTro+cclZZuG7W/AB
D8Mbdxunn6SHZHGQO4ElhnmKHfejf216MyDC24TkqO/x4KvVEfYuTPw3NWBYp48H
tW2e7gPI/l4CmSdIqAwyMkn0fzh1ad0L5DDdHXLnobBB+PUZ6o99nLxIICdaGEgO
Qpd1wvIKUt2GlTRr1tvfj5RRsuYoG72At0+mfjfIg5OQmRD1jnD8G+SMRjwmq7ti
a0WyklLQ1dk0XGnMzDhOqUKKyP9jwAIuR/9uwyyBiUB0b+8w7UFCwnxvSMGP3ULo
yIj2UTYIxtMdDxLnOQePZdw1u0Mi7yz3BVFtDVJjIEoARfr1COokwqlNAFoRveiI
T4ZAQLQoOu9z/bfzT6DrIQjt94RtbPO7lD2dIaM/mDAjhC5mEO8qmNV/YZoDegqn
8ChMBGJAZhliHuQYGcFO3oiavEhdeNxslraoVio1DtENcavHv3DjuYb6tecXILcq
8oeZDSdpDcGMMQUW03a3ueqEVmN//RB+fD1DdFz5nolvy4Bh2soaz45baE67rrtM
f7x4eu8cT31WKclDPY+rF41sI/Gog9pHBNafP07Un3J/IHvQqp0xTBYA5f9QfU5v
X58cQw/9Nozw04fKu8CNwRyF6o92qoEUIxDdatbOX8zmF4o9k3Co+rPTbeYPxOnf
LB400RPUpNmxzGaNbR32M8psUy6eamm5il87/ErdgF97bOo5x1ZrLinJpk/t/6XA
paJffu/J1OKlhLk9kREXueBfQ358HJlYcZQ29G7jXWAEqGRTnIAwGFAvmCe3C5eO
aItF06diaDdEx1QnqPQ+aZ2GbdmaVfW1EOhjSiXuzOI04+4AojhYhMbiLjMtM6rm
UePk7Jy2dUghuJqPND6r51XOuZjlGmoR+P1qHKLHMbNae6DZX8Hbv5utx1NW/z8t
uBE++YecJJLsKpBMQFoHQvgCquHauLr4UyBIt57tSg8B0ebz1qUL8weX13TFINvP
6Zb4jFQPXbJjvdVHqf2hH8nkkl1Zi1tljquHsBoAYLPM/JvixfWYLmosbzlpGFOi
BCDc/TfGtxWgoRzgWdjqm7zH916sGzOf6dx8v8cUth5OagOveb8QyLSOIBPy0yzV
rjkpGPr1Q/acBfOC2RCyB00Gtt/ZSowJaq5hmv1yIK1KuJPE+LrCJ9GieL++Q6yG
g1qLrd1ibuUA0Or3dlIMVZHB1aKKv3RfJ6tQhw74ATLhPuXt3qz44XEejQ6NM9Cn
8HW/DR6qeXWYRs28jOMaCq/mDTlWL504+MOX1h/kEaQY6jSNCDpCJaWRuTpd1qMk
m29etH6I/UcTuwy4JAhsKvxu/ymHJxxzErnRqCSVZM0XD4i8GcBvMhyYqZtcSqJ5
8y1RuVrZ0k58RRODmaddCRHIis28SnlFTeFwzFxgpci7FvYfQkZdpKaDyXAFT0iG
NsUjmJ9riz8WAy4Wrs7x8CK/vDW3Mkienz3MQlXB5PJuj4IyKdvW+hg16M8PEY78
0lFa/DSH/TnB9QDzQALPtbq0l1nemN4j+28ME7WYohIadLgTF30hcsAMw6iyIWhD
RyI3ICaX8mZVWpWJSQevf3IXMKwM7c2HEVQYJGkeu663Wxhd83iM+dJFHXSd+Wvg
4eXcVAVeaq+r1zgyE84YpUCIJ2ijmZ2YetMeL0WNPclkgC8594xHVZKyhBiIO4TA
np+VHZcMsUlFRORYkPZZPdauSEtfE2mKGk+U+IQ5j1BGdviBGZQPrgFjet37GxDu
GiW+y1Z3H2DhyloC8Zmmx1N2AUXj+gQydKgl80KuNvfWOYrmWlh/nzlYBd5T7rnV
t8bgdnn3CSg/mcmwkgLrcUB5vdOHTX8KHVyW7G71xurLcF9iAdhhSquDkmpH+Sew
S3R+T/ViTmLseUPgGIwLJDT9UOu03I256vaq9In+NAsidpejdrvQrctaIEcn392l
gV8tRoJjd4Hrqbsuyv9uwxPA+vm/m7XeyvI3cGcRMSwxuYLwu+gxFZdC61Gd7+5R
eUxnPYSUU5ehzsbIk81xai1G/zHZhYyf5rjxZBQgJpgtMkrqhaHIQSMjgjjK3zx2
KuHiMJiggps0NV4m4Ehk5FiTnXHxh3OoliE0l0b777JeeMLMC2/EpbEPwXLJ3ZZ4
T7YrtlrQ0q+kcC5wk7RK14wvEn0U2FzMg4eAnI94faLh64EFBGjYultnrySC72bB
W7jHehmPv1HV+Ygego3R9qy5fuUo5M8sIDHoZGZTGQTP+meWezsKwECWGBgm3cxj
sj1Y2642Qqqebtn000/cn+dKd2WkhyKpQbStMoTQfUl60/fvevtV23y9oEeIHcpS
xWFddHkYwlqVKtb0UoAvb+CNCtvWLoFzB+Osi4O76OQWYzEPw5nj6FLC4oGia7Kb
tKunLpEZdHzh5LhwgMXLIDeUMoYAmWflBGPsZFJD0osTiY00bs7Sg0I2cwVUIQyz
LC45ZuKErPXPLlBLm5V3NTWKIlgF4Ohu+5g8lFpNm/ER1K4/axD27pLcTvCCROdE
f/K18cBija3Ehbyz580wiDpGbTZF6liE8cWfQDJ0+8cfyeCnfuqABIeS6Xv0Hpwl
SOjwiAm1MUWa4/NusSwtrG6/+rbo2E1XfDiGJWFo21x+MLqlZiT5NWgtelou6Auk
MTbCfAqK3qFO3+ytZJ3i8AOU882Z/ZoefIdBsfMUECEp+bNrqTvEZzWuCEKMg78M
bWeCjFB1zr2iz7Bo0j1pGUiCJqxIs7SwcXf+qsOjxW7WrnouUiCd2kWr71qy8omt
CyunoBpOVBcdJrTpsGH0kyCEpW4fX8Bu1t4/g+lwRQJbJ8kDAtCMYws98gGfQPhB
aThMXn0+VKtg2Xyqlf7e8zsaxF9EfjIZfEgI36KQEAJrRm63LrqOZUGuyVQZJSIf
2a+r0vo3eaFQ/VvWn/4lQSEdtRmWvZRmgXGYfwxwzN2sG1KDXU96lT2SMeCqP5n/
VrbD3cToK0+KupTSOA41819UiZRXfzoHvEEtoi9xSi0BJWJ2UuyVCZWelFv7OLQS
aqAZeId/IG7Q9XdzJpHiXwNTRVypbplXJFO0PIuO+5+B6asbvbqSwo3xsDE78eYZ
PwNYs7xAZoDnj+hvs6ZME4/IN8T2E4qboBklq7eTfl5+PI4qlntzp6HK6DcAbTVT
mMGr3SSQT+QZRFCG9Uftai90SLfic9eTJTgkDI6EC8Y3MS3jsIZeWE2wfUlnZGkJ
jdbuxoaNbOx2/aZAsOOlNk08ow7HtUtCcQZ2duEKo0H+YYGupwskgv1KVnZIUOe7
+Bkorl2ugOgkdki+mvEboAMsqIeqJbcN41p/EibN6Brtx5vmLORTabMt4AdzQMZX
lddSzSNDy16UxdyqbmZALTti/Cntl57pWI6sg1YYR4fqwAVbVsnDLAaBSp69V+fq
qo2RkGZ5sxxtRHkNPhoeLA23JaI1qP1/Edj2eN3AJtd1dXxFFjDmyDkR3/kpwZgn
XooJOw+5gypCrLGfBu0/dMdaiAnLixf75gnc3VjhvGQLYUo1/oKLS8m1Z0USvX0k
1DAF3BQoRZDUfMQUUbb/XDHz2vwRiWW+B7I85f5nmpweRgxlZrnZqJk3jcGoddi8
syKZt62yPDAOy13L15jmU3DhBuDWxYd9f7dOhcgGG6Bd6OFSbEThdHDP0JC8RU+y
q2UsOp+XwJ1fZrfH3+v4+7syu3o8lCygzWhvAs1y3ptwdpxACr1eeTk45nL4mWNb
QOHvJy4Fo5bz1d5sIKqjehAnMZKxg1cz9GFI3ovXMhX5WvxjoqVpWaWHqHQF5ztH
ruf6he2pwAbprXVD9H59zgJYBufzAVRuCk+gpPqOD2+IY1zn1S5nwI9Dxc6RG5Ne
DitKAzX2uxckvo/jICSdXUpfXP+SsVdupm9jGiaQT5eA7YVT683JvUII+bysV8nN
DsorUF6WJYsipFFJ1qI4wS6kq1elnGuCbitvYUkbtz4a0kwYnACE6p0cJ41+DFUC
GCyI4Rta6qLHhr9X2zaj/w4zQSwIH2BzhMtBEJKGNKo9X3uSc/KKQHFgxG7kJrhA
ZdqVH9n4QHvkIVuin2sNmbgztnkTv52yf2mPxZWeonptXY6jMofR10qFpSs/PdOJ
XIbS09DqEmuA8DUxWVjFO7MpwaCT22Avuoz3Bf7y1b811FDjbvS2b47XscisSNHB
x1SvKTZHSKNe5CHDPweQhMwkx15yXcezuh8tHjldOP+ayHxSQwzykxcFLAuibYCu
AL0aeOS1pwOm1QvN90ekSpcIhkeYsssiLqeaoCH/KiJLFskiN6Oh0CvjR2zK2EEs
XXVGW68VlLKfTU075hZrSsJHnbXJGRMeZrUI5MtGl6kv5mxZQGx0NBoTd/NyzGUh
DrIRTlJozIBO5Fe/uyTHm6FWiLQ2IoOaNRPMuEahJHTPnajBbYqDawlWImCfZFB5
k981pI5RKNMpR5QgY4mjGVuw+5wkbGvhocdKFA+S0pAO/Y09aNv7Ap7kgHPL9qJu
vePpfgdB2tPCY2dZs+tb8KNTNRkLTiiP5wLnKfXBx/OzBxX9cuy3HNObuF976ZgJ
0lbLiW/g9voE4nYLJE04YciQ4ubAHKrOsrova+avoXIdCeqAUphryD7HN9Z6ThYo
Ck8hS/qfLujn6NGUHS/fgXgA+BJGQU7AcUsmRiH9KP0Ob5Eh715CNiOfE+B0r0FP
qUHBSxoMsqFKBpuDpvPoEEovPPjKkwmf9VZ+9jwXu0ASOvuKa18B0ssBnZq71XuQ
aFzmeOOJx16SAGK31S7uwF8IYVaF4PusOQ2KOYbqWpknOVF8KF46GpjcvnCvHJ8s
RhVtMo5QmdhEIx+b4Fy2zOm2+xsOf/mdIyhVqUG/v1bEO9N06Nhs4+vfhZ5sXdLj
gFEJ/Sn+0YtXR5lYNaTczGp/pKQDXO9i3weAXT6NcSUR7Hb6BJXF3VHHTMkXHUtP
EPKQQ9jOO4dWdC65dm5tKfqHVizt6WD99N3A4qrjPlFZCaL+BKaIWiaHVLhmZnm4
c2T3a7tX8JQmjRPTnCugzFY1KL3kczWoMWBUDL2Hvw/WCjK2TtcjpPnFW/NpchGJ
F27EHU1Aysycr17iGhxhm+AMrJ57TVcXm0588Dtl8TEFRP+myrZGn1ClEcBhEIps
/LCne2vdC4NycryKzcnzLl5K9qPTpHp5W75bHQrAGg45yCfP4C+lEQLeTPeWeRMp
w07SU6q2SFaL/1Z1q/ab1VWNO6r6NlRHDkM263r9V/+FnMOrhNoN3QXLofXl2Og5
0+WemMOOHUFBK/VAggY1zd3yZze8wGScYTJBQlC8bZ0zWoP1/CZNxP8OCsaq3GGf
auG8bUiod15LTFmsKOegMWIZqY8Uyy+BiAO594re7cMVwsR5oNIq3ObZUEWNJRU3
WuMnrqzxOfFlSSJoStimGIOJudkTBWoqZtRAjX1NXmuf0B2hU5F87y041D1sP+kH
C2/LWO79wgjJ46rmydaBXlU/H/iLt6Eqo0U3jXHNtXUB7+9kz0/rWV4T+TM+7G5b
QHJ5PaeIdq/ns8A0tF30UhM0s0VewV5TBxo4nFc5BVY5OBjxkWWkWMR7ob4gAJgk
P+QcZEnnE7QGii43wpJz5t35s/klSCKt2tyQRIy3R/VgyAHY24j7KLjGA1Zt4TCd
Ney3er1TVIpUv7dlzz83Y8xFw3TWHHjGoYbprf9Fc/UCQaWHfXg8sFykL2VwS0H3
Bqqz0u/Red1GUy9mc39qsVB+NkuGIo2352KdDeiEwtgciulCii9FvV4wwWTr99A+
zIz5Ku56zhmcRk3XVrlcHIbnKYqXJLMbSJnXbrF3IScTQ8s8qhJvQst0A8gZ2Sqk
ABlQdP30CVU2ZcxOJg3D0MUw/kFpRSChfEty4uldf1fTOjHzou2ySjBHwgUK07/O
tPM8Hu3LfsK1nU6V+QsB8ejamibdQC1xcU/L1J1Ea1VfX+jeNlwfGZRcQBUVEVEE
srOGfCwRSKZXZlP7GN8B9lHR0HbwfQRWnhWWPINLlMSZ+7xmKx3Dd4IURidAJKfi
/1SZ+qDDxgrEtsCqIxC4zhljzRu5Mmopf1mDl/6BwQ3itBY+BKFUoFdwk8d0BbDi
QFMkYKDm6fk12YzyUP8TvsLa0TQRHXhEbX+jrnkEZzmGIPBXmuhpP3GSOEgF0GvA
1TwoIYQb24tji8lStyBTa566WzWy4TuKKrDLP3r3Rla8i+lCiWDsToabtgzmGBNc
eCeDNSPRjkYTXlV1Ka44aHn6aNnsy2Rk58Hp2bOQO1P6yMzVV4Fk/7ZAij+m/+xX
6fKFNSh3EmJVLSLGrcuYet0usbwqT7rkTQEfKVYuAV6RHDdBKal4eyfly8X3b2BT
j3qNHCKSa/vZUyu+1k1o/keerVmD6jD25BGzxq6jBN2JhKdD0eTQ/OaLSnnIWGy9
MI9kpEEuzvCTcttYx3N7OZ65RKDDpPYouzgrBtoeUx/0BOrNOgcjWMudGjhz+x9P
kyrh1WwRocLN4sG//eM7n637pikNacO4fEL2qYPMDcPG2j7HqoIbUl1TxZvczWRB
NCLOyTdoaNfKBYh/VejVm+VL6pOl77kSGiBcmydtfS4e7UIIK7P074RtNM/67tEV
SA+HG5Lofh7sp7caxpJQnI4Q6OIAD0lKYDinPnpUJ6bHTG3VaLBMcu5otsa+xhBI
Wsu61xzX0s9CJ9do+2N6pcoLtpQMBHiOlDtGT7l1Aei5/lRFsaOVuk9bfU+rinsZ
k3ot1UZpKOAkn1B35V2AMVYDS73ajUpmJkrJjUoRIwHDfd2t/3SFnNGj1B/KSIZK
8v6ODBZ33nvI8uXaR7La5mowB8fbNlnSCLQEK5My+3BeCfA0lOI4R9AlzoQcNAX1
W76BGFQxBX5DyTu29VVWm8UQ671rjx6rgj/h7zIxpLFDYhAUFH/hRfazJ10BHhFR
IUNyKjIUdfEjcDZmo3cHBG8JPOwCn5kKFNQjHrFxjq4SqPdmrbgUMpCdAlcd/oa1
Ni0Oq/d6Sk/B6/rks6p3PnXjmEaxK73cdOFJDk0eCpsWqGvK6yzoC1f4RPW3BWVo
EPtVHblsxK4vXLmpZkanMfr8FQ6r7nnK0lCaUFCyRBVyhDQhjmoxOoO0a3K/slAT
gqp4c2H1kI0NGpjiGTcbvcQz0tT/Ett4Tnghh+Nc+fu4ZESgmTru3jj6gvmUp1F+
558OanfOeiVa4kcVv4HuptejDRqOhAW/FM8DhL5kcHL7gyu0YrcUrDwHOZv7pwad
jmUk4cBQUhogTDeV8kW9asrR9Y476MqDqDse411CZNf4Q/63Y0e57+W7PGhv8NFT
QPyLYgoGoGrIbhUVhBFXYj1S4kSw5bJ7Ax2B22tGRrF7wNnwPXPezb0zEYYvRYEV
UhQwrMuFCQsi6hAi/dv9wR6Ma9dOEKdwbgxPi5wZGIu1HP01vZ52zrGz71w4+1Kt
iyY+Dwuk+MZKs0Hy+ur0cjx6irxSvHcfw0RwVGfup6rd/SnzYSi9MjawgbuTPdzc
fVQ6y5jfwG94ebaCkM6IQP7gQ5Mq/JhdGSGnR3Fit1uZahjotwjto/Uaft05C5SV
wMcb8/53Aj2xUM33T/x9hQPu2Coj8AS1yI5CBOLnc/8J0QtmaGAsLfpz9q2vfyek
Sljub/8/EG/RFoEoD0yh7DUcOuZiZNvnvIPHUr0UcNDQI4OPIjoZYATw//fjL91T
a2GZvoDGtbtobyjwmzFJCugk9xct0VFhPgXaZu10GWsfSOZeVobnPQPqUsUt5tSy
jNA+oiL/P52w6Oi2fpxMCIKGajVYIUhkmqZDL54qrofMRJTg92bENAb/RCjaOQUO
766PfqnmQwbiSUMo+88X/BVswrVTtB70r+kCoBHVSCnwKOSvOUUzJ3NHiXVAXtgx
idaBj31W0n11CpSNjOfryiQUumB9ZfftfiVfQjBYZPQyf5J47t88lxXyXst7aqls
B6mDKGNXFGRyYjKFjU1P7WgnRL7OvJm6QrOT8Wv02BEhVjP6nh3rMbET3gl/kU6A
IZPTLkYGqpopC8u1xwcFeleqqYkSBScBnfup1ltWyeMAZxqWJPZFEE8lstKnV0aG
PGKx9H434oY3j+3wugbJQLPza0n064CZu3VOIrlPQrVwXnW3AFCqCZnMgyfQ3RCh
Hp/B5IoYnp+GzcUYOLueB6BSfhkh4xcXrwCOIdp6appmYL25SRW8Vk3OVuobPJK5
UvJeKxqZug8yLf31oyE5gJiiAYeqabU1+xHwfC89zO6J4QHLxzQEZ483gyGhEHmY
+/nUvTUOwZMIsdTa61RqqOu5S2OKMD8gFA/0g8THK4h9Lw6k3ZgdBMaAPxCa9hD9
MH78V3zjx8u+BwWzQbrugO0XjnTiz1fD0qPL6W29IfOIlyJc05G3uJogFdN1LLfO
T4zyYptb/Y4OvFY6nqmJHEEh0iIdlG8tRCFmmN1pQGm5QSKWBxnyEDfNsBaboeoi
pUCD31EMCk5/gN2ICYZ4Q9X0IDM5wGMc4wdwwCoXy+lVoA4ltB6PNKtmoH37o25Y
godZJUwK8Px31zIHczBsYKu//BJfeGfuGLOZhyqmQkNSDtEo1Exhae2eGAQr2FjF
cn6KlB7lk4MojRxS8wjaSt44Dzpz5+zZZlyywuwPzVEZC0y6418vmE/YgcSjnkJ2
ea4IcMsJnbM9WOBpDl1FkEuYVo4KP7RLbmOyM8dDc7/mSLvsIU2zxwQ2GSXGkZ1Q
HAwp2mgOeakgYffQPGmYntGzthn/Tcu5fQf8qbX/Zesc5omA3Jx2Crsj8iU0+bk+
hDu1EdL7PmtevpDN+S3/qqsEHQre1P5kpy2qRTD7NwECCfZiSJc8hTF0tbdXE2F+
YKt83+0NAoS8ditW6oKMlVBxCofAiUHX8ag5neERcRDDeV+SyB+ByZsrYAWlmkbA
MJ0QwST+Rxz8ky2nHiQtIFgMr1Wpz9cuKgNqGkdB7w1ylPJMeHGOTeO3Tbhy0RBJ
xjB+H7cJ9jKmiH9DsU17uJfmWARf58nO/QLAnWK3JHQncR+NHolpO7HPGLdsnpoz
Kut/EuSW+GI/N3vHPXcvma9fGZS0Osw6PCsD0I2h9mF2rXoK0Gtj2yFOkd0xK9F7
RAATAAsY6M7sord5VwsJ38oVBFHtbxXtcgrgAbKchXlrhOEcTy1pByhiS8vtIHCE
cXr0OplyQpYLKXRZNasqw5eengy55F/q82du5lySstcTmP3+YV4Jzmge+afSoXZP
nv5+o6kj3mJr38Ceb3RbaoytIAkynCx3+dpiVXNtiImhKUxpaAwDSXlKwyDx93y5
twXQphEQ7NCJqoTwIwxEerhggYvaEDxF4UH3Lm3y8qqQlI8gKH1hI83qs1Qh8HhV
XcdTQ34e8mSV+rcG5hdUrsZWHAe5Zaa8sToaCpvgCxvKdx2THveDsccAV1zTtD+B
1fGia+2IAGqY4pyNQuFmpcABttdO5JfW/wPy2+GMV7izf8+2kgUOggFR5StrpYAs
6Kka/IZmzqRLwmP9ctMpGh7lJK99g5qqvALwBxybiJxZAvBZiyHIT4pt4flfQxpa
MPP6DmcAYf639DwcK2GroEb9QAcyFciNWD9b4+Aq691GkcSNKwEcvob+2OS0ofn0
y+osBA/MklHAe4hu9Eim4OkES5Jw5MqjvhKVZHHWcaRLsbXciIG0W302W0S78Yky
TIlNiatDgDQJ/RzJYE/vH8Bkbr++sziGnQh7doaCQW44lrpxO6Ik8uqAgxNK5NVK
426dMN+z96ho7VupfN0ihKVeEi87ECYeybBB6CCuH1eQp2sLYNDTNsHfUL3i+G9+
GC5dEJDvQAtXoGJVYIC6K82VNDXFuAFKP3lJGtZk5k/lgDvKI38MQYRUsCF4fknH
HgE4tEyWhMqxVDAFU/jBex4Hgs6Hp/IsPTHQwv2UoRKy+HKOwFwt0CkVW09Tqx+h
nX6qjj9sy2O/+HqDxdWlpoheH1jjjb1pfTxi0+XTfn8GJGke3ctv7ztTAWRHp9gn
UUyTJXyA85f//3aeKMxxuF/9oEEVpNQuVmfa6aDhcdgT2SYG+0rBrQ8P9q9y+5O/
vRnMUemKMtXmqo+jfzgbQlbSe0K7UxpbJA8BlI4+pjywbj8Ab10+IgEtNwNlDpk/
DtsKCztSiSuHNXomE5d2ZTqpFoIsyAlczVcNSEyqTHudk8yafoWT/uwqV0R42r0a
2PXm0u2ISf5hepGVJBgxknSH9UBVkwtFQCYKggBomvcJZTUW+Cixf6snRbskb/9A
1NZ+P9Rriz9GHZPbZlarfMpKh0jSaX6w6sdg2h9XhBJ0yFyefAO2ruFiFZjLbs7B
5LuG6x68Uhy87hC8pecIi+RBeCEribxowvXlna1WMIymzN4juqIBeQ7K0F26pZKz
md9tk68poZx2DxwbukPepgQPVHmoL8QPC9vBBuKFIMIRnsBCgew0B/bizXxUXO0P
06ABudGTh6ckbV5T3zwNj46Isv7KqkvGPYf0Y8nvmh5QTWi3pOWgcla3j9Zw5dWM
u8SNt8IKBQ6RpuPhQ6NSY5Uiq/7tIlrOq8vdLDmHogfeKmbkB/0TaBh/2YQHjKeP
sNyawUeqtdIpvzQ8K2coKZUwN2mYQ7j7WUkIdmR9KuDml9POiqUoAvxHVi9d+rr8
9WLzZUoiPtGI5/R1PeWxAPuLtj7cPlWjbRhdvTtQ1tGY8+xJ/dZEj3o57AsVMoXg
jReuvuVTNgVJsdZtyq7Z+JbARBX7gr1fZN3M2pBKyLQJuJX2knZpa29qlH/0juDz
1LMriu1gs69vmSmTb5QKLzGA7QMXjPlg4YmknXCQJ7zJmAOH1Aw25x1p3gz340YI
bG5uRVXJmlS1ICeA4g8PrV/RqI6o9rGuh0uvh8luhbUP6EnaQX9BZb4Vx/8GGlKX
QDHyjVZtroqHUT4ckGpva9/KUY4xOStTh4fXzXXPoQ/DAPz4Tb6hkNA7Rr6XJwQP
AKqytFK4M3O/zHtTgm7tSUnHrSzn60dH7mQLN0MyfpYuMvKa99RUZkO567xIOfm6
8byj5OpDiKNaiFYDQbBOirXLxAOv/ePdadrgGbDjXb23xq6gItORYRaEr2VRjohq
FdMlDkshufbBaPPCwombhW4Tq4vh7PmIPZTKjSYYyDTi3xtCwg685CU6QxWPLzI0
AuGvGx7G7orEDb4dxpyRwZMlhpvlDOFDKOswtUxx8lTMY53uLz7VSXqLwu60ZcR1
aRXZGIQhStu0bgnbDmqoUp202Jz0iZ0kea5+DocHkh5sEI1ZNIuzHk3fgPTdYUVI
lko367t54lakomO2dQQaxowrODrO9ipSu8fFUfMPEAH5irHX/n4XUN3YtpGFt7SG
pflF1bmf/LgI7wsMAHBBipSTpG2UBVx4wTQkT7SSKazh5OXgRF0OxDEw3LC06q8+
MxHSlUDSC6Dn/hI1hESGLSmolcwDGMfk1yTiFt5d+xYF1bL3587izICE99c9IzFn
bZjLK6pWJRh9iUcn9b4ECDpfPDCKdnsdZoG1szUgBkCq8/ehxrAkgBzXIjGvYZad
cdCzGbM97ti5Ynnc92v2jOMXeQK+Ia5fyurvau6ioHnqtZ3h/97jwkritoNtOL+g
0mpNag5LzvtEDNZ3f9B2C5FjxREiXYzQoVjUTbgIgEnxheBDOx0PJKW1kEio3ukL
PU4VRZFNtWwJs4jNiy6HaWGzTosqmB9JXKN+g6+euLe9tBwNE7cl3s42qmakEYy3
iNlJD1QVjnEihjb8n3xCChj/4vLOrEens0M06UZY026dqb6pgEw4f8mcMvovYE+s
eaZYieEksC8oLlbg4/Ctd3awFQ9b3NGBqJ3J9gCRdLOLCraEsXMewOtup5ZqTuSA
lZIP4Zox4abtwc799yG4qt1f+hnGvCBO/pVryLETpnE604aFsEftztsvmNPsekk2
/M4OQ9j5eafp28B564TBFInPhFeM3ytG8UdkGVhw5Z5upL1fW3blVBnHRF8QwkKA
8YUH0k+dYBlVd1rU008sJi3xmKUziPfi9wHlPyY12gT7F3pKe/Z8p6vU7/2nU/3m
s9T7zNEU8dZ1R22DG1RgQsLVYbsKLw56OXMmY3zBgSF/bWFNlfAOlwgfvpLeCs8h
/G+2TUEHvVj7AEo5Fm7IgsX0hcrFB3dbfmpmaYPUZvirUFPtg+YBc/TpUsDf/7cz
MNW32+VHrzLZefOqVK2r1XXRFcn0vYinCa4By13vkqHzhrqqFyj83xbPP3DdHD3g
JJrEKT9W3JztF8yA4BtHvXaXqud3NhXLyrHk3XwHveEkHPiVX/7z6V3bfdJwpp+D
qpLpxoxIf/fBmTB41QEReMI1ezF9FtinaT3ow8ZMzRogcVqVteCZKh9RWBhzggl2
xLrl2MJ6ELcH7ooHT8EW42RcH5VAJJPUM5dAYIFdOEJCKKW+XJ4tFlRI15+3mO8t
Nnj9qv2OzgN4A92/b6mAhqK3tEUveU71ytY0UOV7vFMnGgXtq3b4fjHuU5np3jt2
DGv1LMw3piIgvfxsE5A9gViF85+1zHvz1dBm7q2aE7bwbZ9pQVYLa/eeuogFMwpu
5Xk2BqDqpqq5S0yrEzgefy65W2LshIckNsYAqNww9V7uC7d+4rzJtt4IZ0XzNO0/
bOpD5DJ/tKA+GOa41GUKuuXCtdKwQJbcjzE9rgXfT1qPCU/Cy4wK2NU7N8dkd7Zj
sMLvn1mh+YIZNLkNCnewdcOVge3AlVQVPPqL42ABIh53ln1LKEjDX6hvSnPXdZLN
yFVeQL4iyHgP9DyCf0Y+TV9EYuvZSZ/vplKpkvLyG/ZJinyMzD5wIoMJ+yp8uxp9
cZDJ2jz/iJVkoFth93lImvXC2OjJIZlpufMT7W0sS3j7LNQ1XxWQRO9ScN6BxZ8z
FM5u3OfII2L6r2QTTgmwwRlOS6EnnCosjJWLEDXzzmv8SAB+JfGg/myD5hkPFtwN
rT6krvKAyDCCjKB0Kt8+YTS0ao9eTRPGeM1XAJ9EUOL7vGbZ1k8ucXKrQSpDDEd5
Pdnti51fPAikaASPrZrNkEO2b4n8IiL9g6UNrgvvnZ/Q67kIEUlTRCCQOWDBkz9D
rM4smv3EgaqPqrY14TpLpS8+qsulcPcXlAh1aGcZAf4eqBuLLIdMlxMxWnF7keqN
ROSNfUX3F/1+d4BU8+kkhiZ4iEfGZ3CkC7MdJJxO8ru0IGpfk2lXozqZl+mZJXhE
KBoj/yo/EeeqFgUAuvVITxWPTZ2rAeEJ3otFvJIB1Cu9RJZbaFDu/dK5cGPDTn6L
m912G4YOtH3LspiErTCufOMMLFp30G3Kt7jAO6aft3Jk0Z4q36dZUoKfQKLWLFiC
qnhMKrJqIRHrs6/zMCspW0degslvP3k/Pw7Q3vL4pK+fBkXFju4tJvxskcyuTKP5
7MuzzNwG7kRNZHy1jttkuQ/9XBdLbTVcoTmdzyJV5IoTcd2vIG3iIeiIbHmqSImN
O1lJb//mIOiHysVuNiDeGN5WuaRvq2/uJPIE8cKm/9Xs5UwgAySt+NbhdEgwQiEy
zkaLOSJfpeThqjHbh/XnUb9mzHAzaMm3XgJKcddTkHgCuaq0WWOvBRg7DHSvH/VU
Ybq1oOlzk0+s2ZgqT23yqygB/rQUnK1EIHGXOBcT23ULoXsiOUg7iC5NFXYmbZdD
0xSBpEhvOcWLmFl00BXm5gkBuoyTX1nJ5XZvWLiYxhSZBeFKVh6K0hFusXrTLcCR
V9vAbfDl04S3iM/KbMZcV/vxgxqMoS0oLClb5Bs7YYs06l6yyA1Yr4bMhv1Sp9xE
+7q4XgGn02nWT1DOn9Z+dPFQHaWfKdm0eYKt97oApo/tb9eVpTn+9C5I0eLFTWBr
lhAjcxXiNkSHtWUmWGlbOW7KCgk159/ScG6uw756u36pd4COvwnOvikLbRlT8uA3
fs3xPcHkpG5LZOF4s/iHUePwFsOA+MUwJb9VPoUTuvUMvJ2hKqofLPEXL10MwKpP
L6qfCuPbA2uvMEeEN7O4hwbDWdsl4MTu1mTdDlnrr71S7LXayo9ZdNU2CWiAt6vI
ZlFEQpIEasuBbJTNybHVv/yxBQhfm0+XBuBnhDcoDYrXoSTvV/5O9idBovgaI82p
NM3wlhnfKTkaCLt/FLluH+BPLhKnj7xvA1gay5s0t1AsWOry1lDKVjwE+XGzq6iO
w0bvm5CQEaStlec2Abno7ASPFA05dLrEah2ygoJV7XKgtva+qdKldna2Tra4YWKI
xe8EQ+RpP0i9jZh9YHh+6b2Ix3KXLD6OYAJmVF7GztE2rBQ4aa2K7GrSUfipMGvj
hKzgZDr8kvWkkyXPO68NiUpyX8r7rTGe0pohHR3oLPu08lfHdhUamg+Xf//UiFHk
SRNPzdFAbQn+4s9BIGZb7R1GAKvo8dD77VvHTUhwHQvwsfNYzXmfy3U/v/OE2uq6
oIaAU63BSlacRg5VjPGM5/DF4LqWCiNgFKPSmPOEJZFVaopjN7NNIouLOKEDJ9s5
3E6iRX0n5AkEHyAlVT1UJZvUw7OemnTr1F05UFEqubUTZgYht/kXy4AspNqIUaTh
xSVnEgpiD5Trjq+rKrpV5hFHWQ6jPpnBWaXeqGzuosvJS85GjwZ5XZ9wzLTCiEZl
FU1QCGKbX/ubOmboAQ+21iYv2+H6na+8kodilj5xRhQS7FDbfoakpltSQyMyR9GK
UpHPLHj+tORAjKK8Z+ER9BQH279fsK7C9coS5zsy8uaWDenTuJVx7dWUi+W9E216
o/oe4I+FFy8TSDSEfOTSpWcIKlyH4sHchMqW74WDoaXtH4jsLZkWWj/AW+vveslT
MqBttsU8Z+4Bf8fSogbwrEsdogC3BNS3KHfxBX/g8Zce7zrzXjD1gHQu4LRgGRUz
o38jm1oniINytHXyQljaGmGUUYvSKL6t8mskbbebkcE8IWKh8lEUatS7s+OxgMrc
Rk9VFJAQhpPW/EL8gMfd63dXkmiGEpjEZ/PJnLXxhYftBYdHe8uuNtWGrQ6TqeRs
K1ij9J10JGt1Xn5JDZTgRjFVB3ITYzNu5HiM/QSQWK5H+zrGFU4tEuFixVEzi37w
LFGdsAvx5/RjNfENMZaMZAyV35Y9xNrSD6r+n2jgCCYeebHhPpSE+H3/7yrQR7Lu
ADcX9LybbI4oX2IVAhiM1vCj+9gUUgpkVg6icg31Hwqrs+zAAAREF2NUQ7sRDSpe
BSIgx5CgXRahNG8AeBiKTjl67x8QylBCRtDYJfWqZv3zvK3ugbdY+LmMMSJoujV7
OkMX+Dkn0A5VOcYTajA1KM41S+suhrecJtyfXPD+PfvrWUpPgqXBnJjL4lVTPKom
t/a2+7ux4wr0x/DKLMshoCqdJXVf0+3asuGE0WgurtzAkiFjqWb2nSnwV81LHkLO
32hDycSblTQaVJs421LsJx8qDuV6kB2z0bnh20/M/vk4VWdEmNMbWuRxwd7S0OmZ
ICPLFaTowQmy/j70BUggmS+2pKf8FcislovKpC47X60VeGl44I4c8D3lcihwccpA
hSQy7UL+GILIPyPjUnD4XUjUGqlSBSM6mhYBO/e0D4KArSwXn6bc8AGsMT4/JrBH
y7SwGAFBwpdaoaqV69G0OS14KrW3AMU7ONkeXFoKYmK/ynHPrVUHgxvXhmLIFYOr
8HR+4f+8n36IO/mbzH+EUZMUwx2F/vsqbZJjfID4v2empn9I+1gQJ/4Vo9UZk/LP
/L1pdv2LG5EfonSX3rlOWDn62gtU2o3sDsmIy7QvqzEpdwt64GRsoU+mW1dSy69a
wJWPtG1l0o5bgpCTGNdNuy4MACoA5XJRnIjI8DnsxGv/RFjxLWZOdSeDVl4zcEMn
L1PY3FiPqqB7EGB6qn5AFTDjc2VghooGWY/P9Ue9/L+nAJrQUtxduKn89qP2f8+T
RF3KYHr2JgW0mx+N2ThdkvxmSSJG0d97AZC5WobS1DQo3bVzgqZZaxKMm2QnWruY
6JNeX/t2lxX9fc67EKINb88hTHs4RGTvLycHGunhnf+zh1YI5DlWItAe9+k4KsP8
Qw+uFEuBqpVUAevaHSGzIXTXE5WKDWVy3McLilFJ7RcZkUT7rX5yIgvcjdhH8VtS
QbVZr8HXNOD79/iktuEbp65x2IvqN28zlzcWVN0DRUk28Ul0kxc8bHqR5N5JfEge
Lg+eM1FkYxsKw+IOvefq1vVAOrPI4s9jk3zhusSzT8FusrYwMWrMT0cCykwclgQl
TVgRaL35hkHr8KHq0dXIlfCrjER8FQ45KYU3yEbwmf6Un9EbDMboeiiIu2Qzo+57
jz+EUJRAWCDt5ciSPkh4I2qnRXgk1FVCOt25rOIzrNgx16+uz2bDvmZtJkbG3RX8
WAXR4ksWYfEYGltzilB1G2Yagx2LZe+fo3HX4ajQ0ndny0RwNHA0qomkAOJEzHS2
6IRRFHH3k8IhH2q/5Ki7VLB7FkiabMlQJx/DdG4hnq8q0Nqhstoy2YH/gYeNztGf
sp/rJopJ+w+UG4/Fe5fwAAo2BciXXHpW2y4cLFXm6ErGUPFC78tDQTBtpPyccmwl
yNF1yf4fN+Vkms4AYsqdkGzDNe0A5NeyXSkHLZArKTrrHYkm1f7KwTz1c1b7QFTe
cU01bu0rif+cRrA+XUi1bEzonP3DMEskEocBpkR3dPax6kTjRgNsYHvJbJrl1qGw
hQcKw1TfhfbWpRylwJevhyBZHGhPCr2q4G5+H8BfedrD79u5IxIEEJm8HzZIkp72
ceh3GDsiyw2UStEcp+P81jCfPNT3y1wue+r3E/aln8xUC9drNg8fuvhSMRr2uqxP
4QshephCJJWxqe1gfCIveADCRtHs9DrLvwZha7SIsWC+b0p4jFxYFCVmulUmsC18
EX/poZkn5mzQ7P4GZJxqFBZllTEiqpJpUVWYKkmDPv8RdualwBU018nKKyKWFwiX
Vjghl4ByLU7k2/WpPUF+Xr+bOi8oQKM7s82eqvDAcQxFK8TpIV0FSVWGM+72MqIW
jIG++BaGM23O4JqAUIBxN1uOQ00sGJ6nrcNGFDFVnDn+U+7iZFrSZCbJD1wLBWX7
tSoiT6OuUw8j5aIb9OTfX45HOvogB60dcoKlLv9ukwHgcdxX01i/P8jVO1obXi/k
7jA3LjuoMeUEslMZjpFuWrF5CEe0Cf3Hyx0glFuTEglDCEHP93JukXLoTTa7EnEZ
Dvb8jg1PzJjEzZzMFKJGDMvNbfF7cXJS+GylpHn80YX8176QMiuY9BdotuFQsymo
eucykWjLOYQejmX3Up8IWHMDJ/hkohu9IsuDedHj2GO9k6xcpHiL8fcqPpfbtms5
wUUNWxrLyeOAYYrL8CBoq4Wav8pWaphUyjOJtNtCtaqb3awg7OxpS3B87BupOCGM
uKZauuxtAIsIz6yQVKoQuQO+NeK+eFH1Iq5F8s6+dqBV4PGdDUCmXLN+w33tKJuj
L0zbq4hLyn3xu1rj2b/ujAkxL53CMx2Z5LDu/UgxlGzc/h1gRNWPWX8G840B8PZ2
6d+r3RswimkXivbIWmadsY8Ev1M/NSc2uC9t4NuBCvWHM0CcFb62chlmb062XQxz
mkH0WmYmxlIRvgmvHlGp78FLCkCosXGXSZQ7SO6mn76+XhvySP1sYD4xD3GhccIv
DU/kDDaeypfNUfHpjqnwgii1EqEe/TYS6Of3NRy5bCXpcRnS3I6sgdBSSEM86cNN
o1N5FH2b87/dX/A46VDio93+DYFyupBluXk2BLcp9PsKcWSSmu7uO4Boo4XXwMI4
IdvUUNe+ccd9nCi0J3nqYBN4zIa0LDVVw2XQZzyXqJs574oIFkmSUbum45AhXPIA
ShXhyPzmezwr0zIBQ+dDT73J591ConWE/v7ErFI+J6sk/oIQ8C4g1d6VvryPI5nT
IIv0De1Y4tR8bOSjcuWQoDxwcbgdKp6OMu1X/GLpTcq0p6Wt50WHG+dZyRDHQ/8G
YjDPAtx6Q39FZlqX0Tt6FzMidgL+266iFzVFBdiEGlJDWRaO7foqHlrswPu4mYIk
+Kq2mix1ScBOwEOn3bXy1DiIXms9jQi7FUNu5FE/1FjrQCmnKAuIkoM6Pn7r/kfC
MpxlN0AxC97lb6f6HOqJMdZ9ngCzQzKM4/nu9rTH2bmjsLfAXJOWX3WDLzbAon3X
20d+YxfLsssFISx3Sb1wFEHSqT7NmkqODqRsBmb2jF8drqCC0DyyIbYgrBKvR0FT
Moc9S2HrbWG71wdv8Qjd28VRIdLMIzU/wOYuZWhTORnHUZ76njBFGNLaDCx9EbB2
Z2lKiXwv1/xZ5U3EGiUiaItR8yOa4+7RgiphJDNHu0lOlNS/MMZmXrVT1a+BGn0D
mxTG9COqQ7wHGCZH/Oap16MoNj69UxTukBEO0gYHo2+mWmupw6XTPMUIT/SymxVY
jGN1ZApbBt7IHYdYzcYa3+C6vjLmqeJ9S33O4pgGgUfPdUZdytV+Gs175yea+MhR
nADKxcChvTsGu/LqY6gRu3hS3tELHGBQ1KEHczgAI0vPfddtAohff+zIYK60oX80
+g01o7xCQdDbQAsxccURcEhfvE4Yq5RKNJnI3V3oRtdVEPqeXnQa8U8Ek5vnzhyW
wTsU7Hmr3M60MsfkfjuUjJLUzFNv1fOzzXHnpv3IfmajSLoxfGWTGfaSJ9n/OepC
lCJfai06wIdcaO+7lIqGbtC2EzJ5NndR4dTSmm8klqc387aK5t5HmS0tmMDvQrgb
hG7RJBpi+r4b+kzlOBB8McCmbXVtQUXZiThDiHMkoIvHE3JGZJDbHCN/FUyXXJt2
N8FlLxlObhHS+VF+P0G17Rjra/Yu5zev3ftHsvNRl3Uu5wId/I/RlkgAX/PzKHN3
AoRDSqjspkv6uTymnux0/sx64cnss/hJQiAyedVSVm/WpPy2E9L3U9CVaPz1PMxh
hnDhb5oBnAmXA76+groACyuoLC57aRk2PPzcTl+9wlTT67LKyNz4iBNCV1BTfsjD
jgmPkZKhC6mPPJYT3Ww7AkqYu90Sob5sG0HNX1HT+l7HYJs29ye+fgEWGc7d1rp6
btbCf/LCuOG1aUuOO957JIPa3LNGqNyAEIAD/EAtY/N36SEI7apqX3BPgWwwPtRa
bdTlDO3fEH9gf+WBVsyUd848JgSfBDdml23IQfH02cQ8L7HgUqKf5WOIpZO1ePJh
qTc2hfPW/4yT4NNCRP5bgZ6eCHClXv8ntPxZsawkwHrufkUgrumyAJYmsIx19dWN
jOrnDk7TChRJKKP2VwNr5OoCmJNiJyfpQFSaWmDRP0Bd5rAO7XwKl7ccQpk2iSVY
+PtqsbCIWBr+6JuEZb21ebUb/03bZ4g2IL64TtjeUG5ZBYEzCDhkMOCoAABBS7C2
0m3tj4wwCd+oCeVWE01HiqSJ+AnvRxt2Wfl4XXHW5OY0V8iWRtTuAy7BvJFBCchc
R7/jG/UMmrlnJnb0vK085GWUjp7AaDKxwLbdUjtKaGq8nCJ2jFZgJE0r/yPwdoAs
WGkeC5XYjnTNfFBKlsuy908MLkr7T8xPJLPH8+f3yxw9MRiq+QDXHyfGCoi6UoAT
FnBpZ32Nq4fO4ZA1mXPg9D+QROSQNfOl40FL0cfDX0qsq/B6wHMjmmzhhJ7EPqgs
aCS3AiBwpM5i6XR4IFBdS4tjYOX9QSZig23eQ42wGFEmjl/RxCH1o+CqGICwSYhN
f1/AdxEW1JwZgsz2pN6cAZaVP9JAm6HbCUOra5xpDFX+YxIlIMCiVwmG0q4eZhzh
rU/9QWgGsS0hp2kRsDvdfDk1o1mMyetfbLW3fkQ5ObUD3B4RnsJvi3QuuNhKgdYN
c8l3018GlZNWK58okTF8nsTYHPfXhZVzPtjXP3edezt9HdqEwmosGtUfLtnvhotG
gzKwpqYlJftqrGG9nyc9DzxpxFcOTo4SWvbS8TBffbvB2qIZodnZAguq6+xrukcq
L9omQ1BuW3LgU56tws9y16llK+VO0wKTjz3H6TsFjUnhey5YoGTEVAhwe88HKVBA
85JUdKk6N5D5volCzsVyg6s/GMdDSVEi1OlptpBb76+3tQiYrX5hZaFH8qv8MQBC
0Q6GpiIxuslGQ+CeTB9KJ9bbLKTTrehNjl3v5UPJXxfojH8xFPkJB5PztufB1Zxu
jHovf8GLsFjVI7E1oWnChzrZyzZgcHd1HwWxc5YB/91C5yFSuLOVL9jqa/4WWvFY
lOJ1ZMKy/KSMM4l7oqKugIiUWcwpNnJjtWhmU00c9ENm7n1Ume2jpfXjEE07YD8e
fub2oyq9tqko2yV0OFIeodOU59P7ltrLR885Ctw0Xi4SvbYdzvCImbArnXle+kdS
IUa7+0y/OzNlnzJVhOIw/kVEyso46rCoTR6FXzVcpm2HQE0amxI2BcleSQUQdTBm
n5kMi2vidWtvoa3gbTRc5Wi/9UvVODUwRVYTkw1e+V9ZEpeONtb/ejTJkXUH3ZpG
MNKBGmLe49+YG0yHdrCjtX1VunKqt+treJt9R8TPFY41dlHgi/2YVtJv9DjKf1jM
Gos1p8aOACfSSJpOsEqEPkjDWFgNiTreHTJE39BFQeEE6MnLMMDs5oDGhiqYAnRM
tHX77Qj7MGsYpE47wA60pRi9fdQ2qeue0v/+HJtd2FVl3sZPRJk8c5fiFsI3C95x
mPJQ7XFjJh5bg9YKYr7KmDE0nAl+4lP2eXIUP5N8cfhbMeKuMGTmBgVph0uBgrGg
g+AwF4vSLriiDzcbORF3I5aC2RC2ALZuMRaGDmIJNuYo9ti+lcFP+ueUjctPj+Ck
GkCgYqsM36IFfQjiRb+tvDMQXY4L1O1svy8nAvAPWtng5OVD9SQiRcGFkhgDKMl2
adNIgjeppDcddKq7ZFQjdtmQrHtxAyl+7Z/lezwfKWEa6GB6CZjSDCHn2LM8ncSC
AvJN70v2MsRO/uldkSiAfGplHdppuaU/VSA2X49KYsv6p8AMFlPdJRVFxvGSFCt5
Zs4mSZS4Mtz4yBpfptG/5H0a8Y4Yr/tYcGTnaTrMD0EMluuj72rsoiVon6kxqOWC
o7jMS2Bfv5SYb0GGJUh1jUvONxlGaadmu19cjN11VC93C7IhHvmykbLHT3wRQvgl
yY1fByux6n0RO3A8BrL7pXH4NeVUkQ89p/FKFxZbzf7aMIsLGAkXv4B/yhdGY7xp
9uVME//xQjePk3AwQm/jwTKYXy+wRoDybjm07NaImZE5LQ5+domJcgOBjD53y1Ye
/YbtzXX/O5SBUwMG9uAW/+bGN+VXaWPPnDegj5NIeX5dyJVPf/fMgr/6M0vzh8o3
xwbYesuJclUAeu6Sm9aFI1vd9ked/j/cHUmgRnqqhPbIFTSxI38HVomlufH4TbSd
Y7O4fMgWgEBXhcoND8ORMe8Vnd5+pCekZrP1JqCuiKFjA6FUKuhiMKuAcXIFbW4p
+L5E95dj2KrMMJ3xicjfdAZ6qVbmCMcQQ64yvZY1ROonnlE4XemrtWDFsDMvOfVC
pi98sGwU14yQ4Hcz9zjWHKoijujavzfgqEvOKrp6KcljcDcbkfN08C1UzM+56rfA
1PY9cC3pBGU8r4J2N/9JJrLmmWpsA+ZizO+dBzNSfeJh7w3wk1i9ypee69dOCda5
XeyxPsFybezfQT4tmcD8CfLY/JnCIMqxMSFuWmFPVZrw6w1bJIVqtRNrBeLoMTeJ
DuJA+ccH4HK+dAZk37956XWvz0agD2pvUze5a7b7HaTrbnoSlYlGi/iDHICytv4J
lOytAvCr+HCX2QKdCl/pJFF+pbTNIantBNngNAaDDZapfYT0P8ypd1HqYSCgEJhA
m+CXCHcMSI1r2sEwJBZ+frCNR9RGSO7wMg/qSOeuzh8WzRxhFHrlgE+Aa6w5UCgq
yqoEac8t8awaX7t9LwHN62dlaqLH9TQEwotOCcHUbkvD1/YqxXT+IRRzNowSTRrE
aRKDiFvu8aaa4eVpYBevnGCUqzFqtAzdif9KIPhMHfR5DUY4U/CCnWJfTsmlnEt4
RHv5TkRDdAyshnvc1DYNkpWsnzQQeVrHUPWtBq+Bn6ZTqxEBqUM6C7iAhbxIuAac
J6HBHXHO9JrrzWcTCZnX6os/Gj8Bd8vL7F49Tz8aPmIQ9Q3WJLNdTIOhXUwDr/Ju
J+WJnqqelLwULRw8ms45VWujNFprmZc6/E/hAFGyrpG13L8i8JiPWirKaFgHj2RS
6oyREV6axOgBU//DCBoyhzFQMGP/ou9p9DKDV3CC+uL5ZMxekiFwqR6JdaIFi3dY
2w5FT11vD4yUEEXDOS8naCqBh76I+MIlVbofHuYjbfkv640gI9f3HWtvFot0uEiG
eTc1V1Zdb5uFr2KeCRtnGfNZ++TNwybMV97L4RfyKOj9bLnhNJFrHfXwghQ4S3c5
rauBJD2V1l7/fk0Zv9YjXF83I+CKHwYPdUtEKZdv2dIHg0I5cRrjPjpFX3M/vprO
WoLQjJLS4ddbG/Tt6yJqcLe530d8FBXoDakcZ5X/G+bgXUf4cpsVYgCHBOFVX4vE
bJ95QBAKB9mN9VIV9Pl7k23IRKyLVSb3yGT8sYYaRCnptq6ZtO7OWOFAyqE+nEN7
uTsKO/XqtkyRV8DjzR6lOywalfn1CeuMKn40Kp7DPgfgNa8DcmNZWqnjq/rUNWEJ
yfxOivTD6hv4V/6AO0apnhsFhUeDbBulTyJqaEjxfZMsr406d+SOt0fZRBIVrIK5
0LJ4YBf9CdUixbdY233d4w98krQqtpcqnSXCX27DRFSvq2cEUIrB9JE9iU+cVpOC
aECX0Thn1DjFtSqC9QCjM8pzbX1GWR4wYTeeHneod4LPGLdF8AgkG2Vw3zDo4BF3
YpS7FFJN2pFw31GOdgt8WEYhlxWN32LPkX2VO3WZ46dOW+LKn/dE81hjhnqjf62G
jBfMn3BoleMZDTeV9O5YVzFN6Gi9WKdunlVUF1bLulcG12ZWQ65uY8yqCe3EYssW
XeC+1moMDjx9TIVD9AnThdsH3aWUti4mail3LhC+2zSLiplNT5hPSNMq96iQINbo
APmtbLBu7BMAzagM+Tgqnq1Ja6exOqKg/LfzF2XDoX4lMrv01yNpZNK5x/DHuHZU
cMEx2iYx1MVWFMbD8unF8wrsT3BJZ8wtXw6nJBxOi2UGYtO/dkapjBAuW8GN0Z+e
ARudna8H7VZPS5cUyU/gs3TIxKnfUu73rt5DOIW9R1UzHC/VUdbx+8a9SQ48VUvz
2zIuYNR+slk9ZZwitBkqQuJnEUwoV/FHGkLFlWTObAHZ2EHsru2sy093hcpZToj9
fbq9XWVE/SG6KCA2w/Hs/J/ym5tkGFc1hRRruTGwZ+p4Y4ab7Nb3LGy1aY5wNTyJ
kMD3jprbJwp3x0V94QQaFJu0Mf/S5HGx5LaonSr4FGertDrbJHPRLrvI4J7GErNZ
2xWa4X1SkBMGlSeqHousDzmteSI0onl5RffEkZwxmgUKQH9DLs5QKv3T3Rr+RZIb
Ld9VfnfbCzJEi9PiTMKnOuUgDIzqm+WT7kj+AFEhvzh7N3CiOPoQ+mB1osRJENJe
hKYLyK+frW+nmG5EYU3rDx3nxu6sl6g9GFme5COP11lqOeY8O8VpmnszOJhc5LeX
fHlhUrI0UIa2tBHHh6FAItJRd7MrPbDV0EKUxxWouD+ICjWHDDhrWPz/fDcC0Jje
ntDdFxHyl3lHaqKbJmmDQKV2uoRlLhchNKYvmkpvfpRc7xsxQn9STSE4ot9V0ZcY
My+IbfQY/ZA37JZMzw4MAFyBj7pa5Bw1gFxAAXvYQjNGlDooUKnKIFKXCx7A+RGV
6ss6JpP/MBcleQYG7Lln27k20Y7E+BDZy07eR01Ss+qOppVHAxfYxT1Z+ntswtjy
qEHldYdXFc4cziHgMe9ilvbhrG6w3ECsKiz6leAY5awfhvtjwMq5A3iNZFaUJA6A
h0u0UzDaa8bgHoojm+kBIoASR/Uuhq0NvhXlm8gvofLMKLg09A3Ir9iy1Rar6Fmw
AZfSQzNmLwalv1QPh/3O0Upj55yRNaIG/YxieYmAWXiECmjhncepbnYKxVUqmZqw
OaU3rvAuXsTeZoTaH+LOkZ2WykVruPobQK0dIPHpqNFZGYacuujfuzMoGx1fKD4h
F3obqMEf4RBzGklwReCBwLLsNCpX4Mkv295ryBKmsBDxYXrmlUANNBC0yZ1lUOuQ
kLFHXTCJmYh2YN5ANN5FgWY5pAqW1QtyxpM55bEQms82mj/2W15+EJbCR75OkGjD
KvKLl1s7dMpZQxYuwy5QVkfTJvgOIvzM45tFW2SZRGD0MN4WyVcoA1rn3AkcbLsq
eQdqIw3unIzFni/hQwCmRsxQ3Gnqz98NNY4qwVBeM/hbQjktEf8162QXKRubUqsh
s/p9HbOnfRhnBC4f1Pr/4D3tQTahuJzbYJ4Wqa1/Kdb+5IYSsCfQsQnQetsIQm2i
U03We8t3oavREEVevUvdzqr/cT3dt54W0I0JIMV3HHfreKEcAnwBvnGMhKRNUrZd
bwyDR/rFCVP97rrNm/S8VXkY9kYDtGQQGyAnUtHN5HkZemX0gaAzmZJS+mkI688v
4hNnElszadMZTlm2yc+NA5BOLHRXG0f0vgfdQmdT1VumNjYlBgmrrU9FNE+YHzvA
5KwOURBAAyr335T+HR+ZruajNsFVNQFNWgV5pfeP6KqYqYHYg84Ozz3jy439ddES
0fzNzxoAjNwZipKADwBD3NdkwQzTfXPXQ46YSHMfn2yhpaOIK3HKLbcwgaE3+Xki
F+UwHV5Ehk6WeNiJ5SGSdLeNI70YjIHYyB9ABl6aW7WjaeB5JZgSyIcpnwqlwoci
QiGJTIh0Ez++XKFSO8xj8m0LCLzly0Nq21Gianqmr+epfxWOSaD+Tx4OxgijUJ8y
MVf6Pbd0ehw7O6YcQilge8sHox32eW9VY9gT/0lxBJiAyi/HF9FXEGYladayHCxy
NLkWETIbYIZEwVv88jJbITvEmR4imXnXs0+xDDaNkqMoTSYziofTxNiCg2IdvxPT
8HYBKbzUbZed2G2nXjwixOe4LEAprpyWdx5bHSz/YPGWLxX41ZflyMnwdZZsrldz
LGrygtziEDqlagf7DGC07+wlthmjuUI4jwmpfz55avL8YZH0gBS+2/CRI27PMrQ/
rnV3o9ATIhDp8mItat6tsrdOS/SW4B5VQX6H9rMdE4L0NQzMeWjc/RmlMl4w6eLu
ASHv/RLawBxOPgOxAhK2YjYn65daTFTkXVjIuKXwzpZYsEP7GOvzCedn2eVl3U6m
ztv1J9KOJAeJot50PUxkJgfuJfOlDwPCqzZ4Wnh1gNqBq+We5NvqpRLFU5x2obx6
/MZOkfw/aOVOsKafX0sFRvcBWScCYv8KPcrf67LYLIR3XsPXgEZRSJ+aBlSL7VAy
Ae6jdgNBh0KZrpP6JcJw9CKx9Dj0UGRJwDratLAC0Zx+v0PWVuKDmGuCMl8xZPLg
i2GN7Kclgqb9j8Ljxpo5YubuYfI+IA+2Jg3m+0vHsKjixz51ITx61pVPr8W/yQF6
LZyVDbYybztL3o6yrpR5yWYbKQRHBG+em/SsIe4N0GwVHcA2AtA8fiiFX7dvDAZJ
kHjCP73cqFqv0eFAPurfH/dD4ExFSQcGu/YOWONcNqcMW8wDgXO4as2gRz6SQq1j
75rQhYzjMraTWK8zvbRSnykAWe4nfol3QxKmWFY3ey0sQjxG7WenSiDObhtIm1zd
CKcka/nPvAAIwW5qFuH6dRnr/TxGKgcgAvnyRRacn0B1eAvus6tzhBaeggHxMvyP
Rpsb1JoYwnjwkcTuMBliYxaY4bh+qux8NQcS4vbumwSO8f+WbDegjiH8wBRUpu9o
IJv7oJY2lfCzTTQAG2SumQbmo2tO187TyaxEIBckRgY07wmtnBf01wuucmvEkON1
UotZM7tVvH/Ofe/IfqDW1ArC0pL8DjArUHKMUW/iSpLRr8OzYh0qDUJE46lORPUM
FpD3CX49rnEMn+um7qtCblMTCrMy1kZR7zcBsgQTPA2aj0KDqisM8R3GDbYSHWxX
BhR3iribapBfg1TV43IH5H8lFffPNfmjYJpbxRO4lPnuIQILQgFyfjyUvGr1H9nC
YoFtF4PVPb4W9+UncJke3fL0EM32/X6T1gL7/l0pZ0GlOB7EK/pOJ4O/cAYm9Iq6
C5ObnuMu1KMiIVIw0QFIZfNT12AkWjVT8KQhLP9kS9ZhK74qFIKCJxTsEfq4iYCg
Pktx18EIWwXGSHdCF6Ja9O2G7LEbAPmrnFAZgN7cfFU9lANi0RYRVm5tHRaMsKBf
Bkx58j2j5IPjWOAe4ml3ZpG8PExkmFfocV+zwe28AZ/kpjrtm0tVLxc/JjWLgExp
6aggXOc32W2xKjNFiUe4SN/i1Aoz9WSZNcy6ilMCrOta8WBOLzuJ16Dx57WGDdbk
b0PLfNucqTLggBtNK6htO9LnKlsAus6giW1HpnnXme+VS6YG6r+nBfeT3MyOWwOr
48R0IfU5RA/tOCQjriELfV9N12XnN7gSyn9c9bHYgaoPJMeLlu2XxraF6Nn8D27I
faCdc3vs8GVzekyW3NuI2FsotC+WiWIrK8JvOwT98Zx/uG4/Ff0HZSnsi6tSmzUH
EpR0M6bnEdzRjC3JMqNqEggVZKk4xtjhLu044EaED1mPz/DG+EiE0DWE/c1HaC1m
jTlgbW9H69IjF7brfSnqFb0FQzkAhVU4QnqlT5sJ4na4MN8QiXYpaajnRuyE7Dg3
E02FGsSuRpC7x5aQfVcv0BX6KtU30bU7cCJIVT3NLOq1Nzzkn6l2rQXH6m+2Kjlu
seMKvGmxiKeqh07LmWtfjPqJJ6QDmc6afjPstmYK1Bcb9bamVH57eQpJJy53pmBI
wgngzJoHN7sWDtRG3+xlgFfRNSb1fqg8qcFvtA1BWZr4Q8UQPTJshoJjj9lDeX98
JUOFfsn5yKSzixO09+rw0Eu2l0cVidCdUG1gU+ag9iXPEplWd/4l1Mdr+TqTjd1l
pUhhiWZFpdDtSNJ/bwilggMcKmXQ3tY5xUqDnZRa8jhO7xozs8SRpjgthKNvlZfA
LmW38k3M4TjqICeAAmdE5ZaUUf8tNTSrdwS32padxzWSc4PaBIcssecuZQG1/1uV
SgXljR567ANg6/O4e/tLrxvr+yhi6F0OaSjUXHbSw40Uxp5upXzFj9SM3ThNtxUz
i8qPIzSoL0l+UKts1et+EUPyuYApW7Rbox8v8RFHGzWhjvtYxXLWdhKF1VzIA6+2
Cff5NPtk2uxLUSUwofLzmjM4Y12XzXsQxbbEsFpeFlLP75Mqy9XeBbW6BnBwtPrK
n9f4rzfcTt6rlFGytpl0dLlhjFb7ZdxanMeK9cxkhXD/mx8ZrZZT/MvVkVPBH350
Z8ejA1RhK6lnQLt6NHtNDXtpG34tzjdXL94rJM+fdrConNs9LQ1WlL0J6jq1zbSe
VC5pC72HHoiOvHWo4XUI7xteAnPctl34kgank5+TpUMhM9WIDOshigd5yJcKw6d2
TTvXBglnkCKJML0phulLVQcBXOo+qU7vM8fBj5R/4Zm4OR0JyIVo6+1gcgIhtWH8
fe14Ob6VYzj+ov7+uRNXsrSnlW4gq0C7upbG4oeRys97b9A5BcfmuplpmawQLg7e
wrcJ1FaFiumOsKbxDsu08jALl+8EozT4z3Cnf1QcBm+x+rihf70HdhzX/dDvM4ne
3vAh2INg8pHXQaTZsCXqrtcPt68B1KZtdl7HWR5xUnCBIUJ9Zvz5xHMUHmsDwI+E
amh+8znJsBEsBxljHcxjPm6fVRjE7YpXR7F09xfPGqmF+mSKh4Ae9/b3rwFzYEzL
+n2fViRb0evKOW/BRQOepPuibWSFWDbcs17Xh1K09Ud1Pm/JMJlOk1EtHt9zbxdh
pGygSU0uP7915Z4up4bYJBBErDL9yijBWPS5+Y657Et+iq0ZWKuVoBlrQ8/0UIJC
cl99ZPG2piaGGzzBMztjm47AXr6JpQug+tovk5+PDPA2YuKZEn687M3oAyfikRSv
AslodF3WAZEJj99RategdmjOZhGbVTAQYls+I/tezCPyvldG0OUCrQ4IIVCPCIt1
FTZV6zdeDeWFw8r/Y9+sjps8EvdSW/2Co8vDnqwIlVFipqFYcLLsuRal+XDiTxJN
ggqs/aUBNFmOYO4xHT+otahRW9EModgh+uCASvMoQpDxkkeSwfDvF9D6YyMWDaE1
7+CJKsa0q7zhQci510SOiYPvcIMXM36EsYco95QGW0oRmwB8FdSOc/uL1N9QIt7i
uTsKw2Upu/s1FyFgz2S5x9XEF6KcBOjLcjITYGuEOLnl75bP82lANfora4fhgTfK
ry+CmuFtpVlrSD6r3ISzcyqMVLqcxw/CEPMZOskgtN+tOcw85aLZN7TwbhgL8eHT
Fyr/M4LwvoOuPRM4OssbP6ST+Y34z4n1S9QDMUef9P3V31OaxlLmkJmkebtzx8qx
dSNlatG12csL0U7+Z2MRz6rwElQ6MOn4EsusaMQ6AwnIq3HeNFdvD/T+Bov8KuAD
JDsZ6heCUe0rTn2rs5imdomHidKJ1LX0ihOpRCd03p4cmL8GlzBPyz1S8CPz/JX9
QqsyD8ExlBZgbAqP9NMcoYVaNZ1IfnIjiv1W02u9yCIACT+VhP8tX302Qqxr8x9v
AWW2Fmg0YPZhu/gyPnFcpdfT5QKZPvQiS4rPjdEMHamotbeERimnjsdK0TNRYeTp
r80fXqSSIM5AgMF3TzlgYLEMvB2meDC1gfhXG55lkyciD9uZAyPjYBpjPYcHg1nT
uEJg4vAdGv0BNznKnSK4axwVodBu2C41kFCd+6ylFcQLDs6tzGPZKFg/SK38cp05
JggrxzacNhEqp8642spj0C+rZ94QAZY146ntBhLSWZPaxiGsraUvwUJt41W+kv9S
1IwK8Oevpzv4zNHoNGwEPc2dOLU2hbUY15r98rH00I74topCmemOGtXEXPhOr1sG
pcIe2mbpTTD6ny7gPRvWGxNIjaC6PDzkyEMZGkCNtBBfGympUxioBXamaPY95ekK
nwpeuOkukfAVdw+/2zBPkRPU4aOUNejNC142Ms/D+IC+LQ14I5KD59Fb8P/Ygda+
Ff20kWjxeeKdz+kbiz4tTX8maAL3NypYc7FR34cxD9o95B7GVvmnFN17jUJgDqVn
OvgZw9AAzMw1U1R0cCIVYZcUlRf09mUjy8Bw3JyzQY+gAgZ93IIvpJ2ykEq8isrF
a6F7QfgY6WT5xv5Lh3soYIRZe4ZWQAu8sflRwzmPMgjit7OmtduYBDCNkH6h2y5H
q6A29mwcmfmoP9GT3OJmxmE4RI0Dc1sUBmYtj2yF3nTFA5LkmPmaY2PC8coF6Phh
QoEUJMCn1KjrzSptKPAc8yUalgKfsT9E8fw0jYMh+2n5o2I360nE4K+k8IDyObrb
xEILnSp4IP4lghAufdaTSI16tAIvxPS8K4oYY9OhFTpB3xnGI9wETFw7fXSJTPFt
dqDSA6/G+W0/dESMwgeVFaCDF9g9Qi0r4JAvdBFdROm/8Uv/nMh8fMWvIV3PSl3P
qADzMqmDnYCuQjHDHGnpfGRsO3Km+cnigb819jkKS3j76cTbG7yXL6sGgQazIeIw
PuJxoI7000MW2BQTA+AW3WJPb/p2utY4gx4qSVl4v3K6xb+3aPaphZovsUL/YwBE
JC38PrQbe/5Oqqfm2n/JYBKQ7hOfCRj/ZnakgjHe04nraNOE643SEJHwW1oY3QSk
Afh+vAX8spgfEYYMBxEjzTSwD3T7nho8iDrGdIGD58q+bdC1QfOhYzuQ5qqBTnGA
WW2oStCXe3letmVj3IUtCEcOBqOs8VL0YbjeRoCPOFouBdic+WVfWW6asIO50bLe
DsqJE4E4wk6308ajFgUC/QjPjS1aVokqo89U+nfEc4jrPxpfjCcfZsdPMkA06Ejm
xwAhc+xbXgrUFKVidhZ5Yv5lyMo3KaN6zhSxsXkZI10bWEfrpY05vLuMZn/K/se4
iGZgp4AcIlcVb4uqPTL2Cnr+MU9yemux4KGL4X8KpfDyQ3y6+QmKmpBUG6+v9kmp
9RIDaONZHnmsIsS9DysC1khiDxPoglqvSJOcEkWZj8u6x8SJ4mqhynUFIq/qzLhf
5vGBl+k8Ku7Fzh1DomzlkD35/d6VWMbBasYaGjRbns528yBdOoKQ4bgM0fFbM8DI
PDcPSovlci7vrGZ8rj+y9cbE4x/5AxX+R7DIuFTFwpjUsXnf0SSex6rZiDlN2CTn
wfRGiQL6DA+7a4Qaj4EtFLeqeTbLqNYHkogzb1hBfCDMaC8qD+PuOO44T14tQ8oZ
PPMwBMb+sTuYshi9PmRxuHoOMyxq3d5un23InqpBTpRHFVD9fb5xixsLIhmJstUK
byROIG6AHW0ct5toFoPQxEER+ITxx9hcNWhsnsA+091tJBMA4k8XZQ0EvGfAPa4z
w7TBhsgKaes3UiYVi8Gu6Gi0+L/dTJXXjHa8l3ncRxciRNzYwXzzAxJqVAqwzb5w
LcGRYmvF0zixXj2X4zmColVkbLZWBhzCraug+8gHqK+S78lXN198KrJxKx96iu03
U3/6TC59x3G7gY+xNC2Qa8DldQankXvOGEvGPItthEivQnQ/cVKcnzMCzB3Fn7l/
qv56PFzKELovXpFicJnkuN61ZhG84GL+1BpUP24tdXShX58w838bhZyl94x+OqBf
phSnuimKV/VHBN3bd3734jyT2LV1nEXhYb9yXzjIAAVSwLz2sxSMvnRd4mPdjIKV
lKDV7og+8Tqqm2eQjDrzQN9TYRhjBZChsmoy/AzOkqfjojB42JhUtJRZAfxPcGiq
Wllb6jlbmay3+ydF+dC/4F+USq0etFvxjW9pr1CrYOn0/pfs19VCuW2UbQjlDmVP
CiJtUMd/fGmIb9qyy5MWH56joez+hC0geyviNqXl6WiiB2OOG9kTtDX0E1864epG
eH8fQLgqXjYCHn8W4nzIYgJXm3Iz+WqSEP/w2I5wjLqQm3WZzpYxR9aj2/CfbLDq
BUJVF1mysqsIpkqwXMkoWcl3FeS+yZN3huIucIGxJGmuEkt1OXt2+S+by4Lz6AlG
kabRQEuTTfQOf/+YMiHEzrTSHawaTiYGtcOhlTPVASKriM6swc8j1mH+M0h2Rn1d
vwfGRj+3KU8x4oBLciXurbqwWgUXB2BcTbD3gKfXog3GeMYd37gFdAqPbItuLc+x
r6dbCjeO8hRcK1gyqquhCcWXkSHhJsRc+FeOtBaHDpDrfGXPCoBIKWvcdClHMjOq
hAr3GJwlToYSwzY2wmZdFoKveKErWZf5IvTd/su4XEsDaEpfGVROTVYSWGuTtyuF
4TDowcepgl5OFGln1dBYWuigdx5n9O8U5zcMJT0jntrMmcZnQkEj05O6Sn203Iqe
ji8f96txKdnrzhFbtogN+gOzmGm0e7pkSPShtJD8KS7Ck0IzAq8STs3ZO7mZzOti
SF0t92TB5J90loUgFcCR5/aCyJVIskB5p6rgxCiOgCmTui1DQyySpLaWtGJ1OWSO
9mG0YnVrTR6Xjh1S+KEsKY7k50rOP42iEpbiV8F52+SFh7D5yJcTXyCTWrKlC3DH
Q6Vl+1/yQFCblS2N0n7lECjYfsu15GymEwDBhntcQ9tQ1E2M4aMhBYGR05603vTp
bm51lFkolxCj5Xk3r794tbsYT0uFz+qCCx+14aBnKC07b5dwVG09gcmaq0ct8QW9
PiZQQ4B3k41uI/UJYb4oZhcG2nCnwHU8Hq/kr3v+26xWkZ04B9t3GrZOek0785q8
/FSwaxl+vgQ+/YgkicwovQ2FMHLROxYujKupjr1LUXndIRHhSsCuiL5dcUhljSR4
lECwiVnYrRTFIU8xLhxEC1iEk4M9Vmv7FrrFKLeSP0hdkVz7LrXJgCK9Gv0ZB2a7
kEQ0b1dB5ON9u/eSBXNQXzuBUSrkrThv9C/soxln9G7dwtGu4RE/TjCOqPWEpAYU
4yrifHlzBB9xCLAWPpK1TNJG5wncamZ1z7x70PEzEVHWxESx+p1jGqh3+LV+nn44
3i4QrwXxbrqsQ1X2NGKQ5JO55HSoJn3DkzOtjTrA+K7J/HbE5rNabctcgz2pCDlS
h0BVW0xGZzz2IqkBDVVt2eMwMDzgCCjOi4GlXqC7UjMY/psN9WK3EeKQR9VjCUI9
2pdG4E7Dsl/MOWuLKrUpfOD6hVCDYapuItb7H/r0lblxRqiYMnHqumUsyAb0clDS
acAXbrX29c1hpcNAmDUNC7vAHjX96YVXQDIiLkXCglUr6dmqjsiovE3V1PM0NeEt
y+Nf8kAv3JR/TqxfAKLlJq1rs+KgQgKLEFaEdLFfgGDjZqWOcKsG515TSSz3eU/g
mfunBD5NKETURicmOrhKJVmmtrHKMiM7MMnD64hvDgJGROWBtOpdS6fN6kg6/5P7
l+mx+f4X5uhWuffamkOagfARabUGFDJQEkKUPPrPSmJklAoUuK0aFRCgFbcp6HKn
YwZ3msoJ9TqmqtXQcQ5ALTE6yCmIfLu5O55McS85N/zTQpIAuxjFd2ZVKjb75daO
Uq/fedtWIiK53YhRWMNtz+ZFH5iNZZ17mugntsvu3FNyNWgT+TMTnhIOdyBLLoq9
2iIw0vsNP3CVLR9OhR2FldcOms3hFukCSbbwdIGKbu9dLx6GbqYPl64JmaBESeQ9
ae0JAGOgyJhDX3Fl6rymvfUAw0szmUzPDmCh5g5TlPWh3wYqjP2bzj66X3qJ5FQU
/jYt5Wsao6yOpnRAj5exL/6Of89ywc+LMVAb04trECakyFMPlJSNic5RIY8e/IaH
sfbDDElgatiQOEJzYMkL8gw8bszrizdmlK8+LD3QuCzrF50EnIeLDSrp1bduwb3T
/NkoZbkYpSy5MJn9KYRHjIOF8RRMqUiJUc96tLpqsD2QwepUggcyxdY52JIwudB4
ExT94oP10c8MhH8eXgEbQeMA/ilitNdXMrm0xCPQE6Cd/Xh9kfvi56rO61hGp6tZ
VkFRPB/MTBlhsMVAVWZSELzAZe0ZcjzXxibmzf3dsqqO9OATC6Mn2uwBB97d5Vj3
RZMr99xPWgb99qDm/M75QAFBPC37fimpqy/rdyzY/oZFTzRp0H3UXExfnDTPu4De
8hOC4YrbsFO/auzAHpihAgRCOdq06ffRYPT2/Fu86QyUI4voF43MkxXgnHyjhasq
owk7xdLQcZYBaQOdXm7zwGIZ9r7LRx1s5SSrs4UgQVbUeMgZGvz+tFlhmr+Uh/AB
olhaml2JkLzECJhM6zIqlyYPGAIl2zL7bw+9/eJJnSOIJel2QT8rRfs5aAOfD67x
z2F6Sm7lo50WgCNZu9ymUG2Pzskgq9ovY5sL8GsBwK+0p+XaSxuVkU0d0xMWuaxb
iYMzRP2hELqThGHZW2xKENhTVPTfh0I5ZymmnAFniNacftWSOVYsztlmMJEmhAzB
HI+VfagArDNk2jS03S3zp6MVfwX4cGj4dWEJFBl4oRSRHZV62yds8GvYLpSTBiFL
hFdgVyAJRXdrWVrt4iYGz7QU8XazuX1Zm4QbttD5kA5NopCzQSSVQfnD46B3BD7Y
gzQqQOp1jLa/8y/gdLT1go7dxm604dxvJqX2V8b9gRf00b1juHbvmcuLfkk9QeHy
1HPEBubsRct2ixA4Ec+qIDwTYva9+Todo2w7+IbVk37w1mIJ045e1BWn5ck/tFgl
gbjimKjpwRg+0Eb4QRD1Hi0ypdtP5je/bugSY6maB1L2IFTwT+HV92mpayRixvWk
EE91GWtHhfbGCafRr2zttjQ42slwrfvYxFN2svt1F8/4UbHUQZf41x1g85l6Eemm
BuUDA4EBbsD7kfA88gNiPO99ozfy+XosWl5ROXxG2CFj/ESWUtEBJydSG0X363bF
9ZqzIQzEQ1V0JB9FgpXpL4mXMSpDAlhlG6f/UlSNKWZFuvUUAxK6gGmyVMAQoO5p
awRYLPA5E/VKU70AVOXuK1IJYYHQog6uuqzvaudnoe48iAS5gWW9Da3tFdqy8jba
qagnk/YLVJF4mj+86Z0jrtdTIAGRgiq7fsptdfE65J6Qzab52I7t7erurMxYI0f9
1kg8ij//3rYisgDR/gM1CC46aJPoGG6v8hbgpPFyhygTDwfCNeIw6cEsKLCI9TFM
koyHVe0nJ+yhvr2451e/MgvX8DIRpYCrU4VIKE3O1pOytabqRZpYZTgBDmxnkRU+
NhuEpnGVFQIYjN8yz5wS+vkCmp9wJVlNQ2vk8rCh8yUsuiiLHeGXjkfMDbUBSZzp
G4Hwc1Ce3kb4vwI03P1expX9uunMdxtQ6A6PlvDT2+5xdNm1ufKyZbU+CqZTcNpf
+a3BnORjkeaGrRpvGKYIsprnaFq/R6t2DlAIyvYmvv4lK6iXAZPWu1WEcIVzhJUM
tGGi9kCC6/SQI2xZc1mCKn8E+eCQd7KD3PRdw7LLsFFrXtfVoGk8wRvAgAI2VDLI
Tui8P/ibEKMdS4q/R5BM9UspMQTr/lzC9SmuMJxOpm+5XC/tFXHoSxXFyEs6YJIJ
/rFwF4zKm1oFABV6e5gETD4VtrM/sH5YCFhqAQXje7Fv0GUicGGazwH0Iwwg/S31
aP9iUgtzKaUt9M3o1cmMEB4Dl3ZR6QAAB6ql9xG8UkQ4d23+omsIMYG2nznUuXFN
19LFAeFjFYCK2Mvsm/op928QBVvsMp19utYXJjaUBbF9qWjFEIOc64wF2HHFEOdQ
Yiu5Qsf3EtvjF0jp5jTrwpQkquMvumDTiV4rtv95DQo6chV6PQKy3n2cC3W9hVg3
/fF7B3RBKrhdMAnlZ5Qpf/6JZPyZq2USMiF8YxD5EVBEGOxdKG0pHn2kHWNKWb3q
3UtJliFk6vzFm0htvOydHEGv8bQYb8D/GHPrJs9RgpbvDWiGwO37Lbw5RFwbryPG
6Nr2UGJ2f5SYuIz1QGBHiPVvGGDqBM7LubmPGGtHorT1+7bAwpl75F3TsMwAO50v
VtYiUh4UVIGmL70tVDmQ8HCa5vGXvDB+XqX662AabTydgSNaUPcX+sQvo+KpPwdf
Zrc2saSWke49tsoxY3XLjdVkLM9ovkwlVeYJVOb49rVJH6KOmgyApnzpIrTzj7r4
QZnYm95SJWZRBQhrsqBS22FL/y5iJ2toXjnQ3mLk1iL+CcGy88NnpGj+Hv6IyZu3
3u6cu5ptVIe5cUAZ890WwFOB6G347vIasYL/EtB5GSPzr0s0uBOhlqqmRj8wT5Bm
ok3NwcvRZRubsRXa3MhT7O2hAAexwJiwqr3Glw7x5zFQly4E6fnHhGDDejPc8qND
n6iKmfh+aG5eUj+cDqlOyukvBuR7cUvPhL+m0naZD8HGV3NpxMndGiO+BJMHjG8E
UaSTzyThCuApyH2+gI+V7cXRElwwynqTm00kknBOHMzdu1RMqCo+mfmcDeX+G61m
Cq44qtYkgPPTl5XrvipI/AKD1uhaNSA2N5NLGwQJho4f1Z522j6YoJ+wjQR0eXZO
FmdXZZRMZ9y110h7JO30xRzQzc/LiUO9WlF3TJbG3MbTIohNmsNxC66aJmqklVdv
sro06FT9kUW/8e/Mb0dt7v2Hbs/+sRaIIGED039k5aTCp3xBp5cJuO5KT8SzKhq6
ok3+9SXpwVNxFi8nYtD/MSA+9/f7yKv4MCHPLcrocVXHHb8WOmw9KuL24ORc6JKW
puPrvXpw3GAujzd4SIwdHbbJeoa/jd1VbpOtLZp34l3ZlMiXKnOs3IVA3Xc73Lsq
Qr2Rd4aUQp5/ptxngBedzZwhMC9Sz+NBAr6JGebP5yHeTWVKAMBRcVPTl7PDHsF5
3jBesXyglEgu5OddJn1AS3v05WB985lavIIJLfPljsFSRWeikNFceGGp4ueN01j1
1R1+AJowXsRMid/+yTorceaofHNNmFaZCoUdxJulGvL8ic2ncYZTBVOYu+JtvyFr
IQWJr8ygwEm55RkpwbW4GQd+U4syLXycfEfsKBGuaiTkpSCw2/Dm+XMOw2BYY2KF
5q6bWvYN/3wwm+gXHfprbO4eM+FpPe3EGYABWm+5N3SnMNgFOZNT8ezq6P3brmv3
GFVR8uTkBwJq7OjsVt/34qs8nxkvnnCvTQekoj0hq3da4BpRxUvQkJQJK2fSM3FB
em4saQbISuACvb1l98xXne4Yaeov6cV2lCQXNcSw0Ak5x22ln8x5Ov3Kk+6HzkiE
lWYoJulTPTc/hprnJtbacBxzpeKoh1U1UMBHIsbePEjT9g4Dp8fC3z8zzBR+Qyzq
MAEM3pBR0bbCCKasEs+YTiZ2Rhi/lvfUJUGIMhSLjP3qRSVyZuXHaYinuxUaiMRo
M3wtMf+OzP0rvoPUuniXmxuOG4BP8OMKyGwTGwum2Z2m984O+IeD9EMvbuYLSCJm
Act0pZ+rkRB1M0rID819mf6S0db558QGO1VJBvS3bNCGnv0eG5vWrPZbXd7f6EkW
ef9/1FFFaeJL/r6Xb/ddIUu2dShk397VrU5v4Z+cCyQzr+xnqh1QuXwpItxcF3wO
iECfo/kB9v49qVXyc8inA+Chy4OScaKcQ89DPQBSS3AB8rl0NnOCJcLkdnkWqVIv
cq9NOWWe3JAG0D85YpZa+r/1ZoW5uzdyc6MDamfzHGBoWrZlP96cn1BN4gJev6Iw
sLlAxvUT+VjaL71NC++kqyiJD0O0TX/1uYhwr8v2P3nJkpxByhDxVXV+gxgHTfxC
bP94fPJVeB8d6dyYHR0nqqkJQYwrdktQwi8e7jqpJfddGgPwbENbj32/EMFKVfPP
4ar2Z9o5NuDowq4nZNWxnpD7GkgqyW51tWM0+IeGGr3mfFZnSTi276S2kVr/CppE
yCLkB2Rjmnt2v5qFYNzje3LvGHQRE2XHWaSIZ9mdy/SE8RjTafl8afsWSZ3RI3Hh
SrTFjS0p64K/SHq/JN06XEdlggWhI0weBt5u1YLFbezAErWAHELaSgC1aUgh5o3m
UhXsdcq3FHMv7SLSgJMONwtulM4VJYakYUV5LvKu7N/AUY9aChBcXNoZGgbshRPp
c34vcniju70KG74V/SL0mrAATP7Q2lFKSNFuUriEz15GES8wJ12uYAFHaQ2Gx2YD
OtIh15UOrStZkPqiih242Bslu5Z61U2YXaHyVJavGcHaTAFl1JymM/h0bkyzlZJw
vo+aIZtsfeqIlBuOX/yhy+LesR4j0wCf21OAUZVdjwSPH0gbO7X9i9ucokgvVIw8
zMSd0iakMVswIanx/48udh+pQwsqsxHgAKhgpe36uNjIDbP1kI0iHLm/zQo9uq6M
I2hj1hNgJCm/4X2z3zykUVH5iMCCgb5dyNa7CZEcz5dVtbbUWHOWS/IBQXcB6fJK
PofE+naAf/69pRrEfuacAYTuQZ5KmZxbvXYamyDnkor1owRCp10mJl8MRajMResa
xrsuyxxPtNu7kgMX42oG/c+1uFYcvEFNIg+zwF3Q0XOyzpg0qEX8z27Fpt4K5yz4
CP0wYU0qJ+i8KNw8gtf0he+gtJvZfm3TF7S8Vrw/xA3ae+EPIECVx1fb8fIkxQxj
CMxUMLei3F/pxfvC3nQ8b6423PQVdBUD6vxnnY3zDJDnc8Zn/4oyNS2JIqYbHVYh
scqYEj6G6BnEGETnfN3+B8fxSHDE/qnINOSy7/5KuRRo5+QIx+eNZp8gNQlUdAps
ArXQZvc9COnWYVp+eud79OqU/gSzkMtXHXzLDSFgbnLy65lVk3l1jgkRqHAszd8a
EDKQiJOZoajWJ0jAXp+g9RbDXd0oBqGRUtHhDHcaY7Q9AWL40T4OR52LrHdThDJb
ZoznN+ZgqPrNCLpsxuDNXKxGY0O7NqntZJGPLQIjd70QwUMpjl7+K8u0GpmPWZi2
76NYi1weNHzAu++MkinlVwLfbs0DD/LigSvZIy127PGPtcXAgK5CdIy/tjBYvbir
d2kO4DRBL3+LBlY33xMszOzSx1VXyc0+HO9C1gTOrk8G+IkcYctdHxuAaTqRZWlk
gQIeoHf5ZRO0za/wGtLypkQP/ZaKI9kxb3MmeOV5XwtJhatU1FiEMtw8BlNqfJOO
rIyxYDoIB5DuUP5hsaZzhRkCk5peNUhPgaKeMCoTns0wsgM81NTrJ+IIhLKe+oJx
p9hz3mzHQmAje1Re6IGCjgkI41a2VL5ccpQn70F30P5kUJOdW74eePYlTVMCWOao
EH93LK0Xb9pcU6F02QfBWtxkRChTCdY+5mTfesDfJOplHdQ39yt32J1WglGbWEXF
5rFqduNa03dKai/VeMsrZticdpjsQHq3fcicF93p1Hmzx3J71kOYXKxEKxuY4rnH
fgTfQtm+sVqufu+rjGx/YYkKUtnwHXY893GsWNHamN/lMO5b02NqzzY1QUXPsOhv
UFzsfNspc6RwVhCStb03GRJ0vcmcYEpe9vhtUPb4k8tibZid1oZP8AG7yw1drxak
D4PaUnF5hKPCnnA/0p/ekPeSsxFmuW5GfBo+HdT0/Wf1wNu4/oaIyho4qn9gjEhi
7k5f8fHUfhBWBghirToJVjfBuEOCpvx5zIReIQbczOdbzidflMSC2FQDCpy3I1cR
hsbjCN8VuNWW995Pl8c3mU7UrYBMErFKNzy83bbMjZsJuYeQKJXj+Xl72t60kd6u
6S2Y+I0hNbtBhJBHcEC32MT3yV3jL2iTonOW+35awPoDsaqjUPrKL1DxyRN/5BNM
Uqf3utroDRRLZ2fF++tqqEPB7bmD8/zLyNFIFW6iFVHLIoSy4VTUIFWBWGlfiQZL
nnLotz57GXZZHk5sguOpIfgXN1n/85sKffBQynqG+b+F10kOnecGAKKVI8e2sWbh
0KZAhQ2QuVVZ+tXYDNLEn4hwVy/PCr31RT/lDOf2Q2jGv/pkEZYcwZ0DXICBO2Bf
AAfswCeBoIpIAxQjVAZM9XS3+0vD+EFr3nskuXpPs9iep9J/u2hBwROiaRDIprI7
dni/cPv7usObalXeSr2KNOAkrchQpp8uCIOHATgiyoqTtsE/nyGm8aEYgwiRIJXr
Pk5q6jnfE5p5rmKNR3vUZV0lo0uoYtpTM25XJT9iFIG7dzdy7fQNIwoBuQNtyQQs
pRn3E/k8fjHVDc/LyB+SPmOaypSqOAkg/JUd30v0XEURwNU31PlufMsmrWr8+g6B
46e9I2HoZNllFnpVsGUY5ujw1Ra+ji71aNnF1URW1DTpLCI1mWTTH+ajlP7CgrTG
cO4Pv3SG19uHx3gJJduEKITwAFtXQeEdx3STpgEkMaLrCZTIYrtz2ZdMOtSjDR+h
fr2sHOkYk7/GuffV9DdJ6G+WuEzaLc7cHG/tW+EEaCOG5kqrCpDWC6QfOHwj8olK
vrkA/aXKk26N3wICsZ0YjOUlS5esbtF4Bk0myBZP1LVhKr4S5Bv207HohVhRJgpq
lUNaeIE6+1AY1iRLmrbHMp4KzQDa6KcU8ugPCBrKLwq4t5kuMivm9VJNNdXgnEer
VCM4hRn+twESVbxvfFcO8xoLJSN/guSs23g7S3Zk/aqjt2fO2we7IKNoH8NiVYE4
UinB9KzJ4q0OjEMY4txnELJA4r9pFxgnPPpB8lV0YzJP5Rsme/z8YwVA44VMbSWj
oDeL0W0e829Ts+bzYz4qNEp+2XhPxqH20C3vaRCoRgDU1GN0KPbK0lTfA/4N7VnF
Vq/qMbg6JQUwkX5bLhHjA1v1vS3Ygev1GMeA/aRDlKXfmnnKTiFYDqwohRAADW2/
4hQ9WchBkfVs+kxF0I3/CpPdqJt0a1n7rIdGPQTWTPNXL/r4R7BXY6Q1+YOfAQMF
iuzv4L2YbBQEIYvdo8XiEsycTjXoJYeINYjv0LxWUyEp70fIogiZZy6gdX1RsXMi
gBijNhP00E1QmkZaFxTESJm1gx7ZhIdzRe2vl+SV99Ga4T1pvkvjeEtE0d59yQ7K
1TMbqPpB5dv8/bY26CWvpYnvAwSc0rqmeZYuaeCGU/m5P52DGXbZxei/mwDYN4VP
akDu88nJC9+1vtTtgG3S3ttJ0lw0vISjihteE33cYI9MOFnbUte92UkzP5P96p7q
5E4KkM4Nm+loAWdb/YY1eDquBQPdsTqjZLGTGHHc6EQAj4+ZBJgp15XcP9g6z2Rw
/RnYiu44dL06cud3md6cnlptXfPWIqZpXqkq5By5SZDP/nbIpgx2yPkeYbVhhAb0
nrus5hYJvvZGMTMvgtz6XgvaDHnNZG4sTct7xP8gA2I+OgRp+5UBSGuI2sC+veb4
YpL/SsZmq7MvC+rOWbky6vXfTKgAvblDD5ZLmZdY1few4eEjqG1Ve7/2RO5f8Ozn
P6zYNm/vrFqXUQ08COYvGlqz5QJiKl0vcDI731o8BtsIMb2LaRQxXKGR5gDAckCQ
gMzAZkqVovkR/ze/bcRqNA/TWJHz6e+LqZs5rMOLrcRgC3RQF1njyEG0gnmQUwrw
b7nWWl6c3FxuDuPfMVvIJhpl/KMpr1G3ssOuXKSEG6O5j8Ool5HkjSv7sY146E5s
ICcZg47tTH4+wXWsRs8jUnKBrQhAOrLeI1r1VxgX6hH9lMj9SWexDntCleAeMFpz
IpogJw1LlYCEopZWxpq93B9w+/uZuMgMoMI5uiz7KESM9FP62aJRNf0TbTGbuxQ9
k8vXJ2FnJ6/apJMWjvuQZOV/hwvPS4VQJoPlwOncPzDq/9N1cBJld6b2y1hkdVQM
nWPFT4L9yJpe8B1rHU66UH2ATjoArnzY2qusgVZG5Od7il/NfJuHpiLHTRwH00+E
Bs8t/OWClesTaA2OPyVTHONHWBrgaJNp2SrcRIiN5NSNQjll5pvpZLdeuvG8jZV5
YDSbUG7QgmlsKOUDSPWvh8r+4/VpfIX9MZorIdYP3sbmXyLbJDZXCjDGGNHaBPQL
EQIsfiDhdvXypgySePk8putf8vnNMMziBkjoiNAMwhQqXKOUoXuAkpKc1KKPyf4p
kra/9wIhSOy7Pm93hVeSXgV8NA3zg2U8j6kpL/FRhzE2EpSqEl/81bmfHX7rxaAc
rmAfHl4vGz2mw0A/IYvcpcIwdCPJeQpZM4Dt7kBEEU8DGB/iqiCpHxrivrleAu6Z
AL1NsHNHvK+5pCJus50sq4srCfU977fFJMZ2/NT+gNbApDN9tSJRa2bn+WxjcTsj
0nyGZfK26NjLtagBZfPmbuL+sK0jxyGWyGiAMhWqdIKtz+PihjQrWSVET94227cw
IPOB+CPnBMKTVJUq7kekAELVWBfstXQzNch5vvmH/cX4qMR2UMyi4vNOEbarFMp5
oT2fplUDJFgRdboqv8GKr27e5Nv3pIDgV5s1+LBJELIQuUlqvZLQMXnS4qH39Z2/
NsMopYeeznAHhbwxU0M+VlDRwrFJK7Vlb71Q4zUdOrKU2zLvSY53SnREJchFKZ2c
XVUYCxgrqYJq71daYz9Y1rjyoU51gGx+SHz4Y5AVnIY2PRZL6mwJDuZ4X8sVubGv
yc3EUcYFXkBowuNvYmSOhy0CWx10EchvCHmOe0QNh9bQLkZrH3D99pg/Jw6L2jyM
SrJCc2mzOXu2qnjRgyIaCpurMNpwB7LDzVHz9gkExdz+Im9inuuTim+1cCN9vOsn
nKF0d3/uTGVtgTpBGdIqPPwIZg7IqRf15Nn6VTIN52f8BHx53OAfEj+ZoPRezFui
TtHuhnMDbmQlzLMx7ELIewHc/eKgOcTRM//qsoahTmY91JvojS3dadButyxv/sFd
YpllVQlHZYW7DPQESNcvN0COUCF05/xsev2zRtFlj4081Sz9JwWb9mq+uVyH5SYY
HLErZIMLHJpo0WxdF+LEJZobno5+gjhIRfI9sTBANhbgoRwIH+8/ce+SxluvTVDu
NzEaF2+eOXxM1JFoLljC1PRYr211pOY/JGXbiO9hh37ll8EjnoxF6FfgzyUyk1qa
KtuJpD8OKRTNbQgL2FAIE86o+qVnkveLYAGGeU3ONvPfXoEAgXF9sbl7tV+bvPtg
vL17sX9RKW46YlhYAhBmSGI1PyurAQ5ABldOu8gKEwSqpwOVPfCnLGIzb7HEe5iD
rVvlTczNogLAm8OCozGMKJrecPHO+Mhqll7JNLhbTY572QUp+IKJlgfUO+sG97oZ
BQAmjWxXFaJr5yKdefA8qjYzk0jJMGwbt5VhxIEgVXo6z1HFTJ0/7fjYZB33z7va
wqyCMVcOvj0udgj/NTB2zrj3ZoYCpe70gWa+60yve5wdwlP9yeEIZ8fqDTl3owNt
6POHcXGUibmYcV9ionSud9VlKeBbrQfk0MZjWLMVKuPVVJbNl7MIsHkSsFTRCGcA
nk05+JLxjxfc++ckgXtk8Q+pGvfjX9YknOUiS3ePN464pmFT60QKUWERxNuvMUsv
eoX4SCEYsSpbHvxDY/bKUZYr0AW6j4QC7vfOOIKVvzocQH68Y+hNAQiwn2meQpOY
nNGNZUEn7vBXsuIwjXuSg5SjMDDp6VeskLn7nYZkNSrEbGrDThP9cfsu4c/oUBZ2
d+gN/M9l+X+KIMedK6W5VksFpApfSoVhFLEb14GZBTM8eqnPB35JAUgIsH/EK+DN
vjwSO3k1OUyN964shVeJju7bzSsPvewd8REwXU4mAtq4b1t02IAGc2amLWtEFCal
b86mzLZ3x89YwbpQtvNpkWaxWTzWOJTTmzEoo4UhrKJsgWhLYS+a7i7B4sezl9uu
tWpx+BlbRlVmkEq1hrF8wruY9BxrvbV7aGx/sczS50BWBJbVEV1+QMpcPOuU7TLS
Zvk96SQ21+PirsnzJftLncxatB2advvBVQGZWkd63eQTsPQFzFqSqH8iQ9NEWZVj
7AvcI4ARKNO4VJ1KOSUnTPZLQYm6xcHeIh8IOkO6xkqI/eGfBqjXBNCNQ7u78nHQ
w+6ryb8AsywAZJeg+T1/dy3caREY5Zhky/xa/51n44db27KVliV3YS8jeIEH3/00
BkLhapNYR5BWPW4og7CymR8M42RZtS7ggmzaRTNKIz67tDwBg7DA5Hp2vLXFu7Pg
AGMKfEm3DHVaWEzMROajDE2TCXO6obBcNZVX8nJGMxKp8M9C6d82XoRWt6D/bSkn
tZ7QNDjOB8Cnt+m7TxJbs58Yd4oxkYq0odPROF3Kk/eHVwWeOnnM1V3Ydd2HUQlM
18Kp1cs/suMJAwRBuTGqKxUCV85SLi+UUiTksuw2nNlnEE74icsrDRbobGXbAmCt
yyVC+biz2QM3OPq3Iv4gHiZIk6GULXtuXwjt8OXAfinsvo/ZDy455/RzBAsnhazW
r+2AA8+sXvrc4i0RctsKNEn9dCTi6iXdT2yf+IOoHj6fGGaHPFuP2D/ubJkmNpoc
RSmwTArHWFrOorHurLyOWdAZ5oS0mkXqAr/hC0WVU5rk7GtsudyePVyysO0/7tlA
nclMym5fD2DaZ4hZK9tbDkBnv70i3wjtOhrmrgvwE/NFnlUWr0W4nvQybMILnKku
P5+r14gjHC283fxiaVpf5Yf8212LnY6nNiHSlzwUj1FP/vTXWTHkerndT9F5gt7Y
DvfO6qXvdcVllbWEULknfvFYOVJwHRlJ6MBP15aUClJ/66uoYANM3cbX55/FIJsM
v46Z7CdxnWmV4TDQFIT1GhgfVTxgWjw9SzQi/6L5kgeVzXhH4zl+pq+l8qvL14ko
HqKRMOVOs3dA65PirW7Gus84NagoPCFiWAF1qmLbQAttya50d4PPJTrDe2T6WVxV
iYQTP3ZH4XYPkWtU/uRUb6BtYdyJrayV+yAE1F+bp0YAaE4q3wuw+WGYw3Cx8BKX
Jeyt9Jcli6Uz1DKlD2ZUw838Y+NS56d5UZ2NDfpKeQ6MXgITbSDOXqPu2T9ZTb16
kJlI2rUAa8OK+UBE729EpRb4ff69fowCGxrMFwDvIQ6KxdEW1+RU/UtpOfIYqIcl
Qk3dnLLfz+PCPvglJdkALGbl54zSgvxJtsTkY929Ndl0ApTLqgRwyriaUsZCFHZS
9TQShoX/HCiOvb+bSp7UwChQuSykN5ZN6+PuXre84RCdFwCR8cpeKF+gyNCzWu1u
zmJheHPxmo49HhffWoE0B8Vh5Hy4QTE2ZxILKKMmCZYKp0TZrj4Ml4fcdRe+zeW9
3uZAEhZmeEhs7hUojQMinz0nVxidDwu8iQsZTve0uOh6sp2DEGjyKm0Ou2TQxrW4
VIcQOfSGYqTVURmDcTj9XtEQus5Jle7otHOEp2FcMSinLo8VFWodK3ok+3SCYf5q
1v1/HFxpwXrMb0g6TcxhVBOQZcOmUSG+xEmZDOraMxLDnZfY12IHWQW51btG0DEp
x4R2h7tjtkpFPzmQEGhDhYZnDlEg2zBPefuIxzLdGxx9fKVOZhZvvp4ffFZp+n/R
jfISKZFzNLVn92AyMe1guFFOc2VMHsInEjqAY0D6Hbeoa3d4zxiV8bPKgvaBN+An
r7U3AL8WVhdvaIwaJFpoEz9Xt5wYDkb3DnFOgGZw27DW8k5hQ1bfRtVrm6RSB5ao
tPZ4az/n6psUzlDWg7Wbf4klyBDqJMKm87dQOMWj6kglNAm/GDVXhSHB1ci7S75o
jd4m00BisXrJjYzHfLNlQnrSrWmI3aGfJsPBpxxGkqXui2aj5O6udNewu2SUu60J
zcSKiMpEktY/YYC4qxklGKZ1gX9fwufVTDLo6onMnJH7mCRDhFGOqN9b+x952bH7
CCsj8QEHcGySBNS9Z7aub+VShAGThPGcYeqZDY+K6BCh0B0jTqfsfZEyGSUtpfD+
6ah9TyEr/PexBx073Nu/75XNHuseSohDIJbo1HovMVs+9EgNUsEBqfhgq4folTgt
ci2j+tfffYgKrryXqRW3ffy0joGa7QBtpXC//5Ule6lhDkDgLuXa+061CO8VwtJH
kav1mRmagRDOosjjcB9rRG4ADekZ2q31yO2g8kcSFX3W+G4U86BAIHoKvU+NWeNW
+0RLyW7m3o7YD4v1ZMI4AFd9zvoopF4slU+9ijNsCX+Ji7Xeb5KuOABfnXKqGi0x
0u17MsxH9wyw6qGcRdR8CJmWlvophzWnOuQAS3MevGiYH2Lo8IdYT9zfu+9vZlgF
E2qQxGczIgWycv6kLTTIDmTq/hQ19zYosM2sl4UeIpLxNa66M/oQIKVUC4GT8Fob
oVvmRhqGpfTe1Kh2O0rJKpuDOtkKahQUEPERXyD6wBQR8+YGTzGW1jotH82x4/4I
CnCv7EoLsJAYKvVdygUuXbv3RmChhpJuylyB7UAzyniEwGXZgDxIZO7UTwKAE5wo
C7LAofxULYEEOjzgtLykh2/KKyaryZ+8NQ6RcGgtekhqOBpToRUzUBLxxbMUq/8Z
eGv1gtVSCKrP1j77yCuNKNDwPgLOlyvYe5y3pkNn26TVf+qVipoc4D6wq78aV77s
b4lhdeyTMWBBeMydYgoO7+9g6UqT+vd6MCzQB14Ub42nWH5HSGfUAJk1Q4sawgUw
aj4tUemqlJUaPg3q16FMqr7JixMYSfnnvsMbwbY5alBW7kcpmVjMCC+r09wOVfFJ
FjloVJ4QDdCtBmATW9cu/XwJSTMwtXRWp64QV2sUjoDddzxXKsNpJoNEY1+bVlGF
/J12eryAV6ENtRyFpglpA8GLQ/iDjXQoxFBqfYWU3EbF778OyBjO2cVGHENV15O9
3JW1U8fRwNczDmNjsM7xxZBmIXFpWzjLBiDB4+Rm+ax2j7R4Mzb12BZJGAaTofxz
Y/WsAWJHu5WEv0rKBcQLHNczzrl2PFv26QGolaQphgpELJLJOGyZ9Ec3TYLlCt2i
ezZBTMjCF3XVhfxLB6wetE+GvhM/1URcI9IemmXEbkSxnMYyxDCCxsnhhjtVk6jT
V8FCrJ+hJbyiKrCMxtrY+dkPxLEhYO59/aq0KF11/WyJaewxdNh30u4wWJxqPHI8
8Lhi26YfJYuANDRwVGfw/8vf/qcc0m0XapSyOhMOe1V3Zwr6nckYEckXLdQLcK4U
k7qcX3dKq6lpfL59f6Qbif6TkqSXuHRtoDTEi6cCWiIQTySmL+W/NEZI9hW6Tni9
gXtjB7IR/1xnXiI8foAUUW8eZ0NsY2k9gAeNsrnZAjIIHhBBHAOUQnhG9DXDSMw3
E56F1ivoSWNkSNup81mTIrPOQojrJBg9dUdVR4WBDR7hrvPedscIhLwYvtIY8ZZI
PkygAFJoggaHveCi7PXKuak7Dax3euoP55yfOLunT+Y6BjccaBdQk8/bZ1LCtzly
4KuBj5u+WFz6+wmLuKglI+9QVmQR7Uf/ICCNAbKrsf/IJlXotRE0ZVeClUFSDwue
yKURu4pgE7yJwU34iIQWlR5TOtlfMAXGP/7FWc7zn1/2JV/1MHAJg1J2zxAi9+cB
omRaQnnXvHk4Y0dM3zl97U7NxeckRG952Z5VIa+Jzjl76twdW8nik5M6wAXMZy11
IrCbxKbLU2oIxLCVOajobqg/TCsFQ3Kwdw2YRlQB3jqVBwIcM0ag9CjLwji66Ibb
uRX+rCGxw+HwCVkKDHGY4vfGtOVc58mACBc4ppWWQGfFgi7eRbOJZ70FdvlwKd9I
5lI7I0m7j5lBhylwNt1jvrxAgMTmmaqRxYQjUoFQPwukLDG5yQ0c4yk+tmEXkd+5
qsu5+dycr8Ci7/oAE7AgVrNuCmOP1+8jAUAtljbkTKB/wWUYRdl6PBadSM+kF/My
OQYfUBoNMxMlalkTfVIB5euV/OJUNGCjwFhGcixhwxpCR7pcyAjxtXGMho0IIg/D
efzufpo0UVcdgvEHaClqC3zHmw1Y15nffk02OFkoOw3YEubROcHlNdjJeIJYydDO
J/T7ktObwlis52Znhmv6mjKFy0+uYtG97+zxk85r17RqiSYp/X6MdpGbNp5NrsvH
Ila4jzoiFdWAo4bG9Li33PFnQs0UYyuxnzqVxolWII8t0YAqHXCSQ6J8+hugoLml
Uobq+F71LpaMgDOLAPCGz9+Ag8fNuy+d3FerfNA5l6hu96dtpUhgCSAkj6eKa7FP
wqUJrsIeUPcK40k7Q8tFz34z/4A6XVSkvBDf9y1aZGWF28Yb5IGa5WnGNkgQtNNb
ZZ9Yh5JAFIWO5Cg34TkNDhbbV03TPqMQysk/ilDxceBRNyWyYDynVi2zEcQDbYh4
mf3kGFHjPPTg7BtfyQLFChfFi5YVbCP3u8t384yTjQ6wwC/QR4miI+/ePU2HUE5Q
HeqHZ18oydXW3lxWDm7XP1azinItAfpmZy/H0AUHzlpBytYFRON78iH0nmezk3J/
HEOO6VzILLTimKRJWlPKJLWTZ7AlfZOP/QsAHQlahwfXaD7Kk17GNw6ZP3oSHupX
LXdianQJIUlBQRs5zbOngxfZyepkncrf1BuFM4GDBnEcQYxSJhD02SnHZCqFAVol
JAY/NfnyOz2tBjycDSp3Ct/yNJKG+ce66eOvKfWfb1WGtkxW2dGBIN1BCeHrqYOH
5pqTLM7qKaKEyNTTW255z8EzaCs4TK08M2Ksl7F2m5wQXLdB+cxVUuh4NztfIjTz
NuhBEp7jSnP7u2RXjXnZZ2LGPm4s86SJ09OKL3bED+3VdspqzqJlObevVTOaCkSX
V5meP8BfDneNqw3pAsf0zMIDuLnB00tb4NMuDcwTQ75pVfc38K3/KV4k4sh03sCV
seAT+NPpcMiu2+9/U3pqld8vfEmjnfJzlMJieeS0N3RGBeCYEgncKqKVFHVoG/9a
uizuuC9dd2aOwtNMwPOKzyGUDtBMLqAtrXLq870q7joDIdVM+zHCNDrTP00DvXgw
SlbN9xK9Z95kUKjj53atrrn7lMheeYIDELRGD6kugcT3dGAmLTEl1jnKpDZixCnU
/LTJWY+H53v42TJmFBiY0YSL27tLkO4rYVcpvYj/mmn0UJZBHG312ax1pC65zEiT
tk9FJ4FNOC41xd6WX9lcIgtytSJyIbg6kKlUKCZmw1wdd8cL/VDajd+OyJBJW2b6
hvdJVD0nnDVebIjjGwvnt6F0g0BvZoD28Xr55xUgaDUuYyXY8LHa0zX/gTSVRSL4
cKQGIrib4iwOrIS8szlijWRlHaILt8PyWX8N3g3jz1OhQPDUcVSUrSTm32SUbX50
A3c7lS3xVnXXvY5w7Kqq+7+Hn+35GuPvRkphLQkXuqYyvJ9UWcNdnFE17f7pgNLV
NcNNBOGGX5hHNUXhS2VSXIOUchTI4yZhuFksROSc2FemoxHNm46bQ6CinkJJxXcv
TnxxYXNqYQrtJhF9qXwQJmaRQ3SoEuIa7W8hRjSzie7ybpdGdwySZoxO6BT9RhaF
ATlKwbBQswVvQLJW8QMpzxCbEKXNpt4SMXRRnpDW5zKR/sGa4OMsryynTGtB/G2t
3ycY8x379EpEKLib+xc7ecWAO2alqMi1GATGrZ5lioKNDmQJ+4HWwhQe310qfQV/
k1CY5vkcd0jU8rhu0Q4fg/vUjcgFUd7RasDB0hPtWk1gsOJr9Rn7Bwqhix5c8GIx
rAMMBbEMRkAnBQtFyhqschhWkqRR96O+dhKyBj7sPavRJu0Ddi+AEwseEeupuSp3
GXR3UptzhqrAIAK5B3kAsfeSFaF/gW2jc9bacN98CJFdU4DPeeiv/xCieJ/pRW3R
+704tUrlKp9WBWFK1Fo4nrG4BCaeDkz2Uh8KRnMc+7L1uo5E161plZQingVUptKC
RH5xcYNKcK94uTj+LYGYNiy2cao94lY9I4QkxfbmUkELXDQWnPXSAaYgtFbdg6lV
Arr/o455WWvirzZk+XlfO8Fm0z1jD88e6C9S9+g31MAsftyZh0A68pfKv9O2E6Rh
d+J/WE8b+dkj96oVoUlseJ0GFqmsJRNtltlotToHjscbNMNva5FIqXzngdV0tlaE
MuEIBKF+cTMOdkeRe0L5hlMTNDujlytyjIOEcbfk4I7GjrWQmlaHJ68Hzimno3xM
Nsz3V2h0O3r4zinlHKhY/1haUveNJuRaY5UAhvCDh0rZwh1Ll9jbBqhEPz/4ZVun
X9O+MbBZ7JV1yDb/QWVoF32Rf8vYZfs9/W2C64OE2YN2tV16pUZm+C7O/ZSsvOC0
h+K026gs9ZvNxoFIprmb9KrfkE/17k+I4dH6v+ONymtQvdVNzTIyj2vx3gv+wIor
6+xVepUd8BXSQajVCQSTRuD4BDlDQka2dgvQellavem/djzmm08lKpttlIDUv93O
RZIEtopKGpM7P+nEN8f9jpoQcEzqj30mZF/94OK9q1OZRbTerswm/3v2gqg9umOV
TJoVBImfDxjT8wY3GmCsUzk9EzYWc3XYCE8PrrByEiqy8cbe2B+pZFgdUTqAbM0O
7bEZAasIhBq4Grb91zPJRNcUfkbv2BlwlvMGRHnKxHI7SUMQVZUVkCk0Xg9rydbW
n5tHl6ZIR+w52RaF1HSbSZ9/mATPfw5ysr60iqvfxuVyw82+YsLnrK2bGIM7Tn7k
0jKuO9JDlzZqWqrVIAGydIn2xLsv+QnefBw81p7fd8atqaf+OjED6Zby7oZVaC32
ku4RrnZl1SvuF0jgA9/Ovwy9Ddv4aQ432gIvpzpOKq45inKNiYsSpyGAbysDL0Jq
Nbo6T2HYYHsvRRIjPWygaE2ugnVwGWBZdR/0QOSi3mfm5TbUAsHTjOpeB+o597yy
etFlDqts2wZlaInNwrqNYnPdHGkxU3DlW4Hw/pv8FUL5yjWn28Y3M3cTex02Imtm
gHtoh6VATuBCYnO+ek4kQqNepaXUwiaPcS8PvcanaBgIQn/2piQyXfqH03qmevhD
uSPwbPDJGaSjvevcyg9F6XoTAaP3vo72vMErW/03fRr3WSuZDc9ehcylLczf4ro1
VnT5OE//1Q9RIGrAHNMqgKcrMxUi5hdbXtbKxzg1FvMCsu3QIV3+2vLLnYLN+e/F
q9YJtW9PeNWrUBB4Z3eHre4rXVBrHVQ1/qaDXkxb7k3mf1K1nrRR1DFcTy1CNW69
Qe1nUnYB/XxqyQL/TG3TcMdJr5Qw8/LoggX9ZoS6+LgBtGw0xazH3nqtuiE8/BP4
iuoqZjLTDOk0X794hM+XJuEbLhVgojLU7aUbl4faR3JdUlcpUojD0LYtzzLuqMt5
i0rop77ZqVVSVRjtKk2biPYGwFKO/a3yZnqVCPwsPCsRAWgIM6ReFq29mIjo7qLF
cjZbwaZcSRW79VdVjuLJpd5uixoyI9R1f5H/RpWf8R6mypOyOaxzJ4Ml70lCG/Vg
g3Pzu4loqYQyOIFn9O/fdzivpx9gSPHgAMSF5YN1LlEhvbe+a3kQ65O6IsHXpeIS
WyUM2IOce92DdaRmYeimxUxCreJ2MrspM2QPiRRdWPvs1fJHNHSPUTsv2O4EgNAm
G7Nj3KmA1jQdOaDYz0EQFMRQ0FZz0IK5ix56ff3Ky0FTQajhIUIpi+eYgBMt67JL
91J0mlT20BAkPXYp0dw9Qvdke8xLFvIWVoQwTXnztKPaaUhOisG7QCHkCGz+9CU/
0bqDSSrcXDsDfFuTf9YB2neohm76qeEM4MwG8sU5HYdu4YKCE3C8Ma2VVvQxYrnR
+czNlP7J+FgwCyGg4c4gAjPoTMVHzgPIpuxxkQNmJQ9m3Dz2X7o7ks+lva4I/P+b
uy4xOGJ9Yr3JXoy/l1p/4XcDVZX5UVaAoPVChPmhIrniGFVRdu0W+Iufkqrn+ufQ
IoS1br8Jww4jRyRANJQY0mChE2r/vBcIyytFhCmH88OrfSXnQ3rsdkZIUrxOhEX6
2RdEvUpvBIQq2wNB2o05vXmQCLIs96bobVUvvPRvKAcVdaAMrfx6LS34UlAh6qkW
unlgrHccCSqKxsOP0TCPZVUkd3bSE7+3X6+9yjpfqm5w1gKRktCj4lVkodAl+IB1
ZYbtpqDgdOwG+ivFFsXWspwxCtM9P9kot60vD8CiLJKqZz7Kk0M00059Wk7WYX9M
NbtjqVK0B0ILGIoCcuaDP/CVVlyyPj8Gw+dCHqEGe817sOWEtmWsq4C+Nz/6k9sr
OUzJ6R4QWaPsSaYZP0hw+i+9EYRUZglxE5rwB5kJ2CKkBJu+Il5mAhGLwaXFD7Cp
Xjm3Mjv1jeEUhML70CaIXd7qfg4mk8DYohs9ShjB2PCNA8cLSZK3gc4r73JAcYTs
Nl4g36XGgQGey8/oEmMGzgYmT8AVlQfcro9aLbCv3/epXL5t5dkIN9OBz0tDjAjA
ZATciCezMVt9GYBR/TmSt1cZTClBDrWnTAW7Gx0cMXbOmvucJO4mX0/U91/KM2y3
X1ucavILCIN7MudUZRwqVJWo0pfwOrwHLWyRhz9T6YdobZbjPHfSqb1HhpTQ/Afl
NZfrz6hjnSx4xV0qlFQ8AMRWHPsEoxbQMeEnBboVWtEubr47gxOC6/NWTq8r3Bfy
WlVTj9RfH4Qn2AUHD5XhJFCjnAnJU0WBCYAQxj45Z1le4wpJ9cPGTJKEKRArvevG
rGkaWN2VRaitJDaKuFedzBz6NMiREImtBMZ9X6opcfFh39ijAYLyLl4MCqPd/mkw
NwNUXgFs2h2EQ8q6SP5/IX69yWVop5EQynGpNF5EFTXBhWLjFu/a1iK/gHzTk5YU
tRAI8l6Xn7EVHjy2u0N1ajz9Vi9Yv7E8fXEAhjZrJGYGbEtdebyTz8CmESbqE2zF
J6nvfWNrhKmnrro8yS9aSz30yxaD+HF+7FTnzc5UC/I0ubqkJkHC6sNZaFVnlAjK
3r0f9Vi7HhEOcXLcKaWEkC+C6lPlaJE1oRWhi27tS7iozbpQ286w6kEuSs1gPiol
lUeK4rvbTmbSfA/Atcjj/z/z1va2z23CMxLQc9ZK9OIqH0fP8Zq9XAMBtSrRN3Ee
n2B8sAqvpmhNqAxMiDWPrEXmk00gPemmB8cxNdsqF+QyIj1PVVFOzv9pWnifrGYO
2hok6W5bQJlSHncroNscudPypkzfJgQQ6Zq/hhiyH87Z1li0EI7F0+uW+PSCTjJW
eGoxaYkGKiZbpQB/3uLltpbnlj1giMEZZ1dFxsx/6q7TihsgDS8UmvJeJzNRBvzT
Hx7xi+tQUMkM6jMblO4IV/RRPEbRu69LXRzmwEq+IHFwAHwNQHvCC8vcMDwmW46s
u42wb0NddrpRRtv8tRR5tBFKvnJrts/WcxA9jW5861tP71EY8gOvyQZrofmMMr1v
EH634Qdy3z1PzQS0tBhRipZcQkDBRGVCNhYFxSObGTL3OJv3bP9AhrAeN2qzJrAX
Qo4DmQ8XAgmQnX0IGWKUEw4qKWjidZF5RJ/mrX8pVqinYpH1AnZOvtNteP4iR/9r
XDK8eNP6nDWPmV5myyDhRcoQJv6s8PRcGIdGTV1wMszbuEKt/IJiXq/Gy9t2Fd+U
NW8GJTx7kP6+STXaplA2rZaW4DklS2Xe4kcTPzJ7L9IgJcYKVahWUiem5gk0qIgr
4fucDh4iUzW3OEUtS7F7VVATG6pAYGsKYLlv3/r3qwza7BZTttqfnQkP7j5YN52i
xb+BJRPqX3h0rzrIh+5MM+1qhTJqsKydbB3wrVJYpobVKD7JkK3Yvfdu0MbDmyXU
q3gaJ0lSTjK1olTS/GuCaESul/zklXsj5A5WqgGSXJ//GfudvFCoC9UZGU9xDAix
IaoY98p8wtJSZyNQ4HxvdZkEGQRAMYl+h/WDYJqw7AlrpeXhawdVpQC1v/NiuC9z
LaB22in14pA31InDUBC8X4xRwp3HjSR1xFDx8LScLo8Ysiug8SdDem1aR6d1VyQS
K5mp2/cn7GoROtI/JLNlzT7XRiXxEKSr9nIXRK06CuWD3q6OXx6izkzWFXfik/R8
AeYU4nilGybdKoAFzmLmZeQqG15nyBaISBcXayOeWbgO+Od79VerVdPLZGQNDcao
hqIGs1T4iRNR5eaJziswxMbmNeReuT2ajJbHFGxw8nT2cZVxJaYstoQTqj/y0VYe
zzS+0/ZO+4bfpr16xe9A82NOVA9ex2wWFNf0VcwBGSHQsUnf3a91sZYU1WEy/RVG
GtJmgckW/JfVBRaY2Mc1gq7Sl6TlIu7G37aFshho+6E1ddH1XYTF6ut74ACvr6hx
lo6ZGBLxhdS2rLRavw/g6oVBzla4dmiHOBlAFYwOrfsoedo3paZevrgGa3hgs8Ku
y5NA3QBJISAN+aR+kNb7tnt9bBsnznSwBVCBFQ11asKE+tn3v5rcSTn/WLyV7BAX
SWmHNeolLdV03E8o1tqVXd/LYJDUDYIgu97FwHhd6f+7/2VGao2T4HdVYCblYzzJ
xt9mVl0oPePMP082cmD4XbnPwi9E3ag/uchrThNXsvXjwq9QAvsEnwNwMQ300gE0
5nXNvh/clGzMg5tixw7t+mArrgSVeM8pi67W3rHhJva06rZW6nM4t7EAHK7X++mm
tcfVornNMfUkluMaxsfLS0Nqw68Rx49a+v/v4mO8aj/OSEWcc+aQeCl6GoRyH600
SjFgDbX/oBjxw1xVq9ZxT+GZo/SR1E+Ndnhl+5u3JL59w7wh4Tp84RE+1E/mwaQ5
aoewTgSYLi2MofrAsa/oS/TRBR2k2qOiu8iUCkZiV63eaFhGwWHcgn12PqZX94N9
XupsA8ulLPAo7TZOaStuSIgVw5afvmQMVbwuUW2AXZLkL+QbX74KixpVc/uoiUbv
dm/wCjs0/OCCaZFpUusP83aEMBTySecefhgiUWUiUe3r5B5GIx42ELb/ugwRlp/O
f35UtZ2qgaZmzA1x25NP7qnVoAeo2+y3ZH08Le2ekB5JGwTFaWOBrYCRcubGqKuL
eb58gOu3xkDDq7kwfRmwohlbDUJFbkQzNexd8vuw7eyY3Rw/HYT+fYin/0LBRjC2
uOy5jEWZAPM1HHLriPH4o+QZBUY0U+FPX+7gULhotbggC3gD0k2fxK5ijSt2FMtZ
u1350vHlGFnwO8j5AUra+M1AA9Op5/xcGmMoLraax2YZxtukAuWcxbCS8Nb8M0EB
622NUMAK7wf30vD6RFjdKTyZWXZzcGk5bAwEIScfYoH3QMP8wi8G8Hhn+xD0b2ip
1w9GcnrviocACBMFdEZdajuLF5zZqV2BacvLb1CrAdanuH+p13zzmITJZO1WEMPV
QCtDRSMfy14SXvLRFih5HGvNcZV/6EQpry2C5x0lWqqohzFvMt11mXgVq5Qw8gV7
x881QlVKDLfSzf4TPCb0W+nQR4lr5MuPvdn0VouaUkmNlCQ3l2N5rLO/QKwKAbIu
ln3RGhuh0GA7kwuF0Qe/4EnV1MSCJZm3Jkj/FhoDlwc07PDKiomZ3LUPITDBGW54
ccLdTuDjt1KEOb4AGQgg59eeHjeY7Mbo8dlAz4XTqygX+l63MsVTVK79rVifX9Ie
f8hINZ/PmNqs8K+GgLUUzd+0KHEv0ysYt+kRBZyV7EyppkOHnL8Y9ojNu+5d/JE3
DlLOA0AI62DIyNjnh/lr77f+KPJyVxBuaGbhhu5QuTE29TlMD4XNg+BgBvmGVeWB
VWoU6p9SWkKYRFlbzAjaDbY6s/fMc5pG+ebgDXe5d6Yi0ldyVfqEEGtInWMz6mJc
tqQXxofsDw1S6Stsuz7ChF3ZFZzf/aU1lGUI7BlQkCgrvb46MsfzJfwG0E+Xwo9f
4aA2a4GM/KCT0mo9ffnTN3Ic88yknFl9Q8tsc9qy5PlHDqb/Ir35f72ObwKBm3FM
jrbnmHBWjysE3EXqYLHFcfmh3B5icCwXgKf5ASZo2GTgyDvmX20//KOjqbfWvofE
pJG8HWdhlnCEBPa0+X6yLt4IzveRiBYwvZXY0CXZafHhforER4O0aGbyHoz+mmIf
RST2gQgefNMDjGWfxrEHkbefyLBzw9sQ+oZA7RZ+OxUYxvCmJGMhBYwF6b5/FfqV
S7oTxTSSecPhXQpyGxoGvkx8Wf9jzpooyerzqkt31pencKguUeS4JmxUjx3Eigkv
GcciohIaNWFQOtC+jJ6luGZq/VoSWCVXK7C1X5Wf6C17mf3Ast6BbDlPE4hn2ckS
MuythJqNlreGSk+yVF7OVeqyeVzHKe7ECsGimMFL4j2cu8kmTm/VlEAmweS3oYVD
9Fs95i2beiK8WsbIb6qj/X/RpDChP/7wdy0ZDFoNw7n6Q9MKRpH1HtfdJ7XTjdrK
xdPReUhUd7Vb2c65rBxY04xxfFYgJoCeF86oYVp5bFozsPmL3kfWbOHkdaAsKyMC
DcFOaK5bXHdRIuOnJSuGtq9ZhnWPoJlYOxGjQmTSdkuLHmYoWKkeE1V6jopy1ybT
ymf+WvQ3B6zknU08ddEcsT9asjUVmMn2lbxiwY+FFllGXYET9ICsgf1Fs0fn8CId
QChwlJVbO+GRnTEFy4cCjgEJr8ZKbRFsz1tmrBu7nq3V79Io0zRxodglMu3z/9AN
ySV7mCci5NvxXLdPfvTmUgVqeMnmk/RVtI9OErBS0xkviEF8XL6cp60ObVSKfQD3
gIkR9WG0yzjSfeP284Lf07V6Urptoh2l24kChBOdjxDSNdurh+ZMIYMzQhcgXXH2
EM5D7FHqFZHzFDoTFejKXJmi+WSafdnGpjCwOcH5w3fJQXqC+22FA4g+ArjjuVDA
eNPpZ1UI1exAcgh0ikt3ZbOl+HyRIbWUFiNhS0jioQJLoBn21feAl8T3b2+BcWlV
VNYSznJ+VxPQ9TBwkHG8L38+Kagi4kY62GwZeUMC3xLWPH8Dqyg7lQ/BTE+UpTpA
nmKY3lhWYL3Tg7+wY75eMGtXeOKbhxyZCj56uU/yQPQIxrvf3jqAWhv+dpLQFYI5
s++GwlOJCPk693Uqr/Cz37uBj31FR1M9wTEKOmfFVjGO6YRKW6PGOrPgdJG5kgQU
JntwLP+RUDuU/G2cGzJRtORESSnkITXbOidPTADJW+lRNzscTTRGw0ET8cN75BcR
Nb7pUDKqPgcZxOGFDl//v7F2msBOZE81LKYHCDwyk0AU9dhMMgr/p9aUceqlHD/A
no/+ODHYRsU0Z2LUWS2RKJf79ZS8x/VN82Dj5QuHhXIVuBH4R7d9WahDhFxqULBv
Ah7gihE4rl/peBUlWu7GWphv1ZepGt6EEGZbpmVPaq6mOp8sSGhqFlREDvgKoqch
exhDbVDMcLYBnPlSj0EznLXUnwwSQD/al/LPT6QhdZe6PduZ5iUS39og/1hvClmb
Ef1Vdni0iIkAEHjTfoHOKLiamVh0SjAetTeu3Thbzd0Dq7XST89AZTVhcYF7Q/+n
aUzlPH5BmPVsnsbXMzXcqMIkSEfJ3I75XYgUjSPoaoPRkfwV+d2hvbiSfakueM/E
nZYNlLjwQP21oO7Xl8woqRauO8k8Ay3IvW+9PPJqIjNSnwAJ5vkv0/tYWOKDtZxw
kH4Xrcjso12AMinGUr7vPwDOzCM5FWzEBf/xxroQCmv20MpmGcuO68eaYuqGVDpV
6bpvMKDMGvcpJIeUi9Kjl5Spii71d7tDAO4tQMYm6ECgj4UbTgubXXpEsQPH0dPE
aWJ3RXQHxBGuDFSxzjBWM7qvddWPYYxwF7c8ZHzP5zfOaBjiNeocEWz61tpxsIhT
5cFjsbmhNYVmmxaFS5L0S3YOTkjLnC+qpzjTwUrr1/BOdeVfrrLie8glIsJvUhO1
hw2iACgGFaBL38DpoT06CfYMUcb4XkzFi124reLXQyfK/j8QhLaaQjSYka0941RI
5EvTPE/sM0Fg8YGKgI2egpijPNk/0kmj1bR25Q/qS7jdd5kxxXl3CbyPGWs+gD2u
9xTxP69ksE3WVYhJ7iR7ZuIik/fgyKkVRasoc/W7G29YOpBenmBnB0gIzCbPavN6
SKWwZjHxVkwi788BavoiUY2snDZmPnk97hHPdIrG5ddcozilb2ROq+93JsUHHYfS
kppXc83ibcwaawEA2lrfMYQXbsnwgK9G5hDXVix5zoco2RjXzlvgvmCsnhYMNQ97
N4wTGm24bu/Ts9VPP23zcHBnx0wtrVMHUMrSAf2DrW8kET0AAHKJkYu2/MtETum2
qZ56r75pU1V6ZOWfrTEjg1d1/DhtZXhNo/oKDz2I2c5/PI6lLbAVGAmUbkqapJgf
XSLk/LCzWuHXlUhfHI92377As2BNU0D3+1xrCPt0yWLVl5bBmclj9slQCSp9s1LJ
7VcaOOw89zOyHC4MCYqOrHBkKrWWeCjgW7j9uMSGWasmvXGFtO7dmnlGm6rGBiDm
np98JhRUd3KUkLmG5odNNiHWcYfOTHE2mjvE0nm4K0xjWNWTad4RIwn+ssxmm5Ml
Dbf5x/OUZkNWs1DqdwBKMt9jDJKh86NWb2UdChML3hZSvj+mxDD8l55Jqz6i6KbK
8dj5VYkPz197yh9Doujpan/U+1TFBVIacUYDEjMhH9vWS7HX4L7gcX8lNAr3TRzE
2Mi6JMlMpInGW1+U2EKmgZUuAHMSkwXs/e4pm5A872SsDp84X+GlMuqgoQgaMx26
vrL4haTMQRuDEWTD0ECdeegpEprQjXYLGIi6tDWOOKbY1ue6JMjXARqlOQR9MIPj
JbXCJoxu6QNNtU4AD+pJkBvZWop4Tj1Xx0+Fx8qVtC+EQ+4oRevlMmTWlsZ3ovU6
MB6QbV4oWXnVTFoW32PJHoQ0tkz4tfNopkAVjINJOT5n2cEvgngsT69yAnN4Ae7G
SvHUwt7PPX//DwyjCyWXzXdBl1vQJcwqMBkBdGth7fZU77ZDtc2JZU9MilmzAlcx
voXdTuEhwJDtQWAlNQmxjsdLtAMS7IKN0HGTtSKWYH6b+UyP/RA3UUy6ompYbnMr
I6krIpUDBC7L0p5bm8ctLZwaFljymzXa7t6QstndZUneogXHsfMycOaW8+VZYZSf
8S/VcoK7XU7sjIC/I5HvdQnXC4o7gQ12aUd54GNMKhgIO/xhVVncZmr9pxdcD4hZ
gR8d1omaQpoVRnEatISzFzQUlEdHHBo8ZcoSC7oPAMQ/drX/mNoa5R01p6etxdj6
cUy2tRyfNQsngugICwwDLO0K8jEEULnthe3tn5RJ+mbP3p4q2HtebzacDkPdhxtv
1xCim1qK7+63+j+tNUbK1Qb7r0ynJj9mnGcEFfTd3FKtmJPM8oKZKgi0n0Z0L7Gk
vgUQr1+WgvGoXdH5D7aEiLHssbs0iOXBu0fguGGrw9yST7zLTRhfCAklhJEyLm0x
tEl+S1t9ACUjVzc2usYyEOYwanj6O//NU1rhYkKw5R2pZKjTmznSdUAcBGCyKbID
51tfOtPuCtfTFGt0XOA9EVc4HqNo7C+efV4qy0phPuZuIoCA55n7w6jRBNZj0QTn
WRBAoOC3TYjc22amAhOzKg+THSgxSJfplVzgW4GdraISnbca4+jYaY3e34QRC55t
/CLBluxgDeVDokKBG0voBL8USf6u3nUYc/JAGlb8/JGLqhik4k4HE8YCCLFlswsq
uKU5hkmn6ydguGa4m8aWH5p/v+U4m4avF2Nm6XJs7/Mm2qCB3LF+j2iP1BUBmuU4
QLRSzTNDZJM9spRz+kr0DMFtEU5X5nXyIDs7hBM3O+xOdH3L+mmdjaQqh9fM3V/e
fH/3jni/Bd6WgLqwgGGGxg7qt/wPV9m4yg/6UUTzHQfrklR6vfu8nlulI5Fw8LfU
e8Zpa7mvq+snhqg1SHb94rUyDtoKyiMqeRpmbpF6qlBSG4/l8uuCPpiEgvxxQARK
OSj8ut9OQ4BIr05ZfCfo7ihl6KWcmLyqV3fxzphmW0XNyxWXmdy0XKSxfIHIQzwk
i52e2qAZEGVknC8tYIYR/rCRKR4xm3qzw79ZSYy/SgKn6fOaRPTqsaJD2thx+TW0
uALxkO51TSn3fPXMMz5AkYxfYntHxSeTFwH+2wZ2cN3IsdFjXYcqAeoOexo4uyvB
ZPRdzl/wGyUNhxd9Gj8Jkxkk0556U1bF+6ls36/WHgzdCfvlZ8h4QX/wP1z6PNo4
vUABX5OFB2EYscvTKQI7STK7bprJbvxYPYV6dyigOl2OMaVjVbbHVS07SdNDJtHW
CuAiU20XbMiUymH6QOgEOtzgEEzLb4lEtIu4xambruBOHQOFEt4iFBXZy645Lfsy
GEOGFdT3ZHRk+SFQUhwkLxlxefjuEDWrnOg9HOvWDaJJkpTRJMcjEJL/5qlFvmMj
eiOCE/OWKLVoUCmkBcdBPRxqsmfElIlTEJ7jQC3kfqWaKhzIBdnUIFEzbbjU2rj6
DadNmqE0YfwmqajPqeo3G/gpI+a8itd8vqmGzOcuXCHwQoPsjLEXvMlnIQcWk52V
52X56it8PcPHScalxrSlfPUAcw4pNFS1EJyGY3hilR5tQWowsIleHrCeyitJcJhh
w6F0U7hgZjhqm5oPv4L0+ytu30sieOSOPuvtuBNRBmtii7F9/j3dZuvbxnIb9qCd
f6QZgXNy1Fo0Fx06x/ymdXkB/dLCe379yO8Y6Xj1ngPtmVYPvINR5uIpw4DqGXAG
vL5Q7/P5vL/tZi6FKS4LfDgjEyKWPACigVw1jAw7jMeb/0HkvMzX5ELPRMXmCrSf
XqolmDPMuI4KFX7ydPRmWYykL9jlm5C6sWgIXR2jhiB5ATjCNOPl3FFrVrd3cZ7b
0qsDfEcLBd7NgoSyDbBRRafmKUGiyQWVxX5oSDOciSGdxAJaMefaeAokDVrtmEsy
r2w7ex7W+WfFau9BRozzEjFEkOYXTLo2Sny1plCic9MFzgcGJek46GiBep1yxFnt
Im8dpih05tRevhDKNMN//sF+k/XnTxbDZbdJqnINN3+EqL0g8yDYASgPi+VcwqKG
2DrwY9acAqxIqepCAxmJ89B25u0sg/YvPQYV+XsBlyeI7KfoCLuj8hzQOa5JrHL3
kLp0O06ZO7UUGoKHccvUaCZC2RKTKUEsVFJUnX/lLuzEeloQqGRgo2J0CuZe8JPB
DjcGxNgCyllGw0zoj68HNpCwMrSD8Y31O2ZuljdVOgiaEeAQXgS9BGd6Tcy7OQJ3
UTiYuN/5TCjmre855iqZYibCQ1OETyaOTNwkvLMx1Nd0FesobPR/RolEb31zfDIU
2vG6UIBjfXUydZmWIdSFo+vtCHk0rCLSB4UcOTOg0q1IEFiyAaqDBXcX14D72h8q
joDq5NIMzbNvUTi2voz4K9t8lt+dyWTNl8IEEf8qgvcGDclca2+HjvlazQeaXXBh
SqbUitEyejp2NoIFef0pxRGaUFGh4fKPaQQJd46Waz6qmIdzGiqtKz+wN4055Q9z
rJQ3F8WhZXOrRwt60qWqVU2W9R6qp65EboFEVIiQTQrfozOdJhCqltRydqD2OVlv
vNoZstbkkzoDJALzBwrBwHLLOvmkQG/zZO75ln/KkiFtUKf72FKAEICLrJmz0c7A
qiouu+ME3apk3gVOCJIySUsfyaGzGS8oTjI/O/k/+LSr3VpQRTu/Vab2uMPeoE5b
9ioan+RQ403raTTe3LqcUlzyvQtuxq6F9QtOSJMYOGaPQuUmOdvoa0MPfY1/GlVr
kgsPtVX+BuKpzVscdg29d/nHb8qjPvSczq2/zmhIDw7JPwFKrMY6Z8Bi6UaqKBel
iSGmYkz+ld0RuZEnOzCTyk+FmrRPoQVy38iF01GA4UyIMTwV75fDHJvSdqTKOkNs
OkfMHHKHtLSmIZ4jDYhzs1zJ54F3WV0NBSthv6yVLWBDEBRAGdSuf6JwdxqlvZQP
0P4o0eEgWv2YwGt6gEIm6ebmcAC5zcYvvLAHZLQ9vHuI72YwkQuHPmgdr30RDyJh
VLeudFu1Xi/dfOZs/m/yrFFEhK8X2N1C2lCopM1jjuoOzORuJtjw2lMlW6MJLCIq
Mz2CPU+mDWEiBPIdAo1/n83giRnRQp+0P6Z1fTH9igO0w0dhx/cA2WbS5mhpG+IN
mXGrZ1GLCsxLF5j12AsLAxJtm+4aPjtKIrmzSZNcbuD1uYFetG1RFXLeq8vdZffr
5lDN8QGZORqHeT9k1Zbd1LaAmFZAa7jFYegOrwkLkCrrQzoxn/C/NoGHnv07mbRH
2CuSFjlk9N0nDO9YCeLtRhRfIlIdCA/m9fVI9G2eUUjE2Fp7fX7lFvmw3DExm3eN
hwlQD5edh/tYOJo6QlA4wLkzvgF8KkJgzp/3DeTvgUfttmA5QOCDQqKKofgL8Lqv
n1N1oO/tnWIoxQA5vUEXs91ooQ1Bc6ot7lWpUXUJ9WXFf74RCVkoHXIMapPpwW+n
fDIu1KpIm7jUttFU1QiZIWhzWlG6IL3Tv7UnRrhvlc+X6haOmlf/E5ysmUNLBsc5
ziFE8BAMX6fouJAHHSFFYIBdpFmkHXFKHnR/s48jI00rShXa9Ybwd5QyCNt+aCOh
rrmv1GItltEQ3f5/O/iLOIoNJ2fjWEBDKoFk0cOgoHFEFX9y6qaOC+ZA8i55ZfyA
nYLc5RG0dvLv38znofVlTDdK89Rh36UDGfIgpT+Z+JZ+SKUAGVsPlQockq2VckRW
1PqhVLmPane0JrRHFtbpjjVsSsYI/YjSoPdsNAZx2eeI4qgX5nn7n89Y5pty/FBa
T/V0Wj4zfxHzNoDlSu69nUGNPEbfzhh40bgWZCukqQxld48sBtCUkuT41+KA/vEK
HHqQYfSDVjSLXbXaSwFvLTPNk9IYvYLCF3QTsIo8GiQOnh7Iv+79kxfJZgMUCs+T
f2cI05wNY/WF1hjfHAGR5+4wMow+ZrmbX7HMRk6+gR8nSrenequn7/pntqnn+x5Z
zxZ6sRK0DQcTP+KPScmSaiZCQTCP2BCWKxj/qfJN+je3cTl6S6sw7p5ZgInaAGGo
lBfSORCcPGzKXRBFHdW0yOZt9BDAdhtaZfI2Kh73Z0YNx5dDC9lXmNclRgNZzKr4
cCoBPvadREPS75T5nqRpIKYqzIeFvENgRRm34T/EuqiY0yBkTn4Zfd54ig0PA0mx
tWxV0Al4xbCnDb3kDr5scuvN6X7KK249pdyPdv4waU4tLirF+3VFxBYN8j1P61+X
nTmV8KA+R6PVtujjmwuEv0guoiIAtgSC++T6Yxs8Qn968viZikg/sZW3fNGNPvBQ
gNL9foZ30d6r8ABMbz5SIjeqtS/WlCo36iG8bQUd7RVDUbVZaKFz5egydVWkwool
SunB0Bri0GJfmR/aibm98HIxw3AeobYtXR0lOe6RRx24g0dgOS/EQm8YToVTjpIx
Advd/YoolxNWHiMxxF7O2g71ajwT85IXlv9x3rAoF0+0Qnj/LNYtk0M06v/AejlF
Kz8xIgYc8hSZDmFkLrdHLorlPYkWYPnPztltbp71Ozd1ubbutyndlud6yj407cL+
OzhNyPFGp1UWQqcpsxldXGvkiKmfP1lynlWox6nLPbU9tjioqIMNAAbSrwVQDkG0
KOiqzx25Q5al5lkJ147Br+F/Wgwn3fP1fEj4Bdtu11VZ0Qy2y1RqKqqUAMF/FSUk
dDx262Qf5Cd5+2sGf+Geg9TFdhPbsb29fQtdTpixHtt21zvoppgC/qI/O6cOvVyh
BOaiQMR/Nyt/yPPqKf1hwFflAYlWMV22Z3V7AMPAwI8ZQihcELsbCc7/JWbhA1uZ
Ni43G3HnkthZ/PzNVSwAnzEbX3IEp4zWoqrO1YvfDtC9ef7+7AGT0l9A7pS3SxtC
SaTfB71rnOBVooLyDY+0ieH4ef8x0Huu8rLfDNPxgdUq2KGwr4FvpOOzTq02pSc9
vVMeADJKezzh8TrlG+n/GLu5lBFwwxNVIsjJCbH/e5U8ZPdKq1aNSZ05dcmHAWhP
XrH6+pJcPiqoK6SOF2T1+trxQ8Oc4mKM1qzBbBkM5wEe11TdXjRQo6VccWSb0ODy
o0jxJVVg6zLaWVMuyqHYtWg2JxGo/Vsn/EaN/t5pmYKv2UGcs957KYZpZiZVWiy+
XHWSQpZTWQ/INXWxd6ZW5L4P2CqS8fBYiqp5M7UWKOmi3L7OrfqNHfLmAeBFYKkp
ygtegomskGntIdGmn6ZpXQeOOsMpSFgRZUMX9QFr1ZW2SJpHgZE52xrIegXK0bx7
a162dshqkiTwdYuZ2Te6UVnUgOcFrf0/fX9tyjMyHeMFgwDWkx39IfvKMwbZjKP4
t8EA9wYvdfKi1ECWaLCU9sOYgouqQsZB8PjyydGm7O106sJAT3/zdlEvzFYa+l7E
mDZ35+OMW2ak+/QhGz/8Y1qt+O7CIXBrlwABSNItRCuzBqlUbmZwgfRkLt1tz68T
wEyXusEg5OdgFbJP+9Cvc+HXzCeIQg4CDGWoUnFGwbZiEJVEyc4j6O54bGNqt/cy
gKTRB/isKjE4qqe59TyJb+yQA6NSuP7ODCrI+2uxhwsepCQEtSjR/QEVAee4hovJ
YSpzjeDvGQzHRFNQw4HVMIdrMT0+IMIMAqVG4uOCwLjvMgp2o9L7M4lF/NILUIhS
Cnxq4LPL9TNKloWUDQPeA7tn5vzyS3CYxIlC62r/n+7fT9FyxWcbRA7V7mRitp8d
CWTX33KltVtzSqHtWh7OqVw2+lQaKGiL42PxaI5SE9v+7dOwOFPZcCA4oR8/JjkL
TOnvS9vkTLPZd2ZFK7rWZ49eR9NO2VT+xwD8RxCNsHDENIydZIjy/c2xVSnBgbwA
rd2j71FWIil/2Q6ezt2DHvPnQ67keMUrhRodQGkKVtOzGl9TS8yIUFvCtAUh+dKO
o5iJvMppK2+GFIA2hqNsa1Vr+mTDTgEu39KUusUaL6IUV1ju8TG+bpiMrWYlCWSi
cM2qyUnIDewYuhqlKrBYcx3dNCmnZXUGeaeqBFfQtFFWBuoCCPNcBr+ie/T3fzZF
TDtOvxtQPrlqE+spE4MfT+0pl7XWAy+7X6P9+7DJiJ3STkD+6NzcYHiUsbnJ4ozZ
4f8IbzTcXWgRyHTp+RwPZrqbEu1nWYG/DUCD9CCla7PXzXUPIy2EUbe/sgiILz7g
bM6qeizXeJRbFn2wtHFffuK8aVHqhGE6v9AJNsmARdGD8rus13sNmOPorRz45P8K
ZJp8b+LQaECfXfZWMAY1USQARKV8RLxcIkgskKYR9Jz9rRXR4wzK9q7Xz4hKncyp
mCrqMzPVRJXKAJwwkeF0fpnC4yGUAXe1TSCIk/Qlb9p9BvNd2V92PoRCK3YlckkJ
jyJRAX65o163h95ryuqvqi/2nh/TwlNEXreVyZiOERUTV6oBrjMeIRaPpFNlfxe3
oOjn0dLpd8SJ6wD/+yCuZISKaaTwtW8RmZ9V8mEqZRGeXN/j64jVGupgExwKXzQc
MAhgGUgTpGU6BVgkPz27Z2GNe2IdK8IblmQ4u2xjpQ9zEZG8NIRy3KL5Rc3yfNjq
TFUEkE5epMJvNxyrAXALjv2vClja3HvyOguEzgvDDY9xYNpLq9nwAqGObo16rY6W
fiqAIUlRrZwk6TCo/AmJ2D5zd02ksjW8sgFkUSYWQKbJD3m90vTFrtUTuvmPKkeY
b5mqFtAxot4pgbXzsuvGuww3N0MXSD0DW5gd7+1h+OD0cM9rr371uzJPTQtMQ5nE
uN19snVBcMjRBa7pzRa9SXXNnMsVGDPEVerGLM/OWYfZI7WHv4zo9gSpsNC7RInT
CvZbLYSHV7VnTvBRTqX7segYm28tArQcKbxN28C8m3sSkt76qXuC3fauRx84wGLk
gTaSo12CvjySSNv8FcqPucbMjo0Nvs8IfXvrSy0ckW9HaFUOU6OrHQqJkWuuCRgh
olC7Ux2L9jQflrJR18Pm9B0+ftNVUYtbLmAzQzza29t/Fo65ggskOkj5+aU+Gf6P
hUG3zqMZASQgl0pk6U6J7X7W0llO7sdjg8HEYG60vi9S1Nfdc5UcGVIyQwNJMH4a
zOp5YC8PcUUv/hTLejy13aHHon39c2W05E8N7M1wbaVRNoBtq18CuD6Q+ZbXzphb
OyaKeFMwnmYpM7/VRIhdsnp2qlxcvL/P3SD7i9ooesY3NbRPqwuGVU9Vv5MQnEeS
B7TxIblG62qgbpLMBdH/ApYe0/KDlxjrx9aVaq2rk2UoNVI5y7vYBJXxETMrm8Vc
MUXnvAjKvjC0fKjdlPyg+swK/bX2RfMA4n1vXYua0gb4sna0zoTIkh0WQqaTWbyz
GiaS9Vw3D/nPurm1VFrxh10GKtRKw8cEFH46pswopgshkdeEjIR3V4Bi46nomJEX
jgiI4JdHHl5MMcYTCW9ZJU1nR/GzrBw4zQXCPQdBdjEnp/zrrgSMrDf+rOr7hRcY
aHW0OeZ5Nl3LTTo2vgJu13sBod1gB8vXY5FkZJXDsCvCtJSaNgQNkZQ+wYVin8Cj
Id2kmowkkqIhrEtMuBRq0nu9Q1eoYbLOhtMb9XnqEy4diFFQfrHwR2qt93fuL90O
PWM6GOcSAsnzM2EogPTUlhs0sHwVnT4pJqm85u4msJMVa7csiJYEbDt4Ml1QU/0U
0VLujZaAEx/bE1Zq2Ycf2GYfbfmulfCoxSqzRuGykvmRieJzvQuHx9CKHFm4rDGQ
sQ5C7RBh3JGHwzHQ0Q8OQ5JyAO9zscOj1R/mCJytKCPkJ5qcWkNFI7Pt3UbiunuD
0AXH5cdxh5/Y/GXkLdZJCoWkmuCi/30pIFpzdk201dV1NJhfaMXFjJ/aSyaATNdk
J26k949bvIIq/TpsSFWdnILPJd6bN/BCldzK2JzHtDHsLiMD1SevdIPl20n95UOu
tGH4zEe+oJjHFXYAQ1RDiIlxx/8XUGaagFT6s3lQVkhnY/tT3Q17PgxJuMyDqadj
E/zDqORi+KNJpJm4iFpAaoh1WT9qOjDgFZ+flHMn8BnlOEhbuWsDYCFdhMOhRmdk
PGZftjjFdv4Xrh6nhGnX74SZ0lQfCMltOJZ3ZehgSuUXIg6go+e1hNWxmPHqMLf5
SwKG/g+8l5obI0AmcBEYUjAhBY7yvdpEUl8EcJ3hy5+Jf2i/6OegizOl3bZJQ7gz
ggLkLN3eGfbZumHnZbyqt+tl8PjMnsZi0bDnCKdwynPJ04XGPBLkoTlxHUUFAtvt
Rrhan+9+hMdLY3GAnsSo3+rKP2oIbVfg5xj9mUy19lcINruON6ep/EUMqj4QbGAm
jndBsN/zruL7fPdw+kI0x8Gt3QtjaQPpiP/l4nXUpJfFwruyx3TCBFbzi0I5WQ8/
VIKQa4H2o2FvwgOLXPymCSpNSJoYvEboK40j037+et7ixz+daZl5MmOGdEsvAOJC
uOjN+sac1jJgs60ELEmn/wARQkwWuO5Whxb82wGqRkZQtmUgVJC3euRn/EQrCByC
+BGW3eetM+mcVIKMpKgDoafh9Gq7mnw9FZQBts0LF6rAGHIqCNsJJKp9OkikKOc2
lbxiFWqGL0VVTEiiWWJizfP9oG7UWXg7OUbSTG72q9oKmpCVBWHpK0ZVPUvdCc3s
9EHnGCXAHHj25FG4kF+cfSQ+nVbfiNZobkE5bI9IlarAhdVuDOCECitBCbk4eZgo
aSNcbe96MYpB4xUx4cDYan3AwHN62X7pcsyqePb19XfS3sBktXbjeaIye+M7DTIV
yKBWFKu8y5JEHAKb/jTPyKM0xaFUg5KYuosmE97nx3RqWenrPlPb/T0vaHvLjcsF
tXqVYIKJLf9Cfj+7zTBuKTduCGa/cYc2/00QcpQppjfUCrSytISwFZbhWXQTNHFQ
7ndH/gxUp208YT36yL0cauGSX6+7Ny3NTpu3YjwmknLE/oHakxPYJ89c28/f8zHL
PzIOCrW2CqPqJ/Rtxq6O24IjZQemMgbDCtN7m8krnfp90yZCANJMXXxlkrbwBr8K
xvWaXNYDnrKZcmmHniX3wG1jjHwqmDMw4JGR+HmnN2hBZzFGUCj5c/nkiN+yJLlB
faVoW1rbaIGBz4VaZT6X8WqfrtsqV+7xBbuToBnqFkmZIv+aLUkvymE4771IuqJi
CmsCc+voCUBbfHzmVjSnNiCQqhiiD9nLfzQLnT31nXDJCBKex5DRzAH9p04UmohA
L6LKl7t716rzNBoIlterfJYUlWiqD39M9qmC9hUurh+T4MLUnW684dmd2WWhhElz
vRRz0TinOYDQEIuv+rkTk6PJHv6DEN3UxsRwKTAurXmXwRYH/WNTwCL/vU4GzNMS
VPkBOINnMEn8DdVTSJcB7Mk7W42Pq1usdIjluZnYukYRpxh1w8oZeDegswY0VT5F
C99uqhYTZYOhkHzz3CYeABsm8q08vpezjhre9mEDWKF5TOKY/f4nk5fJBck8k9Ij
/J+bgL9ceaPff4M2DtFWhGkzBaZUM5r/DV9GjL57b47AmlNEw85ciLPw2JnhhtfV
vGnML/E37AGL3ZdzKB7yrlC/CXCojz3zXVvl0anDwwzgsOofxeg8iplsRtYLQ8vF
FTuCQgm183xI4j6vk5NQ/hGInwwxFnSqi/pUMc7rPkAfb88jXD3PRYUgkuVo9AJ5
K1Y+B9UT52OUCjcjkx47odZcju71WZdSmdB/1/nBfqMwa2OFozxGVAWHNAM66Uig
XMzdER1hdUSlqfceureeZl5IG97JNTL4tFO3KNzwaHLZYzQPYPTBR4tmJ98VXuwa
zoMFnTbLn6+yK/8g5bbdyBoKTNz3ttbmlo+YWfApdkhs5WOmfMcVbqBz/EPXDV0O
lbfbG3/BRSlY2b3qz+JKNDKQIkDXooemi47sRM/a6vq+PMx6B7VdmK6Bru1ONTz3
uzpBIWXMubc7uHcrMA/TgmVYeJJ02Ddo1TnTUSDhvmqxFBOzBhMabCtFBM5XivzI
tSagJ/yJk3nxfemGeQkRfrmByX8Xd9XJNqhnJ/NE2NQz11NNIcRhOSIfq5d2LVwX
4mTb0tmDJhub453CJBNu2qiyq2wq9xQUcO8dL6JMrCVoYnxFUae0YFmGL9Sd1YgZ
xXQBM4vx2DORr0HCpUK2opD5CAhwPX6Qmev2xglBZl+zg1W0bZaBBv+FRLwb6hxw
be0UM6OSLvqFbQf93FWVRq05Hd+aNjhN/hRAQ+rPCz55vi7nAQleYFyFs1Hk7jtL
lkh2rsbfu74+9K8ZY/s89c/uRMvwb1mBfWs2AaU6WyHiJ5PG7n1lMrHzTUSxFrkm
BKXQxLSt/V0f0TnEm9JSKalwP3hdaKbyzI4i3vLX1p+O5b78x1tkb7DwPC3RxKCc
TpAyyco7j61G1hwThrdBvunJBL0VRmmwcVMFiU3nC0ec6Qxb7+TY3Lnw00m5T44h
KMeKj64e+yT8uOS1Iwyi0parF6HwFq41X19P6DLox6u0thKpqjcLzLGSG4lJRDGv
oBkwiXOycUQsuacs2fS6ZOZ2mAdN8kTUikpWhqlG8ERJLkqH1EiOHDyBzv6oKMxp
08duUO4RtIDMiNY8JyIXtjFBDb04Z/h25ItiXxr43gBAYAUAZUgQ25L1s4iVeeDZ
9qblm8sC0rqI+bptW45cUhHWF15Q2wyePrwTo4/qV79fcMBp0bHNyH5LINxFpdCI
DNh0MB66yNqbvtD7nrqGaabydhj+k+qjPjgUn5sLYPSOFpxdQQpTI3Y81NL0g6Kw
EJ+eyoR9p92/3gYkoONgln33JmKuXo6jpgQ3pWIq0tsB/yjrlxhYgePb01UsCusg
Lxfdksl8JKbviEXmSFdcqL6Nqoj813oaJptbcod/cgBoy4enzIbKiRiucX0lEWdN
uQoVvHKXBSTe16pUn5ylNF/xxMVJOczcyBrlB57iIZtc3WY887wjPY4MdJjjVUAK
qWYleqhQwYr9nw2QpS9TNcMquRIVuuaofstDAgk57VtL2JfwjAWmeyVVjvOyUOic
5UHfOlKxJgyCcvhyZdulM8t69M7o7KLJTOMxozzDHITOliOeVQ2ivdJm0+xHMGB7
/mgBVII30X7P5IB/PRkH7Z4TFxt4UeZvjvLZ+cocBbwXPM6T4nadC09asjwew4vu
9R46sPu7MSU2rriVkc8IsYRXVgXtEKyqJFp6fQuj0EnCqJ5N4NvIdH88e1fuCGYU
g5rbx/ymklhybgAOZkntESVD1ZD2rhHz3hf+gZXvMX366hHG6JqLa4An/vmNuCwf
FY/ZQEUTWPC/qotSloNhStDXmx6leeUDCQ581uKVPiMtkodmr5pSo2BdOYk9HDyO
IirO31Fl5+W0XZVlrxD4wEXphtq1MdeU4vGDTEeAZz6+dOS1eLscRHKYGBDRTx2L
k1Jd6mkVqBS/yT/zBIPlG7pF9WSlyjZ5wQhGZRtCxLTl1xbA/Q7Jup9In5fGhy4/
uHG1LvIshB9nj+iti1QV1uwAXeMnOXXIRFfS/StsljqptmIjKH2OhxJFAyyZ253+
uaX1OILianfBs8yhRhCGG9ip84EFfEN+Syvzx9hY0ZqMXmzzTt3YBNBmAi4TZiFO
9LnqP2NgYyZhzwpKHUzS51f/qbCU1YUz3hNyPcUaQ+6rKoX6qlZo1Gat549ba/MQ
IidjL/aZFrQzKWJ8AaKzfpytqTIBYvCp0Asbl377jS6aL7FJJK2+JPKSJusIzmST
tsD5i3dQm88+zz70cdvnpHoRNDkjq5fcPFcW0I1haPRDevSnPcyyMYoQhmuSTzEi
wX5PnUS4k5/laGYQoPivQnYnplVnYEHk2HHaIioYhb/k6dZaKuQ/QrZqLxCCeYFy
+/7PsrOuZ6B1XYbeYGvZu5QK6VCmnLkTHUktblfEgiOU+UbehQ/JFwaOSg89QAA9
JLB8YFzySsCBJNIcBfQm0PgPXmsKyTrjPf1jK7l3W19N7haL61uYa1lFxbQc+r17
B/bJ2R7aoVJQjQLuvBvOxmGCUQNGgFWnLztU5f8nAUykk5hnLheKvK9342NXQyzI
k7ZT8eL0TZhWYBr9ssiNQWNnQfeRsjao/bHN0YIhtZQBvj2R740ly2gTjgqTVJ5g
rJVbPqoTZdxV1Gdg5pwrrGNYvLPHq1KiLW1IOqh21xNHw4atKhsVEUBGIeDjzcI2
NRe+e2T8xeKo0MAEwUHTES8KpDjeRPfbii0PalNQRSeMEfbshEwAxsj4m+AGj1qZ
/PL5FcNYgdJf7z9ySxrgzAyAKFCtHkC+LZaL3x5qyn44w7bDvmppbvJBWa6akurm
q3ZH3yEEmRESHKKttu0hbu3ka1n55UWb9nLQmPC1IjwiF4Wt/TTRnU+15jL6SKxx
86oJf4697CRbOgWhVTYecr+32WvchHc5106M/Brqnx3LzMYdTEKiRLwc7jT8Wafc
iEelISUCFxzTO5FNjo0pLFnGt5X+CURCnoEwBY00bOd9+BoyVEDZqDT/76LCEUE9
0dayz5s/7/QFSnyewx61aXGF3EH2FMT6rSkYprP174Qb49x8D5uYCfYY0TbelIaP
4Fv6C8UeJoKgvHKf0fnhZuTVG95/m8oR0bhDBM+7DNZj/2BQFj6hAvCkhkRtQLLS
Dz5emDHwBsJnLUXATxkcMb1JP5+FCx1xwjixwjelpAOUgMtJsX9UUGknjw/bWKrm
f4dP3nJ3yB6SdSdRCkc2kSsCFArVbvcu3qxA+B/mm4T7UqJjeze8tr5vOtYGS+Rg
Ma1gMyJyaf+RvQok/IBjt0bAoSBPgRGsFXUodZAJ734ITAn/vNbFtJAUvTa+LPId
y4fL+J6cz0KrJWMX+Hscv4qGpiJQhTtvA0KQd1PDfW7THV5mqsDOTqZMXPHLd7z8
sqh11hWTpqd5dFCKkO+i2PlDYvE35kyutD/ddm1rzfy4nHF6KAbmwG8thU8uiOrv
j75xQnFcUIFYuYVjS+FE9Lyy0e+UltJOGTcoybo5ftSWIkXxiArTJbDdNfK7PZjk
zaDb7s2QxP3Rrwqni7DSqmjzRB/bP1N4pCzZlvaFvwvZxHUFZ6jzyrozaIzhVwaW
zpMasIAWoK/lc/srJmHqJsgu1GeID2iPRbAzOieuvtakRpJzuU9Tazu1fhE7GE0d
BHPkr5r2smWcF4hn5FP9cAcTTGWzQEN0c3xWrHZbfKOTCNI8OhR008qzNIHSBNOg
kkTmpCY9MvP4/GRnI8W0UmgxonfSKLamNyTSv/MP+R57jUoWrdzzn5hW8H7FHG3a
TIITOkgLXPI1UdXWGHlkKQTe2z4sLQ1tddH6O7guPv61OtTZ2IEiM5Nwni53wE2V
HFmwhYajAnHNVwKPbbORmalcklixufogaFs+febHHkW+9T81ckA1J1RHZje7t3RL
6rOydkwWmXwQ366QO90tS81ji6yFXRaOEibSofqyonoNB36lPuok+FUpzgLtRzRT
CLSKkpaUZIARV/Poi6y916NErYF+wTtPwQbNWaN9fXXykRIheh8a6lnyUom0VQHU
+R8oOyXnQya3QqMlpBzgw/AtriqC4FdpuNQ2VtKjZMx99nJjWsAhtOlmDrfxrklV
bB8sf76KfRt+sWmfD/kzUZcoSLctfTH0pi9nuHnYBiS60KICzVjzbbhKNXo6/zkD
hKDR97/vUKt3TT/dI41hMKtSb5/Os9lVr92+HMAKrkbbOIpRCm1cNt4I06A9rOcy
Qzn1crpbh3i35tQN+8WjpLo/t4X1OhTnoKMDR2AFcBB3Sk9VBygliAbPierKpQsP
qx+YN+k3rgERYc1U7NC8tBUeZe4T7SndztwEebBerd9R3AL9kIz2EV0kl5mOQ4De
kOLdg7nQq6W4z1hb4WNGxtQR6ULeOQp+rwJbWGPT16LGaOh5uTBP74ZXA48pJYRr
8xgxeb7N02y/Z8OnS4wrVZBmkinwaKj7yBbnbovnnvdSoHHcVBAjtM/qpz+5wqm7
bbG9I2tQ9vDklc3XT1FdM6qDhNDj+rlVFXNNtzbiXK5hCvhKQR+2H9ebXiicsX9a
FG0DTme4C/WWLOKFCkJUNmsoDNcyyAzs4+0BN2183AXSKSGgsdTYs1ooVAVrdFVx
WsZ53cz5gTzsaWJlmLR4zsnFZVG1i2dnyl03+hft3VqNFu5XzDfk9ZB09LRFiJ0V
1lozlJteN4aowr/vTkXrX0405XlnJaFCQ+vtfMxfmzjB291iL7GdubpbAAec/5Wd
nXr4G7EUmfKjYU+1NnAbsYSwra2mdQcC6tOA7391mj1j6dgUwZEL9O/LM/Ttj7vP
NMtinT+xUxIvrCWKGFnsKPDMZu1jF32rIC4mm1uZQMKYRRHILe66D3spfrenBOrj
iFSIkdjxGtQPfIB0hpWrQA29JvGK4aU3gYBrqOYo2pCIM7rVSKT7//NMa9Cr/KeI
LqQQO4y3LOgqHysY1x5RtJpg7ESJRKqXOoAyOU1ms6z2RG0UY8LAeXBZS3ApXrw9
uXGyUeFGqKxums7G00cnDpCO0+k2byQ1mQLrOk7ItfWoNGo3EFLTFODYP/A9B0GY
feQL5+kYv5ofogE2h1kECvG3GNB2/c4Anb6GcduH7I1sbeSjoiL2M0TTRwuIHqna
rTzs5zS9nKFHkPild/A5nip8BKgJpsoHCX26LqYj5muimjlfoHAm4BNu8+dTR9vR
jL5iTr8j/qo8pnq9LWFG4+mJzFaIq+85wbBr73nitQZCemWY/KocsdBw/PBITvSf
21hWlnu+c65xZ11jTMX9im+NBa8WkvRWhyKzmIAiFIESraIUR/fMuKckMGS489/D
/5Omtw5v/iywHX7L/NCbblGd5WIa5hUgOxbcRa0bRCOtSKd4u5s8s/lOkY1x5TWk
Y58hyYlhO0SEod+Xdl7uU/e9wO2542+nY4Sp8jwLA8xNKPUWangbwxCheARKyDum
AAhNMOCIFz25IKGy7Wb8XGCL3IvtWkYoU1obpE5FaQDFrmYOEOrmAo5zbMKCqXbt
pkKZEOr1oPOd7D56caiXs8TqOgvmYj3ampjQ0wa2aT7aNSyeaO7EZ3ojHot7pmk2
k+D07s3MO6k21fZLkOBJ6RZcLupzUfjnyzlir0gZFvcBx/dFeB0SwSdOZloyousN
xmFQvoC0RcsJ2MOYuShUobxEGRQtkHgplJzUcukjqTXGn4Yqm/Qad0Y4yYMB0YC2
0qMOwMR2VqsmdyEZMeO/Q6NTJL0hkyIB2mU52fUKBoK/tY038oQlFTqUyn7pyh0X
RCVk+0XMFxKMad+pJ4ayPP59zIq3kyfF7o4ba+CJlN1GovpqfiGbaBuyjnVB8gRE
0e1b42WzVwUUgn7AsweI/1NDpQb+bsVVvreuPO+Olpjyg0MjoieNLcSkwn3XTPW7
ltnwaIk1G44Wx3/zqDacSqHWJ/2IoXdbMdk70HG9/Lleqbzh5XYn1W4WuYrQn2PT
jmyx+gf/w0W9njlc6JScJywjgUxQiZVVRD5YMR3i1Xo1lU1wjxy8M+mUAfPcLDB2
9syN+vNerhONCTC0yfulUiM3ogqEwnCmrkcQVUvl5ECuGtQTTC6PZv9xn7IYtk8d
E6yi0YWjR/2+Wlq0TAjRxyWl4tfm8LRh2XAFigogXOR98ChWHYPDflSsD4OySfRC
93/RX9uTwApg+o8+fc+rz+CIbXrCMlf9+OpZjYsYBuoe06VydJIkSrtctHpKk/Yf
oqt7LC2otx3s0lg5EwStKoQuribL38Ny3ic36xytoFG4cVn1TNAqkG772v6Mh9O/
JLQ+Hth61mcF1snk2fQ8J/MlW8DsL+9N6bgxEe6g5ZpGkbM3+C/LPe+cmt4+K4Ib
ZCW4XSJK1kUJ1qBhLUDjbi2s9sW6KLomymdeXVwhFwTsKdikFcwb3DkLFqLQjjHS
m1qpmrRE6ZGItHJi4+XiElCSGB0pyxKc7EduCPTBf7+WCShkHQ3HKWtG1MxTlOBz
E2B9XKQKqp56SOYQNxNSN5TTvXmXUkDdxvgoQwJD7MiQhpM5MJebTUq5wxSJGp+N
RAG5c41sV53mXza//ER46bE+50akoH+0zNsp5tEJsj1YkQthqoGcr8T8VD1OFhzx
Xu4xTijFYL+dsDMxPDDsthSmRk7Dqz9esYE5MLc5Ow0sG+vRXYWQfplv0tivb9+S
nWY9CdV1DD2u0Xz2wGIOjI2C1mh1fcmdl78+A2M6ka1SBc9SgoaqCfGcLem2aoLi
vf88PYJYON/7q/g/i6ES3Kwlmka19jrJweYFxYoOSPaC16ZqAnM6OaCSgxhLpDGT
YIjjVlWfpN8nUKGuPE/bT8MS/NFbB+KREB33pm4PkMrAPWWzZycwq8B1Jgojlepm
x6w0vy1EZMSzckWxAlKNrd99zoopoMZ1qdsXfwn4FX/LWUmZXIZOFKeCOMiuBcAF
5Xkov88ceIWfbct3d9cExA4d6Embxxzr2HNSmruznQWAodPYjIXVZZbWJ5Avcss3
Q7/9qSmk6nq0WGslfDYi5ALcMapPDVxwRTJbYZjOTUYWljv6VV3SpLaGJ9m25pbd
w+6a1BkHPx6WOZ6VuUiKvHJ0hXlF7RyssPdJ6fvrw0oEhGQWkF78cQRefdUYxKEr
ipddLob1AIZaVQf0IQ8+uUjWy6GnFFvWywKh8J34TTZzp+NzUJMsfQoFNz0zrT0e
xpNBbaC89YNdH2ZK6G7tJD9EYPZT1Z1wQ88HVjr2Q5zMbmD6TboCy35T28azutE3
Gzu7TUtMLfOk9vgcUYG8D3QijQSB+jHqa+WBqPjJN326Z7T218HtLUF5DxTm+Xnw
2ZiMWl1I2BEmmh2q6OSkgYM3utPOEPqhLzUY0VLLk3wE7SK7fZQNRFAvtlSq7W86
zQjJPPrfhnM8YfSNt1GpF0CuoLVe/fL5LwQU6tzGz6tB+HpumKjXQckLa2GnC9ug
coc8s7nOjvF4xpvBw4czjE2W6P4IZroudfvACujUh6bN4yWmkOepfYp76WiQHWpD
3C8+m1k8K0OqxRZq4ikf9BJjacQgtNeewWWfsmAz9Ti12iKiKHUq6xk6U1jhQkNT
6fCfGNkvQxS5WuqoiZ3H260FaBn3uDmOW04onwPTZ4FN6anN32sUmpm0hvjeTfWf
h6Ch3VdKjS+dDgXm/9rHxCdps54vz8Iw5QFExPTlrjmsc/G3ynLFHerUMT36dYEo
69iowQA1B1IBaal3Js0GhyGaC0hqnVoTBpG8CWAtqoktCVz+DR5jnpwlPBa3ztdw
SIZ+PHtY2vggGsR1d5p+R4YwJP1AfowC/onYNMaSn2sx0ewpICkh4N3mfI+verFl
GtXErMzplPNPdff1+5kdfBUd/8qs9pY+0FTg+j1v4U3wlRIMoXMThXX6OKzF0vmO
NmvpuzZK4xdG97LL6EASebRRdh+rztHlp/EXpRx/tlEFXmsDNiq+C/JrGDtdKE83
5yzpxX5LDwkQd8TqaLThUq0m/qvJC8T78WzAVT+Ots6O48B10qMxuw7YIL1CirzG
ywWVhfenrdowctnJlOXs1YPoszhMmClZ0RI0vatoNzzOvA/1aDZva9sn4GTriKFY
Hl1iWUnJU+PA/hrDBhvsdka2zYJvtho6sl1ou74WP2T5SqCNW/Uu8dkRj54d/I7u
dees9gl+OGNAEss0rXy8iIEtjROSsq6eqtPS5nKMsla1a1XdGaqfv6Kpq5IuIE5v
ngnn70MXY/MnvgzhXhMeikjk3ijN1LFx3golcRbIccWwmfhod/dRlKx7AfSc6lAj
u0TCQ10GkFJa5cgWnxyd0RdUkuUqh8R23zURMAnXuYd3GgLItVyfrUFOtOkcCj9Z
no31aFma6V5bXGnNzUkLRrgOxeO0Oym5ehYOm1KFBclbJPyi7PHOIeZaONBQGm66
4OGTf4JcJE/ZaF5qi8vovrQT3bi12lpYIMHRbQkz+Nh8metxDAoc8wR+mkKYx8PH
fJZeLXzHtim9OJJApy65r/2aMCbVOQR6dEzY04D3OTF4hD0Rr2a5CzAjYRIgdyqb
djhcsSCKieRiC70inKWEtqeNA3tIqvJwsSyuSNxQfjwGEgfluY7lVJQzE2lFBcyX
1WzqFFOVVjuxI5vewnQXY8fHPqqstzdg2RT3pPPnDa+5NT6ENWlwb4wnRGrBIr+0
SaYraYC6ew4Z9gos690ZAh1hFiBlDWqoneyUUa8WF8LDxFfb8BrSSBNDQfFHN859
YlPDb35R3zzkbIY5/9yxUacXNGyXbxCyG9y7+RXiOxPtoZ0rP9Nh40GiOd/EMT+F
S4gkzoCe79pyN3JoggllBSfvCa5UN1O9ZEOMVugJbwvcK+pnOJRMxlveBqfRVbBF
L/GKur/qC8KUHve7Y0qkFEOyYre0pMhtZPGPkjgsp5B5Qy1WGCTBCnOmt06ttdx4
Lpcb8ZoPwRrX6GTc6dW5FxsJy6DH2OEQY0Xk3gqqSyriACDNsL72sgTMqLPka9cU
XNMUEU8ePwyh3fAbxfEr0Hok/guAx/Kv0tAMRi29lxrlNi1SJV+ikGdEJPmmwNCc
/43xXsHGx+GntWPkoxhRxdHlXoVcYeYgTyrhL2Wk8U+u+YDtVQTx+SEwr0abRs/r
vvWCB07uZ2efKVl542QNR68p3swpBB0Xida4ZOXLf72+BePUQgTbU0SSzQLVHnUz
0yAqudRuAvMKtTOAI/UT/xMABGisRJ98LUv+Ix66nzzn07Sh4YAwRHRyS+UXoRJ0
fcauhYJF3Ci4kf6+KpC7woeiXiwA3YHZu5XcBy2eS7Owz3FenP7mcVyV/KLgWauw
d801M7jKoGidlzMQ9zodfhCO2nl+kDKafWrqV8FvEJuiKQkj1fEzwPD3cEpAXPfX
Sz05pJLcDelyBPBsCYUErw5yOKjE+Klgv9O7vqylWqYDTmajePa2OH4CWcqbiB+Z
JvdtU5wceOXQXRCLPKrxZ5Y7y3C35YIA0poPGBVLabPoDbiH3Ow/BG6vZepKvwWE
fph5Z+rYDqTVj4xp1guj3fJJN9rms2b1sCtSrZ5XTSXLGGVmw6XrK0+8PmTwBXEM
siVIQ6Qz4VBoeKZHL8u5+dLTOp5yQqannx7tDgozt17nL38u77pfGVybngjl+hEO
ujsAlwOfhjhVvWTROTT65AMW0XzNKR4K7RU7LEP5nU2tiVoO6cbrWfesRflg+M36
b6yKxp4PxPUTZxZUgq6x7Kvalc+/F1qGB3ZAcL4UwwUjRVrTJ7O1Kk7z+0KCv+w8
xaPfqz15yAcEN3O6+rek6xvWfipTQ/uZggurUZ7D1qcQ+jYrXibXLi5Nlqg8hl4n
Knf7d9x5xM4Y1h7J7FNexsv1knNFyTI1Q09gWm17kHc2Oz+iXsN5JfN+L9Pp5p1R
/X56yg9DVT1VZs5C+NozkKQbyW9ROVz1WQN/IcvyyH6Q/ROfG0eQUXS35U3vmw4n
Hg9i14O2wXUmPXVqnS5Y49UPuF7TOCt0fsm8Qv1RmL6qMr1/HnO+kj//3PID/HS+
N2vcrLQ1xjnG9OqVSu4Es1yyjxsnS2MkYxzR29NQVWhuxH+9dEdvb9MvDkq9Y18Y
KdlIoSzIltZsUr7L5i66Rj2+Baqn+TRb56fQaVV7iytKmPBZ+lXsh3RbzZ0MC9B+
GLYpJT8XV3JyKQ+6j11SsaSw5PsSsER+m9kUXp6szb+ShbdOm9DyiyvHtLoAqgXg
E6s+gUaoINleoFAcZL6rbMjinzb1YKcwDBVB5yLaPbox1ZtkiSpaiU5/x0vWWfhq
sS5cmMn5tR8NYXvMDmXuZCdIIPAUs7dvrCs0FoEIb1njDE9TV/zbpYnwC/EGA6Ho
LRhb87eHcZHB6rMhiF25cDwCQO7oAqlI3QHEWqFvTWEDJiQF04vb9nAw9nOHcGIl
2e5yIYmRbByakdGvD+mrHXfooOHwxSe475gLw26MYCTcrSePNt7CbPL3WxTdFyKj
YtX9sfNMUkW51I04TtdXVp2B8kVcFohznMOjZjomEnh1YX5VNlXO2MV7dhiHn7Le
8a9mYEh/KXhAAOGxu19r/plO1LRJNObDco6zXoucekHI2BrFJWqGxEmYhv0crNAq
uEenjYSmLO629sonPPtxCSwCq2+CngoT58403IWwb37tApfEfP3VBs7cR+QPe1Kt
NUcFxNxsqwAiSBELuNMH2CZ2gSxlLg5201lNIF7anTabYUSrDUS6IxLDC+Smtj0u
HzSmPMB0+LUMGyyF4RNi/bvchIlF89v0y8CLArx1HlbtAym/o62hJBuDlL+t3aBQ
oj+7W7np2CjcaLxlZcBj/00MsQOTthS3IsHzEpj0lqF+hYPUQzHUxmg1gumj2Sxs
LSfZXC5IqjY5QhdVrSv9ZxkuN+3aWyYzC4gJTbFBd3hSwTOPiEFsVJdjUshGdF+B
E3sCsX0THJ1WbSOjva5iSYFmgsGY1RH0trkxKi34ZXh/9tRz1jNKgHpQmHZhynND
EFD/MsffYNse/JFxpC+oMfYtqnghU4lSyLR1EKNxrmSe7xbsKvlVxS+E+JGdFgrh
75cT/rE0y2DDY8PuhHktYCbx9R1OyRZsFqH4FNxdAz1Uj6t+lsOWUQU8r0mkKJp9
KOD5Uz2qHrZp3Px0eLJu34snd0zFHBDLGN02zjDZP+Mkti4ec1ypGwNWGpxp8agM
oAr1hZR3ZYBLh1ZzwOPobltTrWMtuJDg54SiPrKzlNDliSUpiuQufpV4KtSt9i+7
+M6+POpA+4qxPK59btPkhIUNT6weEgcpcwnGiMTAZLSYlj6RGAc+WLk9y8YPpUbn
/xNY8xbfa/kUFQgtmR7/J4QipkhCAKZrS5C+6TFIR8YhtyV6EBmCnVc2fTX2aZhz
sQaUV4N30np7Y5rDT8YlouZWtQxRhxdKKlX/3ACR0151SbP7OstFYSb6PPqcECYU
3hN+7dd3EGg7whNp++yYCwyq6SJ/DGfDHa91HN3FnovNQLJ9VKffWW/wJdTseADG
etK/5V1mz7jPqBaZEU9iKdN7eu3MRKWfj+bpE91mQA/Jgb0eaOAkl+M4wDem0xDU
SZOTDIuPJdMlIYki+VZGRu9NoWBdrRTdSF4hSN9mypjNGlAa0L401kJA4lNBU8XT
gB0kdKJdVXkpnhU0DvznzdzfV1wEXyCB5JDRyRVBx/4cBDRhfZ4Rsr8IHz6h7d48
GtXqzXJA6G/t9jrs7zjsD0yLtoVoXTr8RYgyjpl4m9GN4cFsrCQMoK5bd18OiXbw
59Ra4mLwHzixCzAgRmNa+n0YY9oTEwzo1lHlIrWyTQnCv/lhp+lFi2DVE/CaIJpL
TnjC1Xhy1p9Jmy8q1GzrhrNTVpx4vVKLR/jMYqRM8CLwqUYSbowyDA0eMhw6k16t
ysVVSZ+h6vx9QzeJ7AfGrgWkNjbErIfFuBBw0Z+IVzQn8lqUIeGvRJIkTA5giNak
nOds9oIx9uqI4LhcBhxx9uEG7+O/KY2T403MEx1Pyp2kigrKy3mVMdO/NwAgGkdS
ixzxgzs321dvtX0wEkI37+iCmL3EH5mFMTUjlhhV/Gd0wN+roesgBaTf938uedSw
TIBqhl609qYOeDWv1Vi612IUwsTKr7M7/0Z6dG22WkSVJeBftq8bQn6foKLCPva6
0GIetWQjJR1tKpYmNmMAZ2c0GEoGz5KMQz/c9MVoAdOxy9rQJPWH+3jUc8pX0fkH
aKLDoXYRMNqhqG5eYAkq3GZ7yPd0cfRvgXXxZa/h0+apW3YfVTC9ufznG9jIgXVv
4r4labvl8rXMKN7JwxlmtzwNfCmkL6qLQv8vwOskZaXowKIkUpTihVfb5OvLQn5Z
n8JGo1E0/trQhiY1ZeHGVZGQ5dOz9OVyU/GceyiM4CcIbG8ljsRb65PPnchP4opb
8JFLxi6xT9x+hXZg1E+awheogE6eFXkLTQWJv2D5LHZ7VW4Q+7ItvTimITVHvXb9
IGmBfv+E/c5sVb8MCJ4nCd1AOQrS6xKTZBkQFMe7bIFYcdrJSq02uVJPUuGKFt+7
5XmmIwOrDy3VnrMwkFbmJ7BuDnpOK22b8sy4haP+ayzbBwNhnLWSF0a0o8773JkK
/Pr0rdlBGFG+WR64Z6hODjcQ48+ctHII1AJFQHUCbpxZhSSy4RxVOPUAge37DkyU
MnEnNGh5asXlb4Q0pJ/uJh5NxW3sjef+BTX4lsQod0gHowpv9coDRWj47wBJpLkQ
H+NiNE0kaM5vwqMFIfxGvZwRoZzI2war6UM8qjAFVq3hRPKIpFTeWFSPQjev7w2X
UC+g4Ylc1qO9c/0Ipf9FYQmVtwpBM3xT8YoCQorpmLnzEheS4cr3wHzNC9gnMnOE
m7tmISgHVHLmTwjPPxAg8EoFoWAfTTn2fEXMJKliiU0o16IKTS2crlGm03P6tigf
bnE61oncBqoaumZZ5j2lqTwCPoNZUqbPB5AAT68DJ1axHsx+ddj1z9dmFkrvSog5
O1S/c2ly+cnDQF720vxtbd2bm2keouZDPA4aNQhYiOQytzWXRHGloSvPigZ4K1Hn
jw4wsbpn5LxblH/o4waNqMg6455aRvyAx8vlLhRIdL4VPl8lkVAJUbZ8ryhSecLQ
TKJPEXa45q8r6zd3jWZnWkAF1vMhi/2HnqSNQ9UmWUHrr6Rn7XVyuATzjkIm+nd7
Z//bGPilP/pcU61NIkowekpqf1YpoRVfUtVraUpUHKQ/JpBHYdKVXkzTa2+Feehv
iXnMjDKfHJunqDSc9vL5K3aeY7raO+2Los3wrE4vybkrX6mWu+caevYN73WorY6s
Mric7Q0D5EpuKNvJDPUAVlalpfdzKBoyLixjGO+yn0UDSE2+im5KD5iZBydcNDf+
T4JcCUIuVbSVULR0eNMnGLSmEx5HOUDGwg99bpd1jhkNyfAlH1cZVHKLpuB2EMjQ
yP6EJ2vTGAV6sjRLr4p1rxWapbrF1UWzWTUdYBCy9y4CgSDoTDSr12LR+Fa6nkQ+
CfwHlU6GpP0mo2REiSvh4X3c7wIntqSccQBRcdQWT+T7BhyYuCHyYpuNYUXhUhv9
nq4eQO0C/ga5wSWB+XQD0I27nvwpZjF8rkrJZ7Cf7Q7OzQPSmijQ5VPKPtd93ap9
eUkDpS+UQzlk0Q5RnTQnRkWDnoSHvlQXC0jc1kKYNwa/Cr9JelUz4G8yGS4aykc1
9cz4OSDmvTKsgotAe0MfP8lUAAzwbO4leybx+EQzX/ppZleVwPgQ2hzlwiWYInxy
hSWqgOl/AvnrRYvgfg3Rs5ar/6e6UhXoAYUuW/95N7CDtX/TqKsgIatgrkVc1ubt
4wo0XC3eD8tsacwa2NxxrhPSGWSkIb5/u2pZR8DUjx9j05Zq1PIP/3AUeB1O57CI
2N1B/NVdI06ZXIqB1Q1QkRoo1Sd/OKuhJo/IZA+1eYmshbMx1MCiYGBfg6WlXWF6
IC6E45zGc7rebhgqC3LBXAGnBAsHtXObSv7Xh0JI0HaJKS0OXl0DUIxRKjBHeV7T
G6RO4zcWBsMwzFQRJ+JhA6JE+LFQd8gGyDkNFjzRIW6RW7rxjM8e1I4doXVetnl8
Vk8bunbdxvKkgFk3+rL9WWvA2OuZv69VD1WxnaEz72VBPlW+WjEiHT9M/4UxZyQ1
AbO4E23FaQ3ao/sXNFaiE7Pk3MFFiOWm7WrF49cOatsgJoaVsVXWCwphw5Xpzthq
ms5SCwVmj2wl2XD/PtMHxaC6qOR0lPN+45SuYmHyw6XWmDR5kBV4XdyOnE6wSCB+
hUp8VsY2ow8l9eEL65ErZBT3h3GmQB2KAyjXXBG4hZCGKhRIP4LssSGkG0cm8mEI
62Do7q24Hilq5hoaHr8pzcGaacBnbelmLHh4gvJl0BBwDTqEVkV9MxtF/3vvSEVr
ZP/12q+Kn+87hXIO1xBPs0ZMWwldJV7k5P7NHIrIkUmYNC4krdBB8Xfe47hzcXjL
850pDgEwMaIEbE8/4kQldc4/ibzhgk5+/ltaL2YMqLhl4QwRwSN8RPKW1XrPEBG3
zqbMdshmCxKVtnnGXOU0l0IevN0MvnD9yovlHcHvHHwcSwF+UTwSl9e531oLonVK
jYp/PUO1juXaROiPLqpPYVDD/SyPjDyro5lzLiULf4QQlXCoLjRyzoIaIFl2x3hm
QLRvIGnfRpXL8QLHNyJxtm8xOgV2kbK/kP8FLz1QAWA719OPjIwSr+eHVsS5xiVr
5O3Da+ZjshYLt40UkwDjgCs6eXcMG20UE880EIPoG9A6YglMZzi9FexE++gQHmbx
MXxhicO6LWC5hROiFRhAyTpVGlpp0JfCaG26tpQH+4L3YLt2z4M56R++W792IsBk
WRUUY5MPHnHoxr1X5SbMACdrf8lUWXwHSnv1Q400wT5DQoJrlv8PLACDOKnHgjtK
34aN93BEdmmz/B2wU9soDfFQDD0Qkgyq3klhzu2vPfDQZ1sIyHt+HiAM2kPjV59v
0eqbbd6O4SrF3aRadT3jLZPqVg5OgdaxyxHi5ZP5JNpEBEgaVqo7WPRW1sm4JSUF
d0j2aJBCi0x3CQy2i3GMBNzi1HvoboxDCqL7CfIZK27BtgjpKMkGsRtAXeeEEbrq
6a0zWqOk9bMytQIsolCwVFBXQ2Unu1Bz1Ny5TTWtVK6SIJ0zha1eDn6v4ePJfZU8
jpE+2q8qWMtNA8egdM7vGdufcI/7GQ4Me2i4WGX4dWBnm5Yf9GTwrXLPTsGyjfod
2Gpr+RkmnDD5pXCegRriGTPc3bowrmjzFv0ZBz+u+xAgVg9w4u636Wx4stH+oh9X
Q0VRG3gopvOoTHn6b5MAlDDN9r4i42KMz8tTrAc1108vZALZbsxY7eMtnf9haXEr
aNXRcmj5Gb7d6b66RrMbDrH0QXWyN7FjgVP1yF7rImMSVV7nmDZpM453JkKpsuTg
FZdsjlP4ZXOSb/cc1tYLnf/paHlMpCR6D4WlGBDgtPa+DMlmf/d/CmG2/yoM8qSB
k3fcMc0904UCv7J7/Qy4enWenQgAuElgqBtStIfiQCakpsILA0eduFyGaWX4HdKH
3hX8KHzzW4+4ZIhoJdmO6tJKAWj4KSdGSDT5z1XJoNaBIuuyqkprrvyjwRlHEH8M
8JnH2RD6JbTV38j4sY/RiDIpH11UnuHNoTbVzDMlyiiUT0zlWJjh3enX81nEMsyF
ohYw8MNDlJXB+NYNOhsutxSsdTXQnnCqp8acv9Nx8qKFTjr8xBMG12xTh/VuU3d4
V3eNys+3RslFWWc0/dVdODG+876nD1q5Z4l6baUdrB27iB9Af2OpfejM8QtLOu4C
NXjz60lsUmLqBxErzhkmaEy1qT6pNAlGFNfm1CIIvYvRq6neajk8lN3oWnzC59mw
OMCrasilIHHpMJSc1TS1WCRLA/znU3ynUfpnDVmUW3TlxtsU7X5ayvAiBcbSn066
XyodmiS8nFMUBDNxai9B3CqbM1UtmMBJ7wYPqLFHr93yWQy1ihw/l8R4aoTIeCB3
vOx5oumJHHxUMV/JbDPPkpXNIBeEvwEfB/tcncu/Ttbrw/oMNY7GUFMmvw3GEO4S
C9xYazolyIAY9DeJggoAPVWB78UQl6Qubyk+J/XoSej6BNnbAuW+1sKZHyc0Poyt
69qvQ9ahb50R+FhZgtXiCdRZ6QC540RWz5C7x0ATUiqMoKAlYjVwGg++/IoYfaMv
Ljvp63XZ/9CI/mEuGNFrGyA3W5z93tNiLvGwJRTf6OdDj10gBYuN4G2oMmAIWrAW
OYFaPg7Lfve3jCe9UIQCU+6aGc41J1IJb71TVNtf2qJ9uqlpEhWmHMrryvgXAgWO
bboMNnTIvRoykI9A2xNaTsrC0zHg2gMY8B74zQoZxzQWASKMjOSOYtZTXASv4EsP
s5/hP8h8IrpbBO+jKLElqH33Otj3Lz6YfUvjn1qvcdyQUkppsmJVzGwnLshqI+7v
P6lkGh/pEBO5xUrc9M4z/21ffcGEgOuSbCNYTAc2eVZnPwgAxGjycc4YY8QdQQKo
mC8punfVfJ1bEpOWj1QQO5PUWXzE9pKEFYki9mVgGYimrNLIf+YK4WLSWPXBwwZZ
AN3cQWswdqQ0NoAieih4QLmoOJOjpUbkxmhPUufUZYsUDTtLlEAT6xnO2UyYqwj/
qr2ub9fHjyWFcbzQYdboDwW99fUAxAJzmHDgYk10M6bGDNR9WKJShT9J1fOj9s0+
UrwOmfPzZO3Rxyp+PS+riUImtP7+eHaZl1IUHSSHsCvW6933uIohyfAlBdEOpNUC
govYmj8yMnyDOvIfrMwzyfJ0MP5QaRBsepbUNgOdLwv8LwWt+uak26XqirzOjNoi
f0YrK9Kso/mR7XQ7F0XTApnuVtv17shsyihxfTOJqkl5gmuHQMZF3/LaIyInsOE9
EUGuixl0QB8bI+26Z1fy9EWwZ/aAQpS2Gr/6hHJOT0op/TuqNxT5uo10wntOGOFs
i7TtXlapF3ZmEbXA1ez1Gj0XjSGc7IseMOYK2nh6Npa3dzK8NwLxFEL1cirxnzxh
C3+R4m6Bh2Gu/8+H1YBagr//5VMGKIj9zzSyuuXn6hzst/J4UDHMXWQgio866IHL
ab4o8y/I8LUPkEl+aDyEvUcGh0uevAwIgsoRlj98lEiOzdYKSEaYp/zrmXEPsC8E
YYiFHvP72NVksWM4PRMYkWlTSZAHOCrGr7k6gyNav6sMcNWi9+va3vDYjJuTCtBw
ZkF9bWhj++pnyMEIyfzAJE+Wj5PGF7/sYaEkQbjqAXwQR4AtCxxBOsODP0/R8+yj
wJCTQcDyuL9+4En2ezWQX9Q3vRe0wPA7XpW+iZd7j4TXZ7WfJ6G0cla4U6G+jPmP
Anl66Wu9J8dNgGlZ2j9IUWFK1Z9gTaWOI8THRpXRfI3ZQEJjHuwSUH9f0+f4R5Dz
dqgAiv9WuO/9mRl+tPnShGsTZ7MNimldkfK9YI3OeWW4ONXa8VW1Or5JQHKjMSB/
/y3HjkZyU25bimiE7NbyOJJwYrmkpUO06HuC1/T4NXfQAVZ57OYwuSvnqYRPpHa7
F7vsRrISXM0CNwuc0bNzrlnZ8qdlQ/eHYWx/XTB2TUVzzu1eLmX7uL5DrI+l4bmT
EdCfGhg/2uo3U1l97xggY0wh5cZAyWgqA/NhIk0tLnhUW7e2xIxvmfzV6AgaoTt4
ZsHFKm12P6c26Vun4EGvDpKk2J/YcqCNPpy2D3+2xYqkv7h+pTxhlkUJiK5JgsIY
Z3Ju6isZhpW5cPOZXZqs/kA8BbFaHU3fDS6TIAnEXZqU3LagpZECSbx6ahXN7Q1X
P2RxGdMhRMxKM1MErBbmT7kw7QE++ZOa0oyTXxXg/e61S4OvYEPAB1ZP+z3W1ygL
juFsRKK2glIpyBeKTOy2XazdiBNHMyDA6JcVHbOXjUISMtYkCzF7Y95g761PSbrB
E/LkIr/gATZWYY1kVW3j6EFXrzOaSylp+LWZj9MOdlT0uLU3xBg9EZUFK3JuoiMk
M2gyNeqPnrC8X6v8PRjLqjNbHhdLOEBLUHTQS4yQUzpvO1p/rW9TlmmqJdW9Rozv
7zQdxb4SReC+9gDjCfIf4ptXOw7WtWwtL+ObgyKACK8Mi/ZGaFniX6CFif86cUjw
5ERTKE2ME7VHxzJNzYN0c1kcfijF96/UjbGWPRnHRGGgfbUbGNXEb8tDr9Tvosrz
PH4n/w9IManz2p0fo1VtPBu80VVyLoKBunTgxSpChgH37r3iPZC7tdr5KpAXe50O
toNPZ6jzsyoxbn45r9bAfuXkS2spZF/XnUSKW7aV/9/b8VKbBEaDRqAEVfI5bQng
9c5SEyEeifxI2BUOA8er2R2Jcj5e2R3+dehdrGb6CdmFtKa+9ZiYppBeRhOpH+XJ
0i1lz3Orz3CjPFNyQM4aA3j1x8J3Qxf9EjkQMirP6xfw3HZWHS94CXOKugMjFa1D
csdz2y7Ajry4Txzab2+Ot6k5RDDvRTzsy6XBxgqt3xox2/azakUY7zaj4bAzr3HE
OFtXOZXjPbNdvxzkFaEgHjqm1ldeDE41uZV8T6le9p2HFtiIy1LlE5fho8x1G4vB
N40SpWhJt9ksiqfvEDKeCWmMRGRYYrXYHsJf1hxz7JI1co1HTeiEh5sY0BR6HNbA
E0hWx9f/aDJ51I2gPrtBaN/QN8F/sfBQI0M3jtlqjNgL0yk7olUAtooSRbYanS71
7XToZSBOaSLtygcgjcgFqyn+7DuVR0LodjVuhLAC3qGrmrFCNEiwp1x/rL6pI7ge
YssW1iRtpCJJw+c7jcMT8EWkHSEoOU4l5xpAZ3EcjkDaDBjV4Tju3CokUYb9Oqvc
rG1ukkaLrb4m6u3hQ09z4nCmxUCIpsIOo6gNyobbZvDglbWI3gOUCmAMyK5lZuJb
Co25huYuW159qV1/UGC/18ZXRHu1zo8KjBz3PTT2YZbhbie0guUEwVicJ6BTPyBK
7hiCl3B4gn7gY9DFE2IJ9puyjL4lxTLxraZwoENdt1U6dpv5PMV+H2GfF3qXNJyf
MHxMJ+ayBndlVroxwFiD3Q3aHAanNUKME3CLM57WJb9fXURqkx33PBGi+gqYhkmb
QkREAUR1a0w6Kr8iZp9WMq2qkDfgrAeOSbyORs9Osm1grpchdZUYJFMOPr/aztGE
JZMmzHLTRaUhKUom/5fqea7WnBSDy6UswYhHJRyU4FmlwX9LOq2zXFqIx6yPWlli
nuV1tt2R2N74aH5j97Vjh1bcdKe8G5LJZ2mnhR8kMJnM2QrOWjyd//6mm3c705YI
k9/0mHgD9Atz01yemVKRp9UWI2vXphdR/HJyVn6GJI9Gn/XB26yKbzrn3mQ9AHTw
YoX7NyikbxTOn7dgdF7J7uYuMQSy//5CVsKlvFVes09IscoUq1CVllaPduJTApbC
juuz8+XS7Bl0l7AbiBGAA5jJeMJZs9+7KeetUV0+EZ76pXwXJ97dfi1G0f9F2Bwj
rs2JGFPJLgsk5cg70TLEnZOB9JJz/B2cQbE5wbRnQKQZ6GH1XX57bfGwFxjO8iTp
TYYcIfDc6dnzIIA6lt1EDHCda98x3VAquVaDwOxyLZIo8KAORqdMlFndY4tPmYCP
G0pmBSjZF7apgrgANkZSohWjTCCjPj4bF+txwKenkb/nseVTpkB4fBLBGnmSVkq8
qx50/dm7bmIUgl9m0+RzTRMahrex7deDrdaCL1Dz9+P/xUhDHUlhJm7++YRsJ6UU
roHc7T10Tp7T6Sqef66BE1cIl6aW938AuoeNdNgnpr/u20PluxodsGLG7LiAkfxy
m3gz5LtudJumOnIYCO6BAi/Pqp4WEZRNcXjhl3FjklUCgeJQmnWYBWSY2xlDdOG+
7Gj4YLLSNFhIRcZUQ885wPAahrMm2mTF3UUPe2s1Pvr/iIUoSan1uh8FP+a6eLeQ
h0pj2YHYObcwoXAbdxme5EUpDjMiGCPHjofLQICMcASIDZh53r/SbPqZDB1xhjFL
ezW3M0fw15pG7GnAz//MH7o/fXihAnCRAo7DMFKvXWw/HwMWVhALZTEM3BU1mx9W
uvA3zP1qkhHiSfuKb0KYBEN8IaTjCSL3Ur8CfuZ0LdMyN3nj2Y7DfXFRf+YGQAmI
3Ufriv2IsTJwLlCRVtd+/2Nb0Xzc2B4vF1AP3Npgvyecze4zuzAftzXHr61M5u6q
Udr+iw7KpzPo8KIWWNzLt0CvWwwTe2EM8R5U0TlHbMKEM9a1Y+w6qNOTxfO+H2pV
EtC0N3mqxYnwRAz/o+51nYBnw50Fml4+KEEUrQ1xd0v/DNBKKMZ2TspNKBAF3zRw
fkDeUaAW3RkNKi5exAP4IgwjuGKgfkgjsHtt71BBIafuUMbkeqTDuw55yPIVJCSb
jtHMuOvHZbUNf0ersx+18lSGSGFyfL1HQXTKl3H0rQvTgNLQqEFJlgrQX1hw43Ew
jlvlVGqISvpUQVQxKgIiyfUzNNirXRr4pL5UyFwSW8ux5J/viSiNy1rGHBpZffff
bN4IU7xopNDQWkSoDWqAuaoEG5M/9/tLl7zBBoTxza4D3Q1xQ45lvzjP93cmlyMA
/3DgyWPV0KnEosyc3efBlUVZ+M0iv+SiLkbIKAZweH3E35Nrh4fm83xfpzmIxI4J
UuHPgDKsyLWQCYxVi0tiVbQ4CNIwaJZ6aQKPxRj9m++PPDAhgEKzph4E4dOR8bFq
OxKO8elOBluZrb+TKu4+3hr6Q3+RmneXfw4LL9wnTYq5Hj+sLF/3ZPvSSRcoq+xL
WGdGqFNZgmgbEtKPX5YDnc6+Vm1xMTK9ZGMHVrI66lAmMME9EbNCq81lep4AyU15
5TC4xZxR8GWe/YP6TnF+r8syl5MDnKt6J9SpSeQt2nDr+0yxqA8aVijcfScim1xC
gi0BxIRL73IFnGP4y+k1W76chNQFo5AQ16nvvMJRoZF/NWTemI4rG/Y99fJW7hbz
Gd0dtB1bQNDL80A6Cngnveg4D/l199s9WDVwNkqOjOaM/SUTr5TmSVr5OrF1CQsb
axAEZrzjwVsDyNblN0/E70eBd9UVxs0Kvx2NRIGU5uaYAWYft6EWsQZr4knP0Oh3
dy5VSgvJGv/eLlnlxbWHoEUM1yJC8QygfHm81M3nF18dBRVtN7bUYkDt4JSI35As
J4AGR4xODtWEvyOEVIBz6Tql6z0Ba0Eo7J3p3sti206shODexmaP9b/i3MXAtq54
FcfJ4/hCfeo6/vWTSAxg8ipnaMkHU+MLgf6DrUBoeXX6btFD99D/N1Tmyje7CTG1
xP6UaP3fWB8u+CAeFLfzHb/5Z5n4Bk91lVYVA/N2789FwDPo0VfBC3YjD4pVXutp
1kF4XhO+pjUvVj8gjYFyj4uTRuVWJR4Y5h2bvjmEI3018Kpji8IR3uxmcS/7B83O
jceaup31Vce1YcKlErXPESwJR9KLEtT2hlPxJ2ImG3YR4sCHyaqjW0hesto/NA2a
94uZ/EOEFye1gs0hCnGpKDyUPUqrUsOhltvDACCJNkdKdZtsM2cOh9A0o6hIasT1
aRygALG9DdAfXwitANm2Psy5sI0atWIYlUMblX/sfZVmji5jQGkObloC4CKroN0J
1rs7AN1C70M3lngT9OXWNZjYeTikhhUzQOk6hjA76G6T4MkEtqFPjPzcePniKhmv
1WzFnry6vsRlirKThsvazIRf5zSrpvjCo34lEX2pb28c1ch93DcANG6rPvYg2xxg
S4kL4Fxk+0IPrd8184QwzFs70d8P/B8zJc0pni+3Kx9t8/SOv4fRY55K7f8Iuh0R
5x9CzeNQvRuqBqwJ6UKYVaYUZ2/vD3jP5qmm0NLu9j5QwN9RugEzkn4YjnGRIEoS
qOBmN9WViM99qu2BXvQ8aOKPB8rkpwLBeMgBUOZr2kuTt3PO34iuGpJHYVZCXawn
oUB6KA9oa3U8ciFvQCGHQR8QmujxptbCh17btqAuGZ3f4HMGEfW/u+LZoU9C1XkL
m6ltfbnAnhbJ1t7D72y2yx0cWGR57rOOKEQICk7/w6qEjqzxAq+dwNf4TwT4cZGl
bNryNWuCx0yuqQk3O0blRWMb0TEmcV64KToq4Ll0A77hMpsQ9wx1afepFhK5g68i
Sc3kc7t7X57m5vNm+2kn3IQt8qpQAL2PatldaXByBxLyrGCDP5UpmJTvZ9X5iuwA
Pv5s41bOdxIaX3y95bXQovWYsTdLJ1k5LH9/QPbmBoDCV7EkwKgCe5hyBS5lyIhI
+OmAOrxBwEf4tfgDMzqiEOEL13zlb68utEHYi/4RNGstrcvUKTCuOCv1Zh9Mlj5F
/M1piuxdKjRgbNJMr2j7xT8W8+g5lVdITM0lguA++ycyuESK86agkeXYPo0Y78iB
5JQHhbrnMvhJBMJgzflTgkat+REJKTGo+ZAb6bkFlE0cR5eZuhVGXK71jyX8mRqF
m9mE7iNI1oAenSWHV3d/4qt1ByBAX4Ms5zYL+q8IfWeP/AQiiVyZyWX58/3/lZpq
o4cdFo1ZNM84eUYuWX2+EZTdbU8JE2OCPO+8LKNPkMXtJf9mU0wWhGbArmDxHp+p
g+VRMRIm2VwyG4TvCTn++f3pPdqTvMCxykIekORlXG+lsKs3bK2jPjqGMq9uy9vY
SCCcvOAQUUkrTO79wdCqyw/YmWEY8ferAGIAc0dx/HN13kcKeci3Tl4RJpcUAGTB
TCWSRi+ZZFAyJfcFbPP6e6EV9g8M2mH7aov0eJkpDuNIWkjzO+gF4xiKD4G7IQwK
e5G3Q62V4Dc5jrAfmZxv8mYN60soIhxZPFp1JYY2upKngoOkgXqtFi4Os0j1Fvaf
PEXsAaQORP3wp4Qm8q9uSijjK/3iQXPyCB+jfKh/05BekJO+5oqx5ZuFBa9/d0rP
Ynhdp9GHQED8EUisBwKEaDDcbql49752Exba9gntcnZaLdjbCxq2lakVVkeBx3Pb
ZcGvs8kMkdOoBFuUtB4NB4bVT5eNaSCIRDF6f1ipD/nf2ekXEVU1lbhgH6ayFHld
w0sRZEmoKTpsKUEBtYmy1KkHtO199/6MiGyCagA0o1YrGqvtMyONskG5OvWAnF3t
oXPNfMSaSHhwjuGqljquFauceH5QvULj/TiZ89eCp+jWjsZoJNWYOS2RxpBYkcwl
RXnOEQ5uGpYDeTzbTKX5UTW0pYZ2kA8WExoL5GyBGQe3x6S45u01qQrxOBc1vSOD
3rluKlpZCTzJQ0zKOJQwQ3/RS1hei/wp6hMuviKWYA08HbdTFEaFKbr1Eu0Wj4oZ
RhO7QEq7q7xKbJOqHqHcnLfd2h2663lC2DdB6RByoZZfkhngIksD8tgafycAKidj
EoZe63/ZX3Ljq93fkJCCCR2Ku+jNNVXJ2XN1yxklhvUsCKTIhI/C7tTxMTTnyMCh
TycWKljNl3YwgxH8PuW6gFII9LUNuQuSglKLIKFJFL/0KRfgyjge3HMlhKpvQQzU
TE1ZfQMBA7pUCDU4etoUiIcJkQTfxERdAwLc0/ZKRCqjxtFtpsG1nP4YRvDefC9B
dM79jf+0uXNnAafk78fBE+F86asgSQb88L/BfSQBwzvR99YQSS4higIBYUQp3mAc
ipczHwxJq7g3AWL4gAZC4k6zEDv//YB+6GmbPVG75fHhPNlp55Aso+aL0WWESd9m
H9OnDpGhHpVz/PwkIovS7h3XpbV73N28Mjjco9uvZg1qbABdysRYKmgC6offX5cy
XwjwZR5NE63psu0gxNVujzMAP12K4F0AwCsU6X/rLzR19RcPh8qFKmUTauT4SeXw
mMJGnZgMDCv5qY0MOSZaFY2LBTy7nJLdk3YgwS0BAuee/e6Xz1OwvBVP1+Bsd0QE
ZboGm3daeb3MQuCtbNIZnWx2C233RQ0pnPWtKZNJCtRA8aviMKX3wFw2/mrLJh3T
4i1h82dDFCzUQdTyi/aTHTuDYaw6WWQRHb5KGcXBYqZf+pILTf2bpeefaOTPGXeB
TFtRKzmAxWEfWph7Ip68dqczipJIf/SwoSsicJfVpepx6nljAYAts0e+4GmdQRNr
p+TE0FCa6X0GQgxOXH/j6JBmbm78o9oIddOYPHA/qXZ+fHIlGC4l8KdJFDY4qFmR
hhihkuRUg4WLdw7ofBP18JVBK+bZSzP6/M+jvSZJGihsXlTHwnp6jeKYVLzGQz7+
HTiZ2DmUPsrjF3wcayzXH7ZQl01uoo5BUBzi9VPul0Hp2YoiT9EDIE5RLUyMDYaQ
6tXFJ8jQQbaWD6IxlXb6mPE2iTudAlkel9nYkpcvAoDZHfOOxSlxN+0fOBqKfgrl
wpjEp5ckjJYSVAjdEtGdgR0ezDzPr+OwSdYPpyg4GfBc7K6yPP062HimkL6KfLLF
m4pRD+89MIpV7OoqBfCHqb8lbI1gWD7XdmMnO3QgKEC+ciOJK4elX4LPskL9dezW
a8Kyp07264aqAr0j08McSDL+D5V538XNYsS7oSjx2J9oF6TOYZPb9ZNfC1OCZtz4
WieK1DL+uvCwk9rZRxpvunXNm1Je3A1lncd2fm8xQ/FmAk/3XxTXbnv+M5hSNABm
QvTGfvTXd888jXOrZb5SZKoDg3EB28QUQQekniziJQ6z8HlcHTQCjYkbc6RW8uDU
mfgOFZ+M6/NyOuXAFAUK7ij9NOtf8aeMGU4M/N8Nv1w5GCRI77F7toQf9LJcK2jC
810WVOsXiBCYuIMvoWvUkdlwMbvQ+mhQCjrR00z5NBksH9IHuYdKO+GI0Yj6BXva
8EnS2mBBdCRRLVvwJwwMtkEPi7mNjU8Yc1LYeKFdFUPJgJyqFXsF5KGR6lICRuLl
C7zgdr+K26PrZDj1KPaqERkGOq+LyfuRDGZTpNmhgQR/s15XE4+fFurROYryk291
mGjh2bn8PeZVmUTOiAlxPjpFUENKffT1/H0X/Y64QKcG6LoogxnyZHcOZFFs6KlE
XMsuLtbNUAkOphLlS9yIu/ZSSq8jEpGkmM6MnXw2u4ukEHnJthy8O/zNS/o3urFp
v3s47DoP/lS5Ut2U/eUrwu5swgG1erlbJfeoS2xQ77YuhpwrJEd8Yjbb+RRt+7jw
Jl+peqxLcSxWE+orTAsFaHX/0Q7M4OA3VMPaZcGaVperbklmo0u1e7kUdcCpYDCo
7/YjqwP25p6f3FhoyFdCiprQ+PUDIYlVBPplaBeU2BYBF12/PR8Wa6VPmHSSKwbe
UqJpirg02PoDvwEi9xd959O9e3tISkeDu7ROpFh1OOSlqtQWNHUthrFf+ETBuL4t
odISlpTPoxayyAeq35YE5VGL1FcmfnzgFWZIdDfUX3+UkbRf+hwydDpqJLsg8Q37
nu3GyixGNxNJCla079HTyvfkFKHLMBjCD4wnc81dI1hBlOTToxTY/4l3ucZHZo7z
XlHg/pnl/5jzxggDw5qCpiAwbqszp6/AMLu0Hq2A+f0nB4z8fMalPpRsBISll9FS
eT3Qn7eOK1f99ZEuFpbZQozHPXbdXhBHUSDMUh7lBpgoTknnDHmLabT+l0MLT1ss
DZHl5oeOZzxDFsg5aYHHGUH9E1ixVmquzy+X879NyZ5pcb3TU4OHPqzHKi3yRJDf
+x+RcakR0WdPHtf+uZ9J5M6dvGCC8qacOS4OebMi+yOTmRlkKsYeVQ3vsE/rkN+j
LuTevoDgyacfHXrbgrF9Ci1qY8Xa8bo1KpdZ7/ziS/edmAoKwXFC96ZLOgN/PywS
HdiR4Mikw52B+ixoKTqUsJr1FtK0dkKk+z0j6dflQ3ZW3WQTXbAhKMPpbRLcA6m8
hZ2RMhuQHIIBo1EN7kUBV8LWNezF2qCbe1HZkkZq6umY9pxYn437LYpc3zP7ak9i
dm47sK9LEpXIfnl89VDzzGMW17rDzYUvFMi5XW6N7GGjFPSNzq0Xuz6V7nk0PSvg
+KgP+4SdraCt4DyXTFzkErWb1Uotr9eX763qScwBsCQ1ymeMAxbWIF0UKKzeF1MK
0BWku2vX6alFINJgHTElWdKjvpmqiaxTn8g1/KmkNeKpjGfVQ0hk5FuqmvHynv+S
2SjGsnl9PVow3CgqOnSngxfBiOvFv7tVUYAIxzzAIthObP+4J+312HKCp4IompZn
drnsVfOhuTZiMEfrV/DfDQlZ5PvCfEwviIJ3gnZxTCvsrpYjGm3rxdVT6QaKCz1t
GUrt1j2AnmfUN5Oh+FMffi4XUR6tXC8BENx57/D8XWfvxTWljcxMtCQyFw13mqJ4
t1RmuS71x2lZp2Szw4wot5+d47ZUOuEsFvirUGSExPiwQXL8luGq6zvRobFRYs2p
W1ljGWVSn7u/XZv0ISajqbVYC0ubghz0gS/TGRMSUCL322uC4lEVDfR4PlQQSXRu
9HLpj7fNDG/jGtKkkwfyC5C1niaK2+++b5i6uKwIUPGLePDe28SkHky+QBdgBh+R
UKqQ3btzZybviVuq7Dstm0xylr+XMIbQ0nrEiuHT2cAk3Wgo1cRv71uMUDKYEp3c
xl3/dESyKIhKuicMoFG9GJ+azqG7UjKRZEAWF+QO7YVtjaIqkBtCcfJ2vKZ/4NOr
YsLj8VWp6b/NsrrzKp1yBqluWEog7VGAyJMeVaJO9VcTPXsv5SAq1hFP6QeS3Mv5
+ZOmj/uGpnSGiOANGjf4YwWE9oT8AbRZpyw6Lrh0uSfMAXBFhF7MIgUU5Tpg5PSZ
xhjzLZDraMuI0O0AgiO8Nr3iMtl1J2BSOdXXLSw3Bin62NAa3NKqMc7pPUqkUAUS
UmM7K4idavBb2nr+eb2UirdgiJmbICKHGHTcrc2M78KKh59xUCXHQVN4BpdwhbF+
g4T+Z1YR+1/Pt2jHxFIBZ7pJVFrTEJrCE/BaWgnHl0E2w6gYfGxud+qQHgoOEVDA
6nrV1iZWYdjvNRq9hJjRUMvzlh1l2LYRcb+ZX9/NjIl9+G/YdFfunwV0AZNZuqbd
1UcINRwAtVVAQuBluVqwrgw4v+m5DkU29vOpdhX4WtFtFO5Fbzb6PGRb+dkz/jU1
rUm7yHi9rCz1kCJOa48whe8jlvJpUmzOZDFLpkMaQ2n5j+WxnVtGdr+a4jizhc7E
uaIec2svYPKCtu8UhakApmKG6OQddUzY8Fnj5pFRJXr0SBTJk48wO47D7TA0b8JO
7eVIkz1EwxzgOTZEU0UvjrI1Kqfo16nq8tY3p6RvA4m6DALf88IefwWFOiRRs4Np
ShRn/uXe065diSe2YeYoSt8VNyI0Y25B6A44Y1azZrAMI0b384AjsTvOEiCJLNvf
1ycRAYu9SWDNWKU9R7/gon14Od0/E/5oWgaNjFbuufaRKiVXsr/4GsGuxZLG543l
yd0o8UXrxYkQX5l6j8bWyQWtwrnqm8a0Nwim5nIe6KJcn9JaEtfkg/K0yVWX8CJn
o72GxscZEGAfsLAa1UkBjhvyMdEEXPRJJg+uTJWNVHJFKxNeqjGNeNMmYHSu6gWw
ldTaS2FhoPV+mVTMWTgWNyQgZRw/meyAJ2C1o2SL94OLslzAVtXlFa8Mfdzqb4Dv
V8etIIZkkeS2nq6p1GUbe5t/f4rkzDd/Zy8DthnwnqMHUsyhKSt0L31qDNe432Mf
5EskekKdvOmJiCM6/uJh4dF7yu9tDIZ4WDpvSGImldnVxTp/opv/4d9SaVQT79Ij
6ttdpaanghlE8liDvpx8M0LlRH/6kK7q02fQlu6xqT3KgoUMzv5NAxawcJBQ4azx
yCbVcV+hUNPVAN8qWBZarKzu/tqPC4H/5JwKfgPqfjIcbIDuMcs5d/DCysxbkFD/
Qr4J+yo+eNZsTGCTLsDm3S4gPJlk0oFLm+BjSCa/2yOazOC4L6AIJAbsH7MDmprK
tT1s22K59uNGpf19vWvNoBx6aPdaEgg5nhdoJpN0KYlLzux188hYT/nZhyMsxJDy
yRqzxIbb6+H+ynFI0dUHFIUyMjbx4R2VLofqnmHgzoBSLI+RgJoEFYjd3Qvqpu3B
4krM2Wouttn2q5iD+/UydCpVStehdKcnXS/WMQGWYZ+VKfI1aEqv8MaT7nwYdlEr
1kXYCyOi7dCPyYlNRN9A9QdFu6tvoeZm4KpVGA6zDyzZpsz6PL+QkkpOQdkB2mkC
3zMUlQiuHzj4tRB/pK491nxkV4//mAYCZhK7Fxn4pr6PaIoRm0FLuVCSD4+glDIX
Nhkn+fEdcmaT9HuSAweLDPBRs3p/ASQXj/jdZVBtLUrnFz9m66t6HeUTBPyuTytP
P2+KiGjZ+ueC4MjyWsKKUCNcb1CYk1MPeBNiGpo8sTZq1cJhmwxypveY6aw/1XdQ
stbZDdtHb+gAL1IDQkkqO4096jTkIMrVfIR+9owlBKhD4j5Spvsf+sGJJ6RJ5nWI
XMxifOIELoQI5vYG4ZV/jMV4vzdOnT2ePQ9sZIOHNOBdM7I56/NhbInb/orUIRkD
VCoExWgKHsqpDzLEjGLqT7D3HtECtePgJWCJ3yQFOHChDeINpT+lmBD5NDLyiJ0O
+mxRxQlceMWgGxSi2aKc6yMrpwaz+9uvbl+ahgrGURSxj1TRrUt9iRgJbMlRMhzI
ksxLJy5LtyIhtouxea/reiILK36e6iEoutj/Tt/t1lCwwQw6VQI4sx45oFKQRoEo
mvY/iZcryzCEKWdDNIWB2U5xaGF08JGKqx6f32No5FFvUp1YoHtyCmdm+xGqIj/+
eehQQbw00tglM+Kv8NvIBsnIKZ1WJ5jiHq4vu3+ScL8Ji7tUSR9fnKwnDhI56lYE
9GoaDgbpzltqlly+xQd8nZ8oxxeVNBixl1HsJXpA1lFcHTQ418qYlqW5fji9JJXn
TF5wNKzcUn1mryHqWshhDg7Mvo8rx6HRCgA67enYwXTXkY4tOiABFnVOqrktLrtX
qW60RsYDEBZYf+CWohaUSZ9Tf1qgvByRKuHx7uGR9PLZ1lltIH02EfC/DWJhwNBw
96s+0NJru1sDWcgTnKtHvbKJCBZ/Jk0JeDKqsAaqyyhHe0whSR1SrhJmm+25KGQ9
VJPEEkpSEHkeMkoRCStLm35j6sjPK/mL29do6B/RcYJbEX3omxME2KHOyUFZZ79N
JKx1f/ovqZ68cUc9Bmzgu21SnXYDoruvQcX0oPViEN65vels0txsS+Q7EpaRaY1D
m5Kbr3JVhJ/ZydEJ5IO3dr9sG9WBN+YGuRnjULwzLeEq0jbxzPuB/XpiIHKVGycG
RM2uP8Xni8neMnqkf+0m4YUfsd4VLwvopwCeZfsxNY5isiGCPCiA3azw0dPf2mRE
Zh8yYuQSG61J0B9HVD0oXMxxhTrNZJPg1Uuqo6+VnfHDqRNbRCDTBWJo1uC1TGDA
eArLWEoXmwESIx7U5AqA5aKyp1G0K6/hdoPJq4rt9LQJMSHBiJVVKtL2vC+oRunP
/bjROLycNhCjCF057//UwvgaxeFbbKbI6aNS9NEQMZ4Ce2ARrAG4ZbHVsnU6TQQ0
x/8uam8wvGeihx/a/6aMZcu++jsyRRpHdUvx6KJixWHLlubhjIFwFflmDuSlaV3T
M1GQOwQnJtvzok6C8+3BqedlUb5WSUVL9rkMHHU94Wkyh8pQNm1b2bsy9531iz/+
3TMyGAIO+tzx5Ci5D3289NfTKHrdZJhqTvrxZLZPfyjrwTdeU5cTKiA1kIwH6fsJ
tsTLdH0YqBsV09MFUKgzMi5TBE/WU9N6zXXJzYVw6+DW2crBxwnoQ2DZ/KDodti/
W07RQcupWEQddjvaKQ/8lnhzW6Pqj9YJ0dRFuL7ZFRcHZJiyx7ssewsMytZksZRx
3h5xD0M2+hKQiO2xNrOwXubrDJJevohsJ1S3YmI7eu0fRUgLJ+n80RYyKKWOanCv
6kOKWe1I9vZ8/9NsMJGlqGcWFas+dVUm7DR3XppSy2Kc30zFOlvZ4owV6T6JRDkX
ALnJUYrqPZexb9tjlHlZM4GmR/rdHflBL9nRwCVmTqFdUChekEeFZ5kArj8EA1Nr
dTymfSvVwP1U9rwjCbQBelkxg4x7ptay0FyHdS4zD/mXkyvfMpJlMKDcu1HlO0HC
nCgbaab/pbEml08Sq85OQ9oqBrXwTALpvBz1e+O/meHGHRF/BxUieCl2MT1AZKd0
+V5+8x7bsrdZnlWWGevuIJL3G5W23je2skIjq9B9DClM4dA6bBWu+zFK+UPJIUTa
r+Qt4K273MHgT2d9XJXEjqDok2AcJIiHgTkE0FSudosMppGIfX4Yqc5JUZH/g/2V
b4FxdJ9/ygR6xjfRg6NNVTTNRAbbcoVR/If5UXdNOMSfktAYGXxEGpMdLFTJ7IPf
SWnlSbpCB4QfXicnKY/3yNh5UfOKxWg3bbLjh40WfRP/RJv+TSqHAoVXKcrPsz1b
MWEBLSP+0Agm+YxQqPD+9LP6JcyBxI+7f6dk/qjo6VRvmZZLaTySloosXU8J2aLg
ex3Y67DGKaUvetU6gnncUE1CMjnd9MRmkuevMJhApXmrdHsHYOtYhHtup0Nk3gAi
2oy9iGdt/rx+cYHE0+HFcwyZVbut2zdFaqcena3oUeOOulpcFLM19w1Kp3MAGHwr
eRosXzWlWXinIN9WEbp6INorNsg9AnfJ/VTLSBrhD9u1ButGapKxNXEWNTwQYIar
yCwYUMlSQ+qc5Mg2pTv07WBOmZQl7lNDhT6enVKq7ljYkyWSHrFWyTKI3WWWEgRz
33UoJkAvCM8PFxxOuDXBlwCo1goN+CvRN+9K91pHWW9WzzDXibbLST9xZ5Izo9B8
nBchdVv9TzBy14XqCksSpBDvW3r6NIdxIaH4/h6c2qK3XhQ2gVPBVZlSpM/Qp40V
5lahCq6l2oQP47boTLocimTzN4ks3YY+EiBsIA68RyZaCTNd2cHZ3TohjdtmBTf3
47WB+4N529i9j02DQIbZoovqhxvEjHYQDjom4PK5oAdO6QLaf68eTYx1tzfyNLSf
i8s6G6yD8dVyYpWkoJCu+1quusF2eAAGKGYZfPsimzAMPl9sU6q9smCZMXQDby0q
Hdchs+RI4zrQ62BC8UkrnLYwA1PTMn0dKPvpYvbK/CgWgRfzrP8+1vERR3436raV
gTZTgt/eZpfP/YfZ1Is98asZujGYic03aZ2sRNSNqSUuddHyWgaWCIpnF/39DHRn
R1z2o9Esz2MHrXNVA56RiIaXYJ46fzjjFZ0SW2IX8+Lj2guFt86QamDbeyWmVlO4
noNYobisHhf+RuZx3XzWBIyRBOHsHZMK27UJqdwnpCDpFugOMInNNrn/SRbToX7o
culhAAyAYP99n1pHjjO8bXCOdyspoiHxHT708OVLOFB4HXonD1rWHxrduQ3mEofY
bQYAhJKhMo5LvQp5Y8fp4jC2y1F1jQt2y57X+aoNKovVQtq1vaXqNVcTGVAg4uPp
qQYHPO4ZFNXNuTIq5OMAOIqWhnhxan9bJjJoAreBoCgAtjGYUBawXOQCiltsKzk9
RvGIuC+Ib4F9qwddk7nyjcAfB+CNpnfArly2hJuGC5AqXC8k1BPMOANZFUFE/IyY
viwNyDIE/Nk1pSQcBj+rhhJxxoIC44oQcUbq7ffv7Gi/64GuA1Yr0TEEB2jHsWqR
pm91nDwMGwiJVJ9syyjHTI7d8K5KA+QlRss5KjKKIeAY5kfbpHJOB0+fkMzkmd+M
AzFvVhMaGyiftGdLitv05F1i+X0JcaSaSdrl+lBPgZxoyFyqa40+FrmK6aYJ25Cc
+Bj2uEtpjO3cSSmSfIi+C0l0+Ekm1t9EYldu0NelK9AeMIfCSGiSPP3Qi/5lCmiP
dxc2vG0cPn3jMQXZgHNtaZ9oT8Q41Sqa+dgCfiTnyPsWIBDlDh3cJmArSHLVYIBU
bdzp8bRcWPXz389KNTVVuV+8qgUbDgEf9MWt38njMf/SYb5VKjp4v3jzFEQmemqf
9n1TtaIU6mBWEQLsf0jqjAFU5JrgCGw8+E6/teri75KvGBRJzxU+ICExOwdaYSzq
nWYWoEeIDPB/3asDYmrg2B0mu4QBXg0XCqaXIhLgzDgGOn+P81Ia58S7XlICwfqB
gz/MH3lMWmTyE4uu0U4bAxjqsl6xLXQ4gYjOpt6sGBBUW730SO8kwk8RM00o4Z+U
kIfya7KJ4dIRJjHjlcga9mhuM1825oixUHc3qTlhVCgF0DowN0vdyQAxsK2SHQk1
YzjPTU9DWMNhPbh9bGGZEPLWaRG5gMCWqN1BIc7xPZMdQ91Q7TZuj9EFKz7q/CB3
Ib9UrV6CW2tytPCY0/0hwoFwKdv61AaKhvWVKyP73O5gUZ4Dw9yhFpgaYtz2stRV
UKjpp9CpqILAy9MT8ED76motOYfKY94iKSz0BBBvxaLQos6XWF/LUA9Ei7Vqlxql
oxmjxjWtm2u8IRZ9CIFgcouBol1FdjtkOqLSPguPa3YCsrXEywJS77JWONkDlI1Q
eHfHPyKVWFa7PlWihM7t6wTGNtdCS67hafn52utFR5CmH0YZJqAGd6ldlQwgi67i
kz/irukPsuXI9nhOPm+YrLQ17Zo0ZO+8HuGbCRuYZqw6WI3/nwzTRuTLYsdU+K4L
vB/L8jLYNIFvMiH61AwPpET1gD7N/DLFOKZTxsLglwcy9REZ2ZDiYzSJr8WDxcuP
IBlcS+FPMQW7rnyXdHo15PgZCD0iigLhIeiCR70tZH9CGKWhK080KsUaJVN+zxp9
aHLfBUTTOYXDeodRt++NP3LPlzGe6vVIs56urzzraYniH+/YWOtd4Pd8ANWa5Yfi
jS4Wk+pf8oEc6FVlcmMzyHY2N55xamgFz0DWaPONVXe7gM6N9vCLe8pX1ru41m/S
BJTsKlI5NUG4Uo5Lo3KuTiy7ABWVclXBtjIpwYcxvFhbBj274ph9ZCzJ+PAF1wEn
k4QnbQl+HSu5ZWPSRxHFZPrDaSxxI1bFPSU3EegKTBRj70WOfE5Eecf/AaxqPHc1
DPTrbBgWnNYdqy/6ZRcVW6ww53ekjcCL22ezcgc0GVZv63XKa7lWvsUuKXaQSroK
StT2cRxsD1h4U9t8RdhreouaEMrwOZnWqUtuDxZZ4V2HHmPNHKB6E4F5TxAuCfV2
xAmnIQx/l8jS0uP/R61f07D7qwWijeQJek+o3JAwiSI8IEN/4KWQH38wHulZjuK9
8+kVK18Ibho6pMUxPEngjF5w+DKIE6YWIs+MhTKjjvVA6FGFlw9Db5MPs/+w740O
lLsKw6Y/YGxE0IkmMXu3eco+BdR0M8hnqD7zA5V0Jwh4614G60HE0WE1d1+qPk92
gYYvph5mPbiIUUs1d4ukxiZ1xTKNCoEXLFUrResNg/ULfFF/Y6oBBE7uQyayJYA6
NeE/3Oz//SQxNOaM//8SPKIzr21BnMjTvufl3uV5c2EegziBUn96AeurrbI07JFS
eD3FDxYSXs0VK/louiWiPUXlCpEPJYnhcpNyEXyauuAVPy68Oma4GwyN22dYuvJv
0w0K/nv9G1qM/VwAyKJ2o5lq3ilr4oDuyM9yqmQ9rxkJ/7m95Gtuiaj3vkBgi8SM
YWAeCX3E9RCx0QmKN7hroSZ7jvwBMrnl0MjOjq5DSl9xKM/hEg0cQf9HQG3T5ufd
KDBYGyM6Cjer3OwOHGPDVz/G9Cei6fVP0R9XdqBBG9vK2cL7eiPeX4ZV9XHme91K
IHNX/zB8QAj0BJ56nW1oM80aQTpFG19W0hTNZQCkojUsJZQ36lGmdrRTcdzPK/M3
BCFdX2vB7z25UO+Poa+75nKJLON/NSDO3nDCo6JdDeB2lyueyhymrCE6TEONFzVz
LXtJgoyIJl2uUR7dI/Qu6j3//fp2s9rog3gLuPQWdIBjedNi5iAWd842Hx+jJLx8
EO4N25Z9TtPbGGmkAc0W2vwQYMs4itcGZGq/WOFlU39XD1247zhUL54oqgyzzFDl
uFFPWp2csPdc7AonaxwOw/ehYPMWvcPUwRfVp5OtvtUQm3+5cLnvLu+c9PkUi6OQ
nNSyeSw2a9vxE27JObHOg4Nxoym5iVqEGNUmJzT+0D2FD68t5LiNfpmbrE7i70m9
PqwrjSXWBiGca0CWEu9Nfd2NR2Z86nhQPK/vK2SYKi22jryPuUd56LVcV3r9iOEB
ZTzcl5TUFUznVALNugCO39IdsIGLiHT3Im6gy1zePGTm33SYThcbZfMWtqyMg+wK
3BndPFJbgW47FGwimOw1NxWQPazXwI7+oR/mEsO+ZDhoqAOeGXdkCTBVDaGO4VtL
xjioobSxcE1oTk4ZpAbHU6z+uZZxWJYUqFS3WGsaaHe8zf2I/rSoC77+6JWmqQJE
STMVFiTJS//pgqPyEUvKXsUp5UwjZdAUAqgop2AsjimndDCvMeqFcDBPk4BUg3VA
6TH3c1VWXbmPO9I5G+vlkXuMQkf04GiGSWsJobFrqw26H1CtC1OtWvjtxXZFHF0L
fdNlBHz2yXOW6TX22ruxB7pl8tA1dmGynF7AjgRgD099J3swbGvdHVZjeSP7oCiC
bhetCZ+LH/Gh2SeV9TaFIkL5F9Ry7CQCuaUkNop4gweFygyrcI0Q8Xf4gYYDmbBF
tyaOdPrkuqTSXjb0AOllPbnneJxnqrag+wSwT2N1Lr9xZ8CakKFNm80isNuVbJQY
hhtBk7+TskrZvMjYdIwZlKBKGiT6rDAA0XWqBOu4PkhOyAsMqSMjNqiwQQOQaAEt
AqrUiewHLgIor3QCF8CvBa33pgOrdhdzqMCS2f9AB5uWOqcDO4NsVzQTU9NheIII
qpsUdRxJbtpj2efkAaXmaIwc73mwMrAu6BPtTs+TaLPs9Sl5iQlIrxENrlKO+sNn
eNqlPx2NVV5t4AW7pMdBgsBhJKnXWMdI+GcWTqeSKGZV9IET9wHr/P5zkai1pa4F
8TCBeBvgPAG3TDSWnQ5xiFXSOelP4dTnPwKxmPO0zmRxdP6ABUC9B4zrBE6zZeGs
etehQgYH1UEh8nmI+uXVch6vN72/KvlEN2aBccKKdUDPU/X16P8iRIs40Z0PuUst
3o6tbPpXotDZ1FdHwsZdAnwLZvqIKKm/u23HksUmE4flPJZn1RBZgjPKIO62Dqdj
7eXkCr0LxF9cWoyGCm/CHSb0EwuzbRsZ8KiIsyJIMb4VMQMMBexaYRFuyPM5/qpq
JFr5ATpyMbHD+Q9B4QqZrRLVZych4FpNVcPdt9x7lFKgPY8nfBXaFSwMwMuU35W9
wpO7U0yOZ47OB4zvahr0gSjfLkbHj+8VhR2ihyLMpkYx9rv38sCCS837atg5MA4W
uL0YB5k/0tklHi0JaHDC/YhQ/AwkNumqW80md/UQz4Oj6G6olhr2oQJVcoDXCwq4
Rb4WWCbhu2aLmLoyBI1Meo2DipFTPRy/JCHj0jnOmM4A+ilHqRE3QG7GrxIVoYTz
iBifb2WDNSXAOD1P8GdFT7HdcBs6jThcX6Vfu9nv71TuroNn81AGx64n4NVcsity
eW0YCmVXK9VnE+CvsNnnDXHdczIN2TjztHFnqInfo+cE0HVKKiYndAAEann10tCK
Q7o8y2je8g3Oaer7rcw7fO6QEHCiS7SyWBX1WRS/nawBpq/sxPTH2UVnAuhlCo8o
YPHhz1hOdhs2VaakDQC64UQ40unrP4ZuD2YxSd6lZFYn39Us2paOOusANX2rjUwL
AAZMhojx0ZR6YvxdTNV/1Cn5hWuFsL1toyw3U7CHV2d/0GQYvTUPGowU+w79wTgJ
Nl31CYdrR1YhRVw4rH6erIOmvNKZSe7xDsJoGefShNPQuwqSOJu30GjMpFhPoEgI
8fofkh1Ky7vJOHT5ACQzZuBnWCryBnl8V9i0jw5XAuEnBGKNnWlM6VD5KcKwnHvY
o+vlCw6D8rs7ks3bH58T9ghFBuY9DrNn5nUMjr+MZoBnvYAWEelby3YBdHCuP43k
8/IXQ7k/8Q7Q8sbqLUYlQPd2lMZ8oJrG3WwWIy7Ki/GnNutNei3fiKf+/y7O0TxZ
U/xrmuvXgV6JJBxv9lf8wMoKw+P4zYcwJZg1ri0CbqdwZOfPVQKft+Vm769YHfuQ
9BqwVJkMS0m5QQ09esn3tt8ygf8fGNhJVIafdu1qsWocAofgzUkths3lSztGMD1i
K4OrDjfg+hPCJTsfNyRb8vsUqFOhWrRrAC6AwPWDmHekE5+hi5GaIiogqJ2WxMTy
MSi63xH3clmUiS2vz5j5+48XMw5kyGKhxkiD8+fcgp/6OFsHfqI3db2nnBriUXov
Ra6K0UsCqnUZjNYTOsiMaw6JTGob+8A/Y9Vcr/W+4yIHqfgF2rn25fYwfRfU6MwY
7aBRGuGV2qwSbz70gopKn5Tqwjr9ycrjq4epiTDYI+ZY3OYVX999oAXAAWEOGfb2
2ADgH61ncVfMZKeW9gP6iCXtmEznZcblHE2pD2S6s+SPW/g+HuCedEI1DFO/9Dqm
vYi1oNuVAEXBef3R7KfRK2wYARLnOZ7WK+xVi9FeFA2nWQY6Y+cjrdPwYkJV0zhM
DJfKxXePDMfZd8l1rvpgyOLRjpVFTVWYvXUE1Lqstaf2V4q83iGtkvPxLaWcIW/W
dJuwWMBreq08CfDPS81O6T7rKynlBEFYbbHr8meSP4nr2DLf2xOG22xCDYGwgDHC
BNIS/ICn9Mj7rji+ilzr3HrGX/PF6ZnmmXafaJHPFGJeQED7QFg5VfyvTdrxBbkB
DX50SE7WLcwdrb0FVBp5IqoZkrsGIBEnkzKe+TEEA74IgyPEWNBZqywKRMhW8To+
jCMJCO/dxsP9VHmThANz2OqiK9AIUSLFmYucxSjP20fvzccsPr05GehT7+oINSnB
2IbVVT1KZzuXe3scrRjVpubtUreu/c3fMbAsbdhR/gRKZD9l7uq/A6vM0qL2ujL6
2VALQGcDuyfuXFigVnIOaKh47uL/5fSOraQwpOJNkRSZbUlq+eChBCYS+fPuhMKg
enOPBlGHopyMR33C//y0HtxV/me1wylujAUMiSwZj9PwJ7w+HBa4XJTNRWuc8Sl9
4GYuV/FI/34n/ZbAwZ17X3lqtcul2dyL5LbrSKT++iVmICFq6ix189zWaBkwSqJu
Mb72t2BVAZ2H5/L4sQDNzfHHdJq2gAsbaQhyFiFU5V0y8nt8me9/jMsI/AAnLiWd
V5MR/yZ4zWISrllEpNysk483OlVpKj0SOx1jj/dnLz6/4BB81GHxNvd3o84RGlL7
C8idaVNX1sn5c8MIuWWT9CjYwgHnAl4OZpcFBDcy+DnW30HlLeTsl0HO+ehsR15w
r/OCuQNTWg5+RJxJClhNziLXMaYrJi+KO/wiiao8GdluJiUlXj7y3U3jJTiqFCc1
p3EDCm32ARCV0thjjMkPuvQKJ8qQDN4Htybb487uvd9YFjmh4bT76r8KigTnRyTD
tQuneZt3mPz0sTGtTfMmQoGqD9DedvbmcqfpdzdxcRVX+HZVuGnp4yfSh2QgtgA7
vH1iHYBlPI19Sp23+nYvNdcstaJ+5AsG27pZgYas/ZzjPAjAQfQS/bVwhTpKBNkV
NGSbTzKrOcr/QRu7rTqAcNUa2zwgIWIOxDIF1tS0HOwCgBSzxtDFIAH+STGbiM02
3KRe1AvBx0m0lQM/azJ0S2D+5jayWiE562t8Cf0s/C18Cv5gCisAdrpfCIScLsVG
ICf1i+61cPz3zirX7SDu4tQTIqjFIPXQhy/Um9rxV6lEVaPg4dRVi1rAX+n77MKU
tKQ8XVpbEfh8t8zdVl9ghmnc4NRSFtal2ezHsI+WJjYUatlx6dBqsUyeVLaWONtH
iEpM3HVTV4IUHq3GbhGjIpOdQT9k5A7UEZn4CjKSZ1X31uUKOHkgfJMwjHoGBxYn
jpmemk+8o81JZFE4PRiPFTpXb6OMMiujvd7xlrg7pT36C8zus4gah9NyaOO8RdRx
enkULA5F4GIF+JC6eCFLADQeMSgoONmasj5i5+2Z6EdqCiqUMNuU+cA8IaeQbfJ9
rCSxagaS/gsYd+0VjT5TsbjmE1LvsFtunVUxiQvfH+Vj0VPveC0elFd6PlQRRHkn
7N6psl5d+ic45M1N0mHgxPzTuTJl5m2R1cp9lUR+jXMGBAodSOlprdmb2Y0kOfLB
72mpiH50GfOoT1vElQVg38XJzfsbCw+Ni+MQ1FQXamrd7+FKEl11Cs3tfRpXqniC
QQZRuRuCG7nXrfIuEVbhXhEKb/bcNTnHfQ87dZmsOyys398dPN+OMR2RPTfl7tTp
VgpiCggsK0S2jdugAvSC7QIx7aHekTsThfUQ/U4/iCxIMwH2hbm/EB/qR5TUOshm
lEWZ+OzWcy838xfvUyDsquUedqFqPVV0open1e9ngSD+oOTubsta3DinjEBuDMIe
6pa1n6o190XGk9KcanV8GH4Zk1ReUyNrV+139/y/jL4n+k6uJghrOSLyypmsB9KI
GOh74HkNaP1PUdxY/UehipdzUXvDenGxWQpiAOfcCrnaZvoCvaCPeKW8iRBcxueb
BIKTQJJXO1T+1WTIxaVe0x5T3Xki7ox4LdHVcJZXM754ZG2T19fEGspvz7V19dR9
ZSYfmNXtrgaGo/a9W3AU1mOnp7+z9zdTJ0TwLfJc+ePxmew1vGeeJaXUMOBO2pwg
qf+7jYI1dcUGOebSvcbl1MVG6CAivijRfbK8jBaqM8Yt05cnSfZ++OQiBAFfSbOU
l08l8GhcesdJnM2GD3m2bIYoKES1Zei9sPiXpAkOmCYkcjDSEPu71KFpp9qssS2v
WlVmWn9g1NEUnm1Kp0zWvlk72wqJEBrUswXb5dRn+92HarQKZycK9NlciniJqSR0
5f4Q1jRZHEQChM6daTrWRDFbPMk/PtBtFOaDfnkjz5J9qFM8y8pfYFcJLHJOBsgn
BQO8EAqeCUopOT3F85MwCe65at4huqLkLosCRWprRrOccT1BVfAKnewbaptqGxY1
Nuj1mLqxvzgTNi+X126Mt92VMhmssQ0g4jcjrNedHNlgDecCvgt6JheAewZ3FKQJ
gTuFsNftsX1UtORaGjumPqB5pT7uXoMb2ugMXq/LipLZKxF0nHhhBLYM9ubYLab7
IeUsoRgH8oZA23n05vw7nmltWBQH2ufEDyBCyaHdwsl/2rwgo9QzDL5gIA/JoHbs
Xoaap6ZI1lQrvPFL53t1VmQoL+L11f07UN85pnNaChNZ870DD/fHxiX39/WPw5LW
H2nXWYf1l7XmeYx1LjZMwTDXLtkqnW28ZBSWHDnZIIH85Wq4sVfz3cBcRFlhXHCP
GUCxXP29rWhTHY1bN7VlhgZdV4xMxzztLsIR7rN92QopdMwD08x/11ww6gsDpr3M
8dH7PNKVOu9B267JvUz7tTe/DIx7z+NoCcMt/aLQvNOaeWiLmM+/8bnmR1CQCfJO
CuoULwGcdtCzsR0yvHHwIDPBsg907g4NvR6mzOnzoHOCqC+9gBLaWq6Ci5Kj73s1
cgbYS4QtHBchs9nYBWRQN+Tr1hRrCxlTOChIhkSu5PygdnerxZ9/f8C8K4+AedOo
xIF3k5421cwBtHHjYIi1kCV9MOL1sbyL8+EWp4nXz4d4mB3E3i4u3vFFjKIgs9J8
9zpHkQR589P9xM53DQsZQ4GFKmkKY4eUmMCS+RUAABHWARHvafr5x4u6rUe8E1qg
KRmjqXzo0IcOxYSaXVtw8Nd9hQtcm6oB1lJtH8FHhptjTLThxWZW1UVl2ulcPl76
Ad1dYJWpK4IPe+OA1ZEGNT8BgsG1LdGmlG7sBTWSV1+ltXRHFZI+YkCV4xDn8iN8
Dn80/beC5BfyZ4T1cvGjnjcu1hI9unzXVpgPY/lr2w0aIGJEcF0yFD0/vRdbopzj
aUL6gOrkFlmbe2rvAESKHiXinFdHcOw0UR70BsMas8y4h7WBmj0HlBL0gFzvL1i+
NKE2DOYg9hHGO0S47FUxl12BkJirjKnFZV/x9/2NrIoebUyzYWIM8H+r3tVb3q4K
D+3MU0nH4VNNPRf5VT/3hQWLfKoy/YXx2naexkREf1SlbSabRGDAK7MRAa9kLnfC
4AKIxDxw7Tem4QWCNEqWwVFOcd5Ztj84CmmmZ8MIYISsLBufj4cCvd1sPQW+oZny
xMYZLRSdFf8Tzvk9Rjhcot1CDS9esgmShzj3bDFS6MAsaSAwLQRUk6VUQstifMcW
nuRHxep9KCjifkU4v+LS+eZSpNovvt9A8LRgu9+evTDl+bS1CT+mHbV4rp/jvY8o
bgBsOjbDY03wK3GEElk9Uqx30K5kVjlU3dV/7eNyKMqomaSE/KT4JgczrVCf6Gwq
QujSZvg89VvqiHT+YvvxsimDmEdImQ01p3NTdjI4rcbXPE1gyZSoDzrlBgtQl8uB
P+d2/Pmg38mjC3f4sAAvwH6BnqXt8h7rKHmSF8gl6IMPlprcG4nAi+cIZSxTftuA
e8+17At50qOzF80uGTdbGnCytZWJLMncDcaka8/wzv95C6YMBA3nl6eL7LLoIwxr
7lLagncjld4iKxu4G0guJkUijm0MuSJfZDnQYdKWCKDITTXOF9fxUELKTCGQgqhQ
PYOLSmj+S42L5sluhLfBR1OENsHjWhLKfA0dai2LZ5Zjy4le8kLxBHv+H/1yCwE7
6klw49JvVRdxL7MG1Te3vqQVCdKposY1Uz2yMR6umnAsMm7DJfOoP7iB94mfghJW
7be6asmUAJEvCrl2jsmz/K69kkKMEVf2P8lBztLhlXTFg669LmRG+GgJ3FZUym4D
MdyhAXOy0KwlOIZW07uLqpTHaf4NkAs0mFRUCsSbERVmBOY3N9bMPFEmBcIzT/ft
xdW1MwZJTYz9F3EsjUoNYKldbg1agSMLSFiE9379ww26U//1x+qvRFDuymiBvG0S
7/SV2zBRlmnEctzCsfjaxEVKcVf0BK15fHROwEq9Nz4Et1GyV8dI1w+S/MUgic0t
OZ4dwgsTtcv25/N4KR9spDxAE1UHoMCysvIABoZP93uX1ZtWilJXzhmnosoRUE4g
hJsHnF9CxOzkqW0j+l5AfllHfWICyDSJhWqrVrWeplTpBdVU9Q8WRKpf9Q1bdCtd
Btfow32XX7TujxzaZfFlnDQK2WkTJn44dBBsywZR/mVmn7kVZn+j+S9gE3Bdw+Af
cu94Jho7sBkb259lC1WM3rVzIPBXiszz6hHLw7FJsUr2/f1Ylti5XTY/gCaGlC2b
mJfjQXT0pzrXGx/IbYNPK8Jr9a3mXfABwMEidWftwDA5cdC79g3VHkxUq4qUhYjZ
i3PkMfsTp4226nqJIM8j+Qj+N6KQhGRraCzt8nfpK7M1ZQv8tah+nppaR8tR4fIW
uv47dLN29VUUkEx/5vzmHCsGDxuEILLWLD4er0KGb3+5xOyeWLISLsFBfXeSeww7
RLa8bz4FHGu13VjfFcKqLIyFSsmBXE9onJPox/fz0wTX0EFsubdN/alwq2Er/5yA
pLSJnYyyhG3aWuhZJFyxRZJV1BBnLYQ/UfUXig/B9Lze9HkMMkg8lw5ZqYF/f85S
4ssW5KKcwF2TxFoo/ZGvWNV+tx8EB2Bg9WdzwdVNqztZwbnAASmhd2f6ERWg+b81
WXdtFskpbcqo7kZt1LovCNUs3W3+1ojfnWPztIBnor1B2Js6tnY/x94PxjTSNEz0
zJgNkaUkVxIn8vukl8AuX+ZhrvbRyMkc/Y+MszQY5FzyVhMUNn6sl7NpaMPTVy2W
Nl2xOnumTKNTU1/Tfvyv1YHRODLoYA8SFkjMKBu+OjLahlbhxvOVy8zdpPYSfgo7
XhyxRkPEk20dTK5UqWdxvb4anRn8pn8eugSaPZriba6S3LdgX5bxjtHHnIJTnZPn
pIm5MFfo/k+X5Nc2p1SclnSjVM1S9ufxL6QgO72fb+c60Q0vwGfiJuIFij5POtln
PAUVJ1UhP3Uk6tUxp+oBZlGlpRi/MhzgU7iaWZVHLdGhQAvyBse70s+0Lh8q83+r
bWNSeIuiwqqo0FtptTANsymnnu5YguiGKktVa124ihep6TPlcWs/D+o2/SmYmvIG
+AOeoIUS4SsSeZQlPn+pYYz6T0cByYPDCUtOjIZTBqnUSC0LvvSf2rdQ5FG3FKo8
6d08KdlZ73BZUc0wIWPWCs6sMxpGm00VUZOCX8UOZUAw+0bOPTENvLdsbwNRFXd7
YK6eYAGZoIDCNG6Bc1TOqHzjQJfU10H571ALD2obg8BPijOGVTE50fyLR7POEdSW
fKCW0W5UHWcCXly1hnL5zSzM5NnBo53lmljlIsO5B0AqtOycn9mP/0DlsPtXxhLm
I6+2aMKfEFfg1/bL4bw4ioFuYDT+HUQXMY1U6jtOPexx7KqkZ3Ix30vI9OxdPKru
a8Y57AgQVooSIk24cHdUgjSv1f6dcewV5rB4fVtVdb/nWvGSj9QDSEdZ0yrztlXL
sXMLFyI2HbSj7jOJDyp+3FNsBhwnWQzAUfbW++XntrsmcUkn8SEa9HysNukhmR19
vtGkTd/BdbdEz0dlA42w23fhyIf+KODiYuUWmvVs9/O44lNnC7ASbtb/WR2y6azr
IP2sDYBhfCFvxc+wEbdLowXQsg6QOz8cNU2Ai6eREY/iRk/vEy8u73Lq80B2UtZM
yQHT920RK2eutFqEtt3CfziNEzGF1OMKvqdsAuDGBogHaAmOLT/nLBISNyeL8L6j
Bm5c7fvib+pid9/U1cW4aROO73yUSS1Pnq9V6vYB7Qz1xxHrC/B8BWTQCqYOk15o
/7amw0zQa3+DHHZncZUDHAv+jBQNGXkPwlpM9V/5A/74C0QQlf2WQ+7t9P0b6ReZ
hGL1M8M2SgEgAkAp6wgS9T76mM6zkZqbltdVa5/QENf+x1p/aZin0+RwER3FcL/4
eqb7jEKu29GqsUR67wEP12s/u13+JJUszVzQ8bk5LcwyS3HZGSqyLAKtz0PSBcIX
ZDaG6gGTcy2Z3DEkw2Iz0PdbQccgE0gKDMUWxtXOmhO7PehBrSjP1VTrLhxkJbp6
s0YISY9FHQjMB15srPA8l1WJbSifmKcxmkJNuFAdHcRmzfZ3dobOi0Z5XLnrQk4O
B2XSDqYhiCxD0zkOMNFJSCxlJa9t8F38RnyGgSVRKg4qpq52VylkjEEU+giwppt0
YVMAAvbhvO3D/x39J0gLhPnCixC1q8Oed5lvWRXISuPr+1YnDgf+2Edh00FiCUtf
SRvuM9r7ecGp4EIQ3yLFP6m+2G3Pth+spG6JThEZuFpKqHLhdHRN6fNrz5LSQfZz
RKmRpEDU0fDb5EQtA2FBd4wWKMZOTUH6adZQpGGmfk8bEwvEoxXqqKNIoEjkge2l
Yi2GMWNHPOg9aBZmFypryl28cWD9j0Ab8UfMVKkw7IhPsy6jb7TKOjbr0A9MG3ca
+sbUeOdZh7OzJC3smz8MmWbwu4875W+G1IQ7DFgaB54JYeSeMElATylNX3RmXf57
PMvypiGrhkJ1mJlNRmv0t9Rd5ZLYYd8dTZ7sES+eYqd/wk6twE2qhznLrMC7Wy96
bbUizdjnfV4KiQgxDzFs8LENp/H0AZmbzYW8Zqzl+kgG4oI/UdxwM4iVTubNOPZp
bkNO/sXPFdW/szXwyHx2oe8EVH0h1mLg1BpQ30FlcvFIwYsCSvcITmZe9NzQ4SmB
WEIPKH83wiDzHwpgK4pvyTkYYt95ZqAsWubv6Y18rnl1VsVk5rOLK5R+bIQSPdTq
QGMEXNdxZSh/XW8EvD9GQqVkJktyS4U48gZkUf3GLhJe0cN02NZIdcMK0H649u/g
KKy0D9XasAC8keRC9//2nAXlFkA9wWJAH3+4dmFD/pXrcWAHEcMp3XrClrWmf10k
acADA1hmZStQq8hXLSUHsOqYfSklKf0u7+CRy4giNwkZUqD6kDo74VV5a+NyueAE
GQpwgCBlQ4Z24VBIhp0Adlv7Tv44uQ3N3t03VXi2Nt0X5abFMHgW+X9uXAffAJSb
78jbgUwrk0Wq55wXdTbZTZ45cUUokqPHeRn5e5/vzfmiUoNjeFU5gJv1rUwqLFtp
HxQgD+LYPKyZGVk7dkl5RZoSCKBSbJ06q7UzjrZB1NMYTEl9NYCdN7YtpdbpU5JQ
lXwnM2P0d5aNukzNCSBkF/MAI3S+LnyQqqoRUxZVIq/jepek2StQuMMXAkSlJcJm
10sEmC2glyUSYqVcQ4d/XdQ9+uHFW2dDbA8pA1y3JQnCxPVbYEY4iVjMiUNnHpk/
vvF40qsLPtLs0xGze8UTFxS51dp2I2cv/hKlVvGHq3vylDiQSpMp8cxkoRylhcAD
0AMpcAoUjoIJotoswD/9wyJ8WQ7kRQO6XTunlIePMobbkkPc8hrpqf+EXKQyVDEJ
GDK3/7XQFFtj5m9IZH3/al3JpSD618UQPFJv+FYj22BQA83VQc3kave3vXtN5Mu1
UHxIRqWWrj+U0Ql2yJAXJESfcu8FlSIJQ+JlVB/jcybmt13yS1m8yPcXb2s7DBFp
8KLa8VYVB/4YdT9HdnU9yi1xCR7RdBBeJcyY3KknHLakWnZNiPAvYw6uLGq7bF99
oDNREy/9UGmcZ2p2XMD3aDH9zr1iJ8nIz2w8wFb0bqkQDJHrnIMDv59sCEnNcUqC
ANT5mOTKWwXAzJBAUScbBKifraTwqsBOkVyaeLjrJF8aYfsTLnMKXJ2EqhZzaA+N
peYhIum3WBgL9jT5b2s1huHRfeJjjvVEhqXHPoILfhhzIXD9GrgLurrm4z8UyH1V
fIlYpymqm7FdDoTX9hxNWpuYvREQqNpBRe1EFFXE6k47xu5SS8usFNSDKE6J76ju
0kXrlrLlKVsYt7aOApdzIH/sA2jL/NROKzxubP8cXiORVvQB3B9cO3d6e2AFnpGv
EfpIxeB0v48++YKYb9/MXpNGElbMtrwCzIkvbUx0uYKOwe7h1zQ5RSYLLa7mUf3+
6xOAuT9wW83+vmBgJeFVJuGy02T0QAJFd4SnBLkRWX00WeWS8rcHGGcRLaUQq4O3
PpZ31zS9qoK3iCdKLIJ8WoDLwXb0wLnCM7bWYfbraopHhSozwF5Y6w17jqfP0Zvc
5EfNfhkYT3evZmltLXS1NzB3DWSk3HuG4LNicpyH7Hn1dqO9JLcsUQtWHuUQzUuY
ExIiBHz+RUFzsjAPMVPus+lsFOvISb4YLZHVv3M7KmfxgtXnEhOKEw2IlWeAz04q
DMKoa1imOGbuHHQA7t8oTOah7kgyTZsC1CQ8VuJI2YQ0TOZs5qvO2qGQgek+5OKY
wYInLvlFU8XdwR1Rsan6xU5WdlvXh7nS5/k2zfAKBLNst0+sNPt3cSNAVtL6gGmt
NJUJxgdush+/6juKB15I7rtiIO/U8kp30UKEXCpdM9XYf9JkXaJFOUSN9wheTGDi
HLLuWvup8p7kKxibhF3Nk6lvrw8236gZarhc5+6WsiqSGu+2aK738fQIPqN48Pog
afPRZuxdObx2AvmETL4RDE3e3K3QrsVJVI/O7FnhwouaNR5nJVjPdnNtkDdbM+KR
GVxuW9DB43Bg2mFtZ9swcOSSGv8WcWUJckAT3J6+06QouFWYxTP/zHzaS9AQXKi2
l795BGTItgUSId9Y+UByWZNbPSnBtJQcdvEVFQ1qXHY5N6xDwF4B41ZCtWMdFD4a
99jOe2swg3jE1plbWa0xmzNUbdWo5fKhMN0c5+5WLf5GajXRvGM4/sSnC1kQT5v5
p+CW/43wGTeUtE67AkFM+Qn5wy5XTk+9Zqx/6s3QnkhknMq2BADl+ghAif4HnJ6/
nCr5J1Y2joLeYX9wXfPzR+/05hoS5NTLzV/TU9gKVQ9cT4YhyoYflopHtWYDfddo
9EoMBMQmBIXInKIQWcQC1fgImzH0ti4XJFiP0bNm5A2boFOnGUujbg+TEDD2/IU0
WSqW0h+Lf0jsusdwuU/JJzBkATO4UfQLn/1Cr/p60QTlLLZNG4oxFiI8wMEuP6co
+fCCwBK0Q7CetFYSun/aBfZDEztLKMZ2+2VSqcNH0rONDQ7GM67f8OsPp2/I79D5
xHJcBhDcpZ/6hqtl1LzXxYtlVzQMhgR17IeL3C4rDtHMfnPk7kubP7u/ZqFu9Jzx
silT7pbTbYWTAwcdIfw/fQehZtT1vB2Wz+jRbSHhQYFrOnDqBCiHAzqRXN+Q8r4s
735Tu67G4VIzJ33AWnWatGrlRJV8e0C+qUMbrWBoc5SlUOx8aZdazFsBltl1UQr9
J3GKNTaSFCg32GJqwovg1bafTerhR+f8grR9JC7mhD96XAXstlOhbriVtD9fr6LE
WvVMCKc6W1OJ9y0PAhmeL8Lo6WgP8wiJI5SsuHfchJkxU8LaaAhNdrQ2IQ5VwsWk
4BXl7qScMNt6uPrycgW4M/kObuMfO9jhDb6v6rjPVnoAGDb2hv4ckQa91yxxG/AL
nPGKocYzqW+X+4J9uAGcKymWZN++/XQdtDoC6xHtxVJCdWo7hWrlr+FHg5Z17Va2
EmKR34fZV8PfGsqfQparbBe96kF9yAQz1NbzAKPxXjJcX7uuJalJTOKun19e4SnZ
LU6ECncOLu+MvIxcsJD2NmQLDBSN84M1nlDDT1O/XP1aE009mL+9BlItvtx1bzSY
f177gHoGHS2QUUv0GcW0cgAM6jks/X2bEwvFWnh9UdwTvDaYxCK02AfhhvT6s9qX
lcjirBc/26CsDQy8fJyvgdfnC/LtIFP+rlnpkeJ5mwBcCGw05T7nSfqnSyPBMYUb
GQwSaliykjFoBCFSejl1GrTEjLgSQh/HMQGNOGTFiJlRnzgaltyJ4YAvsSGwze4R
hhASJxD0pEMadcDHGxeG9q9/Z3PQvXWdMIHQ5xVQ7cVm8CMc4BKXiSQ/WSQ90X1+
ab5uCId2SkwDE2gU2Mgm6fKZEICUX/wlihnMdXPjsuUiRCgNqS6V5ULokq7welC0
v7UWltidfjz1g8KnY736B8PB7NHGVQNootyMDZpG+lkVacDIX4Dl/JFffKMUVQUc
0JcikpguDT23hhNEGZY34if0fJCkY0rjEvvJrA3ppM+ZJ+roAYeUAHDXahN6Dv2X
7CxjANl6jViIR5L9TBK9yS8FlOv6QCcGWQLiiTSQlEfG0qolSPaF4L0s+8YYECT0
YbMKdmfqQWaQGxwEMRI8r/iS9petRztcqVh+n8xYX+/FzejvDrDNsE6ZarYVuUKs
8Tzdf8n8dcHyIIDfAjQsI/yN93t5+3JAnAwK1UbnyAIjl01PSrMBxGKqpXKWNMxE
veRyJrTkUSK5LH0UlMtt4e1gp7C0B72EfhX+WuXNpzqZ53uBl+0Pi5Ck+uaxXGZg
DtHbyWYIWOfAUnsG4qzOxdnustShxj02dd8VLzsjxpSlei18gQsCmNvRKjITyy4T
+nenG1OMc8PwfQ+w+7Eh5iqoQalWJUqIpUXNupJYTcmGfdq4bZWa3eRJ/rkq8dhO
fH8H41a2yv3UA6fCgQOTdTAIHR5yW/2o6+VcForQ+y+tOrNiaiibK/kykaQvC8NB
cDnpmncW5meZzd6uWbiJ4eGevQsjJsezSZFTEUtmtKEwdrvjzoVLPYxQ97AITDV2
hyHsG4ZDqaz9jq+TZD1OqJo56BqUNM9w8upKzdDiPfEQoAJuk2wFEO4C231TLYAQ
pUf0S75/svuvbtY8GLAh0oakkNrjGohS9AC5HWLf6sGlPTWLFmoSmyPpkW5PUA6E
eIz51PZPZLqK/ri6t9RpsaN8cyGCOn/el0WC6HdiEx8013QwYwGtwrvrbb445H0a
6MOWW6p1qJhq+keHZdPW6PGixHJ6AXWCiHm/ewV9+YV6P9HrDEiUWcf73N7hqlwg
sRSji3AVhbljuW9WTKSBv60lB1FSNHk/n1dqhERO7v/QYF9N41x8gsK8FbXO1qDo
NZM91eBMRy6S5hdhhoVuBKEpMFIa+pgLRTkMW1EkHNZmrYZ/ZfSb30RPVpg3jPpe
j+IBUwO6dWvFgGvd7DdtJd8UbEmaVjEgLprSlR9MhcwHuepr1tufrXqyaQ3r/JIX
A2ZFHumo6EHX21eRvoigTWZxctLTazSS1hO8eUBagms2cQ10sQADKfAanVfEDq26
G8aXSwGCT+uwR4EAXlGEwE4KOPR7LXaUU7ShbF7/e6TKiWhSpNITVHRjB0NOEl0o
wdSmDUhdwcH0+W8D4QEYxHbGbpoHyzHiFQiFOptxNQug+zVtQCk/Jsa7pKzEJ3+/
ErPZ3KBJL1QhUszFEoodd7ur7Kh6wmQsdZ5Zz8fqSoNHXUmA2jfKodb1Ew9rmv+P
tK8/riC/3HPDVUeI1J2yQXTHXeK6HnibPkrUtV27FhvItigny/cnmW+/SP9nxYO5
VxwH+AZ8reae6KeGsHrliL7ziIunhHuYUlpvr0N5cOBjZYLsMJhdgq5POdVqhccz
1pqeWOjalOHaqjvM9uSMqZzxHRzhkm/A5yw3sWS3x23ZGAg2Ors5+NFHZVXVGqwC
Y2In39v7HAh8yrRx2s8QZxH/Ws5YD/1d1wVm077Ij9zBijDt3EUGRpWoRlcxyIhN
aVIGgyxYTWdHPZLiaj6WAztb62njAL+iX9JbqbcLod+9lmjAypsdc9u9oPbxglrJ
lCdkDgBG312wG11j7wJw0QfuMuXP1SrhOLRKjkwCOX+nbdsOt1eNNexZnn2iZ4Vf
dyYD3DltRR6TLAtBon8Gt45LrjEE+zV9S12wncmvqr21EQYzyRXZ5W8UcZ0SvkB8
DcoLliQN3arCVh4gPdWhkOtJvaHrkOu50Qbo17f8XoxaLHK0FfDa24wThzQ8slAO
U7+Yojb9HmkFpWOsi/EF/tcBz3h5zDzpUwpadVOV3B2YXzEFOI3Y3vx0rxc+dUJi
ZcVLarePhhhceMsN8PspyJ3WvHF1Ofaf3vw2GJJdPMkbJZ6x1oSKSI1vWzeLrFom
y4jlGtJ7ZSU9A+keuixthR137vP8R1SW1lHkJJL9onciy0/T4duI9HeBwve9NzZT
moq+XLeUwi7eVKes4PksRJcwLB8QFSZQuqADDnBXOgpesR3qDc04xo1nhn3RRd5m
u0zGhDFW0GT+zyK6fORqiqFqlfRKcx+7ACdecDd8tXfiwQdOs2bb4I5Hot44oTBQ
TMWPqtNu4wRRoFYowsh1KBXOOt5qc8KYCDdIsU4pibWrdTf9zenrzH1AAmx31Yut
JIL/p2YosbQRX/F/4Q4Si8d1dOkHA1Ow1zypxT5v7tkP0K8EumiXRsF40H5+tUGX
bTvaZfDPzeZ3B4kO77w8eNGlMqvSte4kR64wtPZXu2lo9wHn4Cng49kNxDI3dZEe
Dl1hfdlYUGeAhldOdAwDWl6lgpavaCa9ucDXRG6S+hYjKDEP9kPNc245HrEoxzLU
ggmK0fdqSG7edmiitBdcVf9z/u8nSzzOGfqP0S9atkC/S/FcsRAOtFgOb5mXNuLs
M6XGzZwHLHwhiW1JJB0D6dzNaf1Wu0JcX2UKNLXhKyxHKKnNNsflxH1E5Hu35NHc
C+udrWd8C4sl8mwu8cAMfE9GlF+rjWcj6uXdn9C6jZeGusQCqgBrR6tb6sq5HVaO
8iQYUjD0IDe7eeKL48Sm7Y2WKZlIMdbN5dsBDez2PYm10XhtxFAvZcj1ZXd+xsu3
4iJiV79iVubA8j4PLCdQth3YlCZB3lz/TP6QmLq46tsLxFOdw9dxdqFATlnJcwPQ
h6rzrfaGI5R0X8pVDF3ovy1z0lOL2Mysmt6uONEJo/lhgzO/hIkUuOxuWAUBFhGn
zqpsRgBdKxXQAAYuAW2mVW709KTkAlI9jOc5dD3GxdNr/ROe0MU3XZ91E+4vzisM
M9ttkaiE0Jh6EXUh2qP1u8XOvEVZxoi16JOUEJ73yYUJfGIcVknXp7S7+Vc+UtGF
hlcP67MENvPhkMyfdrbzYj3JU9Y3c3v/00uW+dh+KxKsVl4+9/5sLIb9j2rzrVFO
cNW7Mk+JkmnAjCIk6YZiSoUhXbZFsH4mkA/VT+TCMa2PpmXyiNLndoNVWLcWxscl
tfENpko8H9ry0RetRuiyLSBUWmJse8zZgYogTIgAXK8rPaCi0WzkQe1TZtvNWndd
oiH3OpNWOmAeCtS4RLgT5HV26WXSHR1xOw3Qy60DkV6OkOoj1gocmQyY3ny9LcDG
xhTmww35UL47uaUU1BDSIdrBxgMsNU91olZnaD9oPn/H17VUsMBJu3JfaS96/n7L
NgcAp31TtNwhKobD8tDIkDwD/dxzDPNKThahM5A3aFV52B9hDQvCRkdmuYs/9368
uvU5sj4QZCNFhe2wUMYlyefEYY+Sl40yYDypAy09wApvVaGaV84Lea2cgAxh2QBH
MR6+H/ECEZqHCmiwCf7WOeVmDqOA8qqphHsSa/JhoxdeIdqtz+sXArH59W3NIWBD
PdvBue0yvaW15Vy7K2A0jzdPpGMg03ezeHbfbYGyKaWOCBF6APEFcE8y0VvkCAKZ
r6lCz9T+OvSd5Wt4fasAz1D6bcDxpHpkVPkVf4/yOlOmZWNWJO99iapI3gegm/B2
6dPhZAJzU5q3FBpoLsBjF7FDota3vqYgqy28KVjQ+b3oQHCC8NPcCIOLGR9pHNeP
DE5q7VehI73byWVha4jLYRnKH+x/UjEthYnfnyowwbvRlwll6i+V0Q4j0XNd1Ofr
nxxECL6fw5ESEJ+xP+Y/JLY9JXczuquiDkL3sjLZBC4qhJ610LnRxCs5pyzOT6v5
NyL+sLzXZEZ5SViLB4pOxyyl8DN+jG7ztf5+RmuyCY1WOHJecbEeh5XQCTbgf4lp
hqy/DWjMLUk5MRqBrejznsbR+m+a8gJoi9sANQ1NPGEQcjcRZuDg2Zz297MXHtvO
T5g0m3WFFLLPxOpNqpwJxGp/glMXjj+8yn92zoxT0Yhyele3eTnwrhyQ27mb0bCk
MVCq3pWMhp2TSMVodwTa3yIvdjqfd8oNjpZEMs/V2qWdz4n4mXuoZhvVhIIrwFT0
OggRGFEQkZmUMX+dWdE3dm8i34yxiDh3Z8bvKvyQqQ7zEjVaKG4nL4scZ04L1rLn
jJzoCRWDQjhZlatlRmDCPO2KoOH39nJj59B2uAIvsk51zYmlT9Iv9iBMSndYvkos
Sm2BMhdUgLCptwOqPZq4vz056yTkwJ8HZxH7a0s97JroSWaOuLH3cd1WK2oCAenU
g0WGrVGp1RRNFROYOvMKtFsts9PchlXh2458n2m7o23Ir4XFa1fvkcGi/lRHERTN
JKNIw5zG1PF1Jf7EXKMRbbxFbbu2tclmizD3VygwNE11X4qR6+pfOdq46W8Nv+L0
O2RpOpCz+aX5ZiSqDMwEhyLSNO5PuU7gqcR/VrrI1vjLWpVffSSHvxyBo8B+HhIQ
00006xZfi8xxdX3S1vOisUobDyS72BAuPbIj6ZDdHawZqO8aztUH18vGhputCmZZ
w7RA9e/n64/ag/5mA/B1nbS9f8C/yk/PxgUrkIPhYqUclb7fuqaTX/Y15BalcLno
Xnk94xK0Z0BZPvlKfaQqNoM5Yo5tNgcek19O9E2Qg/nQxAmjMPQY5X6HjtOzo3vl
13jHatRnCdvdX4fIgGihDVRT3o5FL/+VkAS/+ZxuJ9ddAUPTgJMfpe93KibmLxVX
179sP3+rN9tB9yQHMsIbBtIRSR/JSkczIe0NDlGrG04dlH1CHHI8Rd5/9XMu604z
cdsRgAryQ3ta/88r6gnfMc7L1Mek0TyhPfVGqoTVrr5HKWvSlYQRqDavG133N8d4
yEZLJxniMIwgRR6dIfzWT1ubjVaYZbdq63r2Cf6fedNDhjPZxaX44fkKUIfRggA0
yr1G9v13TjnNd/hmtsTGgUfgO/TCrqvGaDrTBkF5wFyiitG3JwwPppUIcYVKyKZE
xP8Kk7NWq7/hdJ/6FmC8CgbxfXyVkXXs+Ib3PTYotLxxJO/1x9eY+l8NOyEdUhwd
q80ixBCC809oDlL9SD1P67Hvnke3G/AquBObX7DVwiG8N25qCEdzTuGZfVN4lSeK
8at/BFgAfZohTJ9cykok67qBjEBO6pq+1nfQWov68lBvQRpfwNyeXRjYkWpw+trB
i2igWfU5cY7aCk6meOwBD5GTL5koq3DpFooycMRFSGVjfd8y4MZ+engVOl4Wz/TU
jC4qeONWSJzY2vHgPwyMroQoXMn8Rd8T86/OL3XIf4B10dpx/GPZ5+Hj9MAX74sT
PtcJ98S78YoUpG7ZPkgVgJqeYwkCaoTnpBVtpR2R/m+uleGWmxXoMsnDj6A78crq
5pVmULgdQR9G/R01+CogRwVsrmN2SfRy9f+JLZ2TAHLzu0tM3NxDrSlPgM88PGCM
Hj1T9sweX4xzrKCkyhDujGDREMUht4TI/o/zQ4vRJtkBGtByFXN5YAcqr6gd0kA/
CTDXR3ecBvks/bEo3Ht+HjXvMGgqlkKXXD8p9j/AjFUZBR5Sp41o8XpyEXmlatlK
/NDdezY1T8IztsoPkli04NsRPuPtw0jy3t+JieweoVxAoyBGCHVEE615Cz4s1h77
m8MKnU/IDlIWhJBURiR+s0TmkaWeSki2IKW4BOK42Cxuty6btgy7BPPdM5GO31tp
ds2CaoCLxMyra9f8QW3JBT0HvByCRzynKuGfZxwblIQgCDLFl/JpCdgwKmWyoyV3
sR6WofOkdXwNv6b25Rj5nzZkojJ2LLiqK5CmqdFSm6qi/lrQDlHTX/Qgk1iuEWUt
dyfLzMFNRnN9y8tzr7rmMGnYyio8G7xc1j3IJya0vWtXQSYdxKIc5BiII1JEqngI
UhlLBaXOl53/sTinSiz8f1qlEDjB3mpRY5ESkqtqiWR/RggE5UklZgrcaHpbUilP
5xB4rVJQ1VLVBc2nMkqVtfLc13M3rfOjfODxP0Sm/YdfnmYm3gDf0qMXS3tVXwAC
/9+sapYopMrmz7zw2mV03AkYj07tAsh/2PMqVr9Fj+zzGCKryRhw+NMamB7VImbU
FtM2trJVtUxXIO17gV/aesOArO6R6KpJo/7mYEpnFWtW8KWu0b3P2O/Q28kioBw2
TK3yXDCmwQhf3gdbHVwbqrgWcnGhhOiqPbkVFgu14YvrmTIYFFYwCCwmStlvzOw8
Tlo916x9X1/MWc2N6v04E4imcG5pypyqS3vC4TAae0wYWfekwrDzqTWs1SD1RJzr
5SZc58Vcuydeotg2kqmARRxXgkY7VPXhKcun0xi5bb0qQPcmk3Hg23QX4D8aQwNL
3bibWyqaUxwLrIdFYyE2dXkXXEtqY6/+TuIqlOSU+751r1C3FXTxBvQajILZsWPE
k6zEk75N5PYRSIqrQO6K803DKuggo+2JcJPjmRg0z+BGQgDChubEiJMmh9iK5UaP
DLNqTdyTiQexuVkH+IuoUohQjeU/tU4+r0jcGKwGAf5KBVE3LoEia1azRLOEgTiK
KcBN7SiR2I+cLmqIsHhzspeG1nVh+MvDgJQyKPFjVRdlxleBRjl9Leaakq9Jb9tt
V3seBLS0JBQHVeQo4AeuE0lIWjx2qXmT7fL4z7uBjD/RcrKN6+/7i1Wz04iq6aZt
deFjohdhTmd49WyalnzomDZKqeXGjQq84iRuL18hWUQHc5s2HhK6AC7BboMJTfHw
v3/WGnB2wePRyO/zyOL44RFhqjXiIZBLgyUgDzOjmH8PJUXDtsqX8O89RPWm7Cbz
z/rSh+G7C/q4u0dLKiQDunsqU0h3uKSRumZCmyVT9qx4/bNCPGIReOzDW/gdLVNl
crdwrZzQcyJ+EJw0FbgnVm5tei87X95isEQRWHrBHpW9STJxc6eq9QTj7v87EiAF
DjMmjT/mMItSf/sirNuRIUCzBlbQun7TrfXuNclUog676Z87z9vYkfUyN9dtRqfZ
3OGKgF8DeWY56I4A9WbudvxfB4rQ3i8f/StnxgEOw6DGD8870oeaQgVLpwQBt7BF
slHKzTbr1KXPDM+rsFHXEzGMDmwG4oc4mIp4XeRIS1uMvo4EatE5MHXDWVnPP6/g
NkfC94ysf/G48GcYbWhbpRhC2IhXBRQ2hqTw8MJKtmAyEupUoX+V7eG3sJSdRfKX
HF/PNkFT/9jHeuk3QP9+kDtxTVhU8bQIxLkE6hHAWN7nzRIxX2eeun3KBkTFa6o7
o2po7JZcQGG0UHo6Ja2HNIvWIoqyBn+DOLLdqeM0IAfZuN5d5Pxs630b985MHKfE
/sDSeSCioGwBD2WVWD/mKd6z0Xcy+r1k621KKRw0nqgn6FvFF2J2VXgDRbTw8UMY
3cBzDjMfEWk5u6LbJbr4KpPlHNlFIv6HblTvKWP22Qc3s50yWOo+jKWQeb2qCydx
HEuX0EytuIx1FeGmwl8FfrTcsquqDJo1uuCYKC+9c8vWPt3O51zqLNyWXskjUfrQ
lGxg0HwyfuSKHKcBPnGoyA7sOlkt5hQFQ1HFCafkCDZTZ8XklBlRFxOdTdlj/FL4
tnx3sBDeR9WUtOQajGquUMPxMZf4PWO08LAgKoYwIWzatmYGQcrpk7O1a3uD8pdP
vg1qshOtdvn2BMMsgBepkNv+5sTR09Q8mVUnwrYLg1i6hTkgtk3G/xjhi2cRQtK3
WwEHAjHv97SraFDoKFVh/rNqD0EvtRzJitqCWK/uNPOGpkZDV05++UCYZTLlDD4T
Eu0TVnUQASte+DV5k4D9Hebn9uvUXmGkoA023i6HZO39oe9i/R2nwWI5LBd1tUop
KjDPL6Fzwbmzgv6YedFsLoRsuuVB7Hmq7hOdYfDg3GYiLTT51kqW/WD4hHK+UBeZ
BKJYlUpGCAOpUlUko/AxEugbjJGD45QKGH7ylLDXfVGTRUIc85o4xQ80CRo8k1KS
zT8Xgz2YnF88F2Qc4usDOajNYNJQzXlRDbUhGQv1max7fatvXp89kMCrhVetYERH
8EgQM1rVE0DuGSSLzXQDUR9IVJOuyORpXpb5Ww9uOkEZBcxkju6MPljCCRNZfCU1
Y1dqx5ZkqfFJIfBZDlNJAbWwOih0klA0wjSj6epEXmnN+wsUcALvBe6U9J6vxnVG
4sKfikEg3c6q6gonKZiCTycjocnj4S85im+tTaKteHm6K9z8qRslfZ854PDHWwKi
49Bn5wMU/7+3zVrflCip66Q2zqDlShTgFAm7JlLWEEn7oqxdKm3eZgGpbdPzKGk8
Rrbhf6q6sLY2e6W1xs7XxJ/nHZUfpmULBWPZ3HBPqPA2iUm4uCU129bg0X8JcRt0
i+U+FxIOr/RsS3Z61DZGnFnT2pwwuoUVeuXTWGNbUOKe/FguWbQ8TpuG6fs7DFfC
UxsyHlw6cYHpXeBk7tSZ4Fgd/iE/47paTVOtVUMCCpieqve5JqXSa/OO7G0OBHqv
4jbag6HgSteVPo84dWHSBSYhDnGJhhED93wPEA+Q2cD1PoQetIQFi/qa+u24yoGh
hMGj/Ez9oUsWTPLv8bm39jSiF7kgYap1lemuJvsvxD2CZKQluIxeXVFUZ8yFCU3d
AjxvA6BlGUFNlw9faBhd7f/GyvYf7KHKNsD0qNRSi7sEn6P6xP32jVWd4NO21E8U
t9/1W6GMjmacXGLZVEM77iU5T1PJ/9oLSr8ADjQSBIViBmkBxp0baKjitOag/qji
kvLwJat36igNhVdCoEABGdQ7ypoHFq61goVoerziilsY0WXiv0yBwvdvrAfUTXzz
88YNhJ03TIi403WoAv4ECn5XM9vhVXam6rlIGJS8s/iTVCXjGEbV1KWC9dVypqQ8
ejjik7lJmh5s3+FJZxWUgjKQ6j8KXqU2cR7Nd+l6Tj850mJbBpdBnL+6sqwMO+zC
/bmVKWOW/R41tQqjqBG24OWPYTYKc1CLjco3rzY/vcCXFdptJqhe3SQ4uAQ2BhZS
tElJdi3LkxSYkvmEZwQvtZiLmuccSIpOAIDWy0KXXc1vXojiCvwY66H2fWmmrYYu
1Mhb15Rt2Dj1LhnhT+OwD3H2a2Hc8W5DaZ/nW+l8Rxvza2V5Y5nm+ZpVWQulzyeW
VjMhBR7g67rmnS4d91SVFct82e6Qi96DObfidhhyP2rDB1okE/JErgoFEO62wPi0
LP6fraVgjdT3mlHfTjW0BE8WKvC6JLi9C7Wty7sndB58kIP9uK8bvvbdb2qKwlpJ
etGInOj7B4c+gY6PsUuFvJvkw0WFlFdNkckmqnTLPjVPIdZ6u0kxQrNFH2eBPeVW
ZFTbinli99LpNo+wIDs+am6qmRrOfLCLCpu+tviKAE68vSSVI5+LmXg8vJZn3xGp
uANF1VSMfCz39RUvHkQ05cdfuq0up595Y5/NQmMcdmOT/tDUc0oQM4XaKHT3my+9
gYP53YDJZFzIG7TU8Wz9u0XO4+cEF7ddKetP0+TrvFQZBfG0n8ekVw9HJC3NyANc
PKwVqVyCyOzvI3VRpUxEhgguLo7eCm9ibP3sWJSzntt9f81azK6iMmLkcdivTxNi
jb/2ujK9PuR3FfsdAk0vfPy5Z2PiV74LxZZrcmrXVcMaVtY1SL6Gqo/bNPZCHl4b
ySMkKxcobXhvXdbZly7gKvP3fPj1VAUjS83ez84zEONiy4bQdxOX2c2vDvZ4Smc8
4sYY7KuYPIZ+JVBYZh/WEzxDEm8BFq3khhCf/fhE4YwZqUWjiQlEEoxuB/5XqMKU
DPo+OH/l0sblcz4js8QQXgYk5YWBPV2ykOQkKeTsuWbZ0BxGyJd+ZbcZru/tEP2h
lqMrZJq3JduMcRHOS2ok+DH6QrqQLovQ020WOm1FQMK7lsh8QQ2hFAQpA+95/u+X
9mjen5rGXzg3qT+kUGGzLC2aHR91vl6KBVWBlnamOq0oqCgtnsleqhtsYo2xp1/e
J4vclbB2C6njx8RLtjpEzy4uG3IhzTfWKa2Dm3lkXX5PtPKbwHSxtTjawmlJNBKX
lwbbjbvrDRw66khucGLqEV40njaGimjg54fUzTvnyAUgPx57jFKCLXo4wv/l3jWm
Bu9YcFodl26ngVz933vB46lIESvJXW81pzcUnN0RDYadeh+1lbmeuFePYFGLlqLa
e44fzVSwdw8PfYg3HRhOLSgqKKGItd9S4GerPKVOXssmvEgLyBsVeqqbopaAd/Dc
Mh5+O0dclkiNL7I8frWIH9yG7UyUQIpfo4tXROoyBWYHAm8EqDw4nZDLuHF/f6kV
RhqcEcRZt+JKUTNuLtcweR8Nozq36JNhV28L/woiHgjvrYuBDZqZwN3cVueLmdVT
AvolQiSUQa94BOWr7heM95geOoyZj8Wbq5BLmYpnFEsFvd49D8z97zQ7STL6xyxD
8L+iKK9CZG/L3CuiNYZBpNsoG4T2pBYjD/Qt9J5TPmJB0qUNJm55+zjh0W37+bwd
Swu8Nu48bzPVwC/DZAAFIoHZWgpjb5ctSdEFpHRIn0j5fGq/dsK7COugnH3feOoL
KSNFtXIzoDXIOeQ+BR4Vce/enL6L60i7uUsFaW3fgSuXm1hrf5wLCgzRyR0v8vKU
85uoTxwSOKZw6Nivoe8jjjEXmNDtkXOGXvJ+X/eeyjBDYhTw4zhkS/jUigRJAxyl
ZVrvmEbUxXmXHQNVayni3Hndgkl30tZ0TZWVIqG9wV5aViHOAshA3WxvXoCz2qIY
7+hqbosu00knrSARz+6m/O3+WnegtjHwTOTtwgxyl9S8I+g1OJ+0RLl/ncPz8TXH
qU3rmPx7A8LqW09PHgdwkvvW0zikckHFoggCStL5yfwOTcMyAMITxrCI/hq1+uMn
ib1ba99v+yQoGzOnSv7JQm+spNEGGgGK+s8PPLSsQha6Il+9MEJBfTGqhENrzzhO
VFtvl7z1tBDpKyIf/ConRc/LZuITSSwea0B0Ruop1UWrVV608oPe4mz4z1xvlVhy
+eITLX84LwOiXV2F6JpyqlgnFl9io2dOffS8nubmgyuq9fl1zEgVe98oCV8tVmf3
QHpAyTeht78Qs3FGVHVUc97NjUjEdtfHYo18exWdIvyb1wwNU08TsLDY+a5n3Hw7
y8mhOannTHzOZQgmIO4+3OjCzIHhLSfSp1kGOCXSODdudTh6MKccPe9c7dY6CakW
vzw1Qf+XG1mYWQl/PgJvLOWklnQhmH26WEpCvKpBYZhGDS1ZWatDxV5AIm97PI+P
60xxyP5/VrQ49xHRhfSQsRjyadKPxgT6PzQZ8pFpD0y+V3/cSaA4Fe6vV9vP+63x
s0QOGAitkR3xo1zAALwZc7YcPjSL8ZZ1rwi5sB+hsn6YPdhmFA1xvhBJU7AorOVZ
vn+ffeogEG9xrCQa+qRqrbJ9PTBCrkfDzDoZq4OOUmG72G4SnOvzGRO26Jr/xyqG
AnK/JRHA9CAIQHJlrHm9cUYRRWQeGT8nrfnMXY0hRD8QReys12MoTx3tFEnw2reg
kQO2YFFNdlwoIqiEFM3QbkNxibseg7xouZwHjuu79OuARSdrhKG9wF0Cp3HO6+Y0
CMovozpxUxIvQciryu+jFkx2al8hbDY4PMQFPfILDyyRBLmuLDhE8fH4bmHizUhN
7smqsLRJ6ooVCwkXKHRZZzCbhkjSSLMncK8eRSQHB76yRtfNng4bedqZmnTXS6mR
+BkqwuN/UUVqlcGH4vbi482RJx6PSSc4WOV2DFRbKLfmFN2QA21ErNPZ2R5ipBK7
tAtPlDFkX5aNBM6EcckJtirdKRWGAxrwb5afaxLVWS0DC28D+nWR+2dyFjz+aGKV
bIO3LgqwMFKaWUKV5IhuThSTLbHOgjMTABo7MgsLM9TWAESRZRj5bsm87v88sH8c
uxKYtXC4PcwZcOXexwMitLbNi9GB1C7LYVUyQ9MxPQQnPxHT0RWyKMwxiY9LXXuz
Qey7tLtpZacTsQaOftI8+d3iVFtrF3xS+MqIlQoKoSq9mU9EOtTcjrClwvDYW3ap
WmWtvCS8Sj831ap5McAV8xajqYZURg94IJ/djGeuAX6Wa7+wYQtqPPXl9DnvTJgZ
CyuO00skRguLkisqlugd9p3S9v9xCqdus/idjGrPg7dUd8v86iCXqFf09cwgo3cX
sEz1LT2OVFVuzqvAJxBu856C0HHoZIQrbRUcG9+zf55d3Xji+Fc1REWEnv4iIo34
moOZxDhbyqN4u5dQu0LLaZxQMY9xyJM5e1Ph/piwIjE7wAPYyYmTqc3hLgLmpqWA
Pi+1NikP3oEeK/Ucgy+QoOK6lDV3b/y6efZ4rIMKiRqK+F7sjX0kZ/NwhLHrhhZ0
U88a6MMwcIqkYkBgMozlRiCGZDo9XQQBkJBQ3GIXnHY7B27/xNrMzzRDBMoJpB9f
5a37aG5bYVWrbry7bmYO2IwHTf+lC/BpQvM/8dUTlmPalk8mFl59OyN+haxRKAg/
QxnzL74KWeUdX7NtjI8lBi3XoX5QWUao86MvxkngR6YvOp/5yQyqbuSUlG+F23wD
k6FvBcACNILZNRabDdWUhotAFdB+euOgq4cHuQrRy9TOFeTgNA4dNV+TZKFMzEPW
ShyfjnUAbGA0qNdR7SSZk6P+s2oYRYLPk0XOBvY6Qk/bwcOKyDOvGmtTkSk2QUvV
PTKp2kM1GtVtQL3HRwey58dUnmA/tPYE+QgimgUpaE3D+7xewOPJIZWgk7unQYZH
OCXF5stTPYzHoHMxSWqTuIdSpkmNT62Mppo+FbYAMhAAXYaJs7YYcJe1m9STvm2w
gE+niDCLucyI8vn+tZnwOCbR5GvwwiDPFf27M3vKaqMbnak9FnbgnzFcVCn1koyD
5qpfRpZ9Bek5AwFPhBiLGHpC/C66BG9YZVQcHk7MkpwHRYA6ZEG1isdhG/g+NxS5
ah1dPedEtBH+kXjxJ4n4jSeuRO4f4eh5FURlp+gNI1x1J0QqxmHHBZChiERfrzDR
7r3MUb5WMapqvMH0hTjpq7k4piGqVqD/wv7vH0YiaiJ2bux620yWiGEGGSbOCFuz
6EQxh3kuZSBLRhoeJ1/K2HTa/VUWX0i2dEFqRJldBqEydnNUskU4E0RwrZTREBkb
abad8yetdhhyl7eEbh9/eZceGaY+PRHoG6QPqhFoXzRdSknDho8nTS+6LSFEoILv
T9okB7+W+ONX/heRYnUbZoHjPLfUj98zctskyljW7aNSdJI+tyfTRx5dXdGtSkue
v1wSpLTJb9XkA6lh1KziSdA5vYvX6r37ivheglUjswZhSgZz5qRtTMLBmSCvkj8B
h2vRMY6razgooQ81ZUYz35jP8be7AdUGEvJFlX1lgE6fKuTdUXz6YCutjhgIU7Bs
OHpxIrLg2VYvJCwOBVV3SkZrq2v/DxHqady4V7WQk8WPRJv9PksOKN/TlXaVGBsQ
6Wjn3PHdZPuHPttJ5a6DHQwb7PLd/lSjWFXZPzwQjb1CZtiyRYR0/mX0wNgiM8Fo
Lh5sNyYhzuMS4ycNRzXjX4bUuAVTOJY8OaUyYUHA8kLONFUSknWqrPUZKG/Kxw6X
Q6/R/7Fg7tyz9/C0l/UemUvlceY3ZZUw3kTYW4tnpRPrQcCJUl1+EvGbzWsNNds/
N7OO2Amxka5LyBtcmCk8RxQGErdsILkyap5kaCY8Z05ATNlegqDXuY9sJ5eWGgdx
BkiXmmyOAAy/Xz8EBGaG6V8JUDXCTUbz6PObK30PYRw08B2nyeXU4oED/s/Fmc+n
sOMV2UIshO2nQTkXHD0LqzqtVno1GINS+kR+Qyao61At3i1Ht6sFAgX6fMRkbCgb
8cFiMBqAR7ddMc8GjlopO94dHnp3RZvb9O/a7VRQwi8RGpmPSMpImmSjiQ0fZSVG
hs4MmxOOloshu4XdH0K5jjbEEW3mk1STOCHPfx8POtbyaSnTBcW2CddmwKo6DUWd
/D0sWSF7oUvc4KWWovF6ysJ4rj55F+uy+Jq148pciotWNIErG4mO/NbFeHQyKpBc
KPifvzFW/28F/UVLpHrrobg9FTEHOMnMSjKIBWFGj3VMCvqKCh8SrLS3HkuFtBcX
tJw0MJrXjUq2f6VVWc6iTiYNp4sA3nItUYeflg3nRUFJGLgwoM+NX1o/7+W/UUVl
6IjU4dnNMpiuNWu6ljypQdCpYs0/4M0MNQGAdSLM9BaJEL8Kn5xFNiTiYdQmLU+h
vz+9syB+Zjgl5S4VqBxoHTr+nXezpTYmcoWmSC+LWhHW5UaXzoHCWf5c3+Otmbl3
23gqBnP9UQOpA8wv15Bi6Hjb0pw/dXnunLWEimfo6aHzgxX+rL5gsVKOv8Xykx3F
7xpK8bwEQapXHW/3IjLpwtcy/2o6emFCj4Rr9paK32YRMFNc6ycoW7oh4rXaK+aD
pEd+ZuL5K2oaoSy5lOmDL9B+8Y1upZPOqW8/WgstlFNrf+AhCO6LZt/waUgxyu96
9UzyVT3zJD4uBM48DM5OrON4JWCmSh8FVWfeoAEjfabK0QUnjhilccKQTbvAAP1Q
IRc02VRnmlOLsSVhIy7nz4pPH0Y9Ju4VuIHYV4TeBl1bgq/oZKjV94QcRQlMJK9a
tXfqQQ1cNZiod9CXSYrNfg4XbmxuNhJlZ42ADc/R/KaTdI5cLKcEZG1zXZPvf656
SuM/G7OgDYDpnW1IipwT85ebt1MCKX/7NCKwArueCc0Kn9rHrX/7a4J873GXPruR
L/hALdME6BHQymqLVuIGvvw6z4/qtMWTSjnHhAoaftnSULR5enyTr5lqjq0u1sRC
VTjHBe38xIzq2y5H3nTRlHGPdMg7840Fcuq/FdChbQFMWlnzwGnMldiTZQ5mSUux
J56EdxT6grM9Qfg/CJXZmq33ZuZkCRt18ZdzNXobx7/vg3FbhnNq1a/0ELk7nRSD
REYkQ4seCfp7lGIwD2tU7tiT54wP2J2YDRS/+xwNbQbJknywOk13blmUuVR3Hfas
qoYUMErVl5K7Vl8Uo9lpa9d/dc7EPxH86Ky2gqXePzCQ3+l1eShhkV7AqqBaHigv
CYPqMmNUtrWR07hk/CP53kdZ3omYonfg3tGbtfhDPfF7Fh2wx6xqqX1zG0yZS87S
6H3jX4SAQRQqpvuxyQYPReJ/h87H2DGkTGVp0YmIyNWLn+QP0bc482zHjwp31quD
XT6LQkwnfbp0CIwhyxtGIBwmCPFlQXZMLWQPN0FXVUtTwqxPGgal1BigcvHI955Q
bhnIJnu8V+8UPUeLnCQjrXEHBO9Ajt5RKwx0UVBwhCOVLPgPRhxXezkgEK0f6KIS
8ibqve4BgefONEpD/ktZOTzkpDJGEe06VOiSqa1HiieJi+yaNzWl5GtgSVBWcH2J
WbUDtQtxcK1XBLTcjhOj0Znvb8b8AtodFXrl+9GoVgzT/aEYnw///PXWCnPUEvgX
GeH+355I3qB2pU7/CwYl8vnvCA7aJzpZSybmUeg968Xnpc5mpZFYP95EChhe9m4S
4QFdSngcMXM92lOz6CDGYv3d7ethrkpthfy71UXOXi3zLNVT4seDJPOdgQDkbS8N
U/O7WdZJp2yg4YG8k8ElGxSAB4JifEGgvG/tVoK24jVZBhv5MifPBj6ngQYCLoAJ
0x2OMXqlVPOCT2ZyAUx2Pusa4lGQMNdX6tzN2du4ly5F2Rh/DaUeYkcwX9O2/01Z
Q52JBW8/vD7sC0n5sWh4ZirTredm8b4lgeotE44KAGwP58wO568N/ri8YtlCt2w9
NqWMtQHFXTH26ik63QzR4pDlozgic2Tgzhiauv7afvtgaiCxeqPftq3IpbfmjH9W
tsSlmfgdtaQnGMz5N/+pnvmNeLdlC4Vpydss6WwMF/6Mou47PxBdgc5cFEPzSq8V
hm+1b54OaKswf5PU1cWOe+eWxKV9XO6ryqs5fo7iT4SYBgdc/rXnyPsFl4lL0ETN
NZ2aOxVaUhOhKeES5IVaTaUaGm4oFGJp1IRyGZT44u9wG13ddaCkyPwWLiOLUZ53
0XfHztNfzTvhwBgQzb1idK56rWT/WNFxDYpRojBjrk6dVRixpniPgdgT96XMpnzi
buNwuOLvsqOLzbWXe3B3EwzzvAt4cVDK6vpq/X36Q4GxBwowLiyAwoaSP3hYvw7Q
SH0NFAFT0b7yCprwjQeyVfxPXB2j5DR2BFgLi1qIGE+sCSaAJn84K77JM7aNrBne
bGH/8Tqs1Eb7V6rhqqrAsCMJub9mi2jW6sLY5LWke+GAJExuIYUhCg7wFk8uMptb
LDbwpfKPhMiPOsbWiy/3RddSdYaxvWdJgdju69cJEHTakIjGXRV7gfTAwVcCRwk3
EOrmlrhA/MW/gp4MQXCm3FSq24Z/tJUQW4oZDEl00aY2vbo2JM5JqaYayWWGfhcU
mqFcXRtFHWXOhjHaqDaY/6JPnpTdgPZfbxf1yyyTNxUQ6oAX+JJ76vp0ne+oWSCW
OibPCU/XWnQadwG7JSggHvEl+QclDfM3r2R2yVQsmjG6Fy4QNH+GnE+U7Lr2E6/Q
uY+F04HRGhe8ijItCOgFGq174GCKtkxmQ7Gysqw6F8fXbnkKRiyuYQSWFCZx1XUQ
QPNZuNGGLRYrciRc8dyFWI1lSM6LLTe0DMo9bJKasP0+eff10S+qZMyI3GSvslZh
jYRCdK18iq2r937m8Rx21nU5DIMqO4gDtJdMQlMws2sF1A3o5kSiGl1OhbsLlOgY
DIbbbYfxk+ZM9jta73LN91wLIO4rU1YG2IHJ0X/gVIPTioN/LJyj0lKDl8ipVAA2
m01+cl64m6bHsecKF7is3IaUb/c25TF3ZWRF/yPzTniGC5THnxHdtEmT8axhexWR
CM/WYIczqjR3Lh4ozalA/NbIL5rrd6CXuX4IQGBwj2LavsB7OetM+rW11H11pVKN
rHSEWe6zJfhpI9E47y2xSPjVEXzOUdKayBuPApnCkF8zhz0nyqIGVqRac93UznlB
FXz2bCDu7IJ5CECd1FsWJcqVz8TbH8mKyyB/7ZXXVf4KzEeE3QStpOAmu1vsfyWV
hm9yZj6LO2rlNSdKQUUz6K1y+0SXDk8j6SOT1PiS4pPeQbPO+7v99IAnU/Ty0GAT
ox/EhdJIqEAVeqxw4LYXRz7kAU6OyrwD4Z+HpN0s9s4ZUxyri3GY7YylRMHW2SMO
NiQFOmPh9l67Vd+PSAShb2WMh7vNFUd59mPCYAahczpUIVLjVGSVs4JOYzQ2VODB
WPgy+CXJGHZU1BsC6rmqPnzXVer6hjT7yDOW6HV9u/FEOvXDZd10xH72ZNw4LwPB
w+YkFbNyTOjc2v1Fy96FeTKBqRhRxjgkt/QyvhTxxRIPL9BoITB6U8q15BDwoaCa
tPHh+35/SSPB/Kms/rzlkSScbsXeCudy60gGJIrNSJAOj1tVsOcB9EnBvQUI/vbu
6VzpNJxK04jfvJMVIbxbBJ/eGlxQm7e0gHIjJErX2lBL/XK8mJ37h/vtQGuPj5zS
8nTYUidghKp4tgSNbeW5Zkb3agTsHdJJAYyTTL5fBiQfPiIjLIVribnXvwe6t5Qf
sdcXwRZxwiWqBTyGdZ21fqv/y8FR/xg3jpgpZzJZEc3/BxD5W5aBwmc4mPN51iBE
vi88Df6CRgfZ+kC9q7UkoYk32FLyqs/Co8FgnGwfq3ZdyquePzIKxRrRCaNy8TAy
hiSwIiQfNFNoCv6z1g9/PQHbmTjWINH3/0IvBk/Lim9ggb4L7UOmF3D0lk8axV3P
7LeWySFfnlJVF0NbyHzU1Vgwfw2eMAWo31Nv7KHKZWzOFi07ixsL8HhZsOxzNjPz
jd5I+0uhIIPVFiumRHgEUCLezfsVQW+OeLDIxZD3usW4jqAh3FdLbeXuIblA4U2C
m1yTRsPB8vrImT2cMIkJokvXKDi5d+6xN6sPzd5tNrb3c823Nlkxs1VglWVEVBnn
Nhag+sQtOVvf65wMLmM4QX3dJhmkuOer+GGxcK2m6oIpy8hHumLESKXUVZ7tOyfV
z0hMRp0LcsvOao5j+Y+2vk2bPzBBh6OoKtbboqEjKD0XyOcSH5niqGR2IaeF8r3U
dkT/5Avo/yFN/MkIMuHp7nIBFdEeIQfPfzZzsej5+4jNyape/+IYqdQS5qu43DjA
ACzGyJSIi7Ph1gIht4Sywcwr3DUeU2hYv9/n/iL+GnHSjBHKpzCg7BZxSj9hHRck
CyTrrtKZD3MLB0A+Ze6AlEqT23p5s1/WCrcxHSEP43v48GElGCZ7cqsuN19DT+v2
HYiUnRMNCB21olv8El4fsjRCckSFKuAC3JsNqQP71awLH7Ow14iScdXYAydE1Xdh
376Bli1YtAwfZ/66kNVAbtiiqdzXGa/evnWTosd35+zHaOVwl+YCX52CRumx0fFT
nuPWZIQRGwAidXgVk8Uz8ULIhvvZMSDZd9ryweL49rtxRY2H0haLDiuYueDQ9k60
+i+zbWAnBC8OfGie8JWkloL+fc3zLCdewDsX55plp5HUasloAfhWCbhppZhDdLN7
vMy/CXXxl2EMzYzheTnPN5HOTtHm5sCuDmpaBoiNWGtHMTTROJR6/MRrxMM9gy8S
EkAR9Ye6JVll74wh6ZTuXn5WgpO7546C9aHuELpKp6tl+vKH2apHnBjfULXwF6gH
OABMCsY6NbKzMohUiGwVSVU2jXJYktNOcjcRctlJH5qgapP+QmU6LyrVrUt3Xc/L
xwOTknqAYzW3X5WAuXI6HOYU8elyjcqti751nbL/I+SHIPcLbRnLyPYQ8NjNbGM0
roWH4apwVKTxA47BnlmYjPKgBC7ythwoaZeuKKtrxrgc6Mv9lED/WMIi8TwQGOcp
QXit4pdDnw/TPwSankL934QWSuax7d1IU6lWt1xn4n8gmp+4mNTrKtt5O7cv/yMD
NaS7AfSmtFoekTPcvCCPOmDDEpY5EdEz+mSqQUJSIUPXpJnFbU+/xhjqkATo0QOH
Gp8vWT+BjqiFIltyg0t6ua6xTY6sj0j9QoNYKaarLHWk+inDTO5NAbAIzb+XTgAA
GXXRKUuO7bHVybGwf0tSut3Vtug7Z4KEnXx1B6nP34tORlcIXv9WoQMInKCWsOg/
ufh0Czb9tetu9lMKPH1nT/tozSAAYd6H+pyDwmOX67RS+ICF+yE1ThQ1wqoS4Egw
9SZwxyHDHya9w3FSmt9olT/IE7yJWPIT02FaQoo9YfabVXi9iH5B30wzJq8oyjhM
PjKFiFn1XtFncCVX0MDB3gO9Tdrz6yGevrpVCcPlfAsYCZ93Vs0OpuItdHa27mrn
O2WY0vGXo+U3H1VMKecWFyvvDpXESJQYcJIU6W1oKDXD8yeYwqKuv9SwPN5Dk3CW
PwTbDyonHwpc7FYmSYzpc8No8qPJOrGargC2GienDuYCTBiQ90LyWQPFsVHvDxMX
BlQGuop7sW4BXCQbAR3fW5L8Se0iyACK0FUOhDNGfBxSW9Ak0W8LdcrBIsDzwwO6
LPfiKFqHwIolsnzrLzYJ4HMZp+7E5us3uCMqJHq66iFgP03GyauYzJITABzTwcoW
0MwvPjzLKO/STpqwyV63eOjS7tq35t9iWx0zPY8CSo4iexqgAIdSnYUh+libOplw
ASyHZFUEsZVFaerst9YHRjlZlrY6Ykul4L4fA1jpHIpGi8FODSOWOv4EGaIqmOcw
XnZsf3pV2eYUH9R4blvBJdxf8b6EpmeMzU/VWV+dM4ZqYasLUs0KZb4tOjLj6rky
13R2LUj+oqElbm7KvKMuQWUi9JqmM8PVSINoYepMnIPuIusaNzQsl7TowyLcEvGQ
ZYprEP7cgfDQh01EA3P5x1CuwaQ4y7uSzJGeegkmhZUWFH/dPy05SA4gSJ2Brj4n
qMEh3Vh6ZEupPVZDhzI/MUoYpk5FHu85Bx749Nm+wQZtehpVAE43shgfKaGTdyH2
1yj5ZxOb0Onm7rx2kAkA6uCDTLkjPIkH/7Km9KZvpRaGS4SQnCuCKmDRHNsgznHo
SLTlcIRr8gg0wFnr1Wp/Me+q6Od3oHMjAk04riMshq2PtqQCr3M5/Es+1QvZznut
Lj3otGxcj6fI+juLwCZSX8H3suzAQSKQkQdtsyF0Bd90oM+aDM334GkbBX5wLw6o
X8GSR1Sa6UrBKQlIJuJY0wd2wc8zDBedorNaMoQgY1IMxSdWNsInCOPGlu2RMK1Z
A4b9oFDTBs3L/K/9pQnOLDbDWfdnK60J7MpUQdx0M+sZ1eZTaogTbcQ3YYXKf76D
OqVgOs5MayJ+4WWrEpyqvyWoDT9wFXO/nn6TLEZ0Scld4NmGE0xjVRMSsv9yAZG0
tARUT9SznR/KkLP0h8omCj1TN8rn5yrTwa+jSi7IJD0u0N9OrgYtINBvHgIDdVPE
qvzRWyUAB5w07Yg41h18TSjvhh3w8pw0IHBB3PkZAP/G6ooWYhlK+syCqBE4dMc1
CGjbOoo5Kpyc0OGfoIh3gQSqHdTNihkByH2PnUn/NCt3be8WYbyxvyrk57dIeklg
9ie//ah+fV0yJushSlGPZ+vN6rrUIdp+QKj5FG85wI0VkOGQSHz/zr8RdCzFks0K
lVkdqd1IIUYf6DywlJzmb5VXYgEqNBxKH2sOJeMk95V4G8PA6FhCo4PRx4KAsp70
hxA1V9gE+fCJf3KqlWujX1cm2pKXG8brHCHC1+NRLjKioTAWpyqZJF/7xBwXmljy
1HY1SLm6W3HvwO7lxKU4xP51r46xg6FwdOHW+KJwmLJi6seEjIffPfL95J31V1aZ
9GbZn1sNOjzVuQoHCS0IptM69pXQIE1X/P6e3HvASHLVRObWv339NmM3qABeG0ok
SdIvwafo47dOG9eK29yqEee7gN/RvByjBykc7ZJ9Kv1JTGu1GNY2YPMW0T6X0blN
a5ZUefVIAjVoe3GrPg6sc6xcKsumyA4xGEvM5AdnK5Va452v31m8w72WYOsLL+O4
hN9/UczxrddDRXI4RCRGKjzeEVSJHOAiemFvCYbaM13QgJyO+73oE78j5RdA2nlL
oeWgUitiWTLk3fv4dYk7Ke0T93FceA9Uf7ueG61s++L42md7Nmga/noQsavjzE8r
xiRy1sZHNxyw0q7YDmyO8aSPbSCV2/MRnE1ayhhzqUrOzQHKb66kQE4AGqo3WBBo
OjVwE4Baa2ov9bg6Ctt1JYDl9q9kpZlOI9KSUidEG+kfMGwls7PpHIJmly4RV0Ol
ND5yb6P8R/Zq9xk9Oa67mXejhap0gRyqUjGizvpvIfGuq2TgLC7rT5Y3T5y1C80R
6BYeHK9wS+pJju9c1naENAPJlN3H9kt1NakTai9K1wlZgrFPxRNgcjQ+1rQpz7U2
VWeIfpC0lkWOvhinehs0lpyegpx9G3sbjXv92mvpvxkX6hLCYJrN7O5OmpDxM63F
dfD5m5xb85F3jnqEee9QAshIxNVlzV+Q7/F7XoVlBMG3dxHaCCx5ylyPM9tP5u52
i2OPZU+MhoqXre3pucG/XUNgNauk9K0YG5pInMNJUsU1cSuZAcXTzN/Xv/SsBMaN
dnIpPNfHTfuf/bHpz7SEP4XvKCQQkeRiQ/fI8W/ENWuQ/uqS1gHGZipjluKIalkh
6XXkNAP+1cFNXbgdVGaBd6/CvqQG0k8Jh6PxbbTOSzxzK0D07vR3XDAmmoHKBR2c
2QIBVrc8pbOqiCxXT8p1agaW5kqrdU+Bmm/F1dTVLZ4H9ZZZpID2ikmBlKbE4hG2
IyvjMktj7CvY+zwruaeEx+SUzEOZThnFO1rRPiXghnfT6Osl21ghppHlumt7Zs76
NWj4XK/+KB7Y3A+20F7YSURSwKxK9nyKrZEFudwB76By2+U/zpAuTWHbdFavz/ME
7vMMPbh1oX9+rEtYevaMvB15o/S3lXR1nLnZ62lVloHp9jEhhiAUSxoJ73b2aN1Z
fQgzZwUKogdkTbOsCXUA1wEHNUCp2d/1IyEtOAv+mIk4XT8FYyQMxNelPygRYXeN
DpPIPvZEXSBA179slIHTJ9PLO3Sj/IJ3tTq351gDNVvNPjuuzufoPzLkC1FKlJ1G
PscPlqn7s1C0PX7IoX4J+J2g4Pmxk3QJlkAnI9OFh0pL+grwpFBGrxU+ZdPXVVK0
Tj8jpxJiNyUYaZ5SgxY5547dXJJmzgjGWTOTD8Iyhp5VEX8SLz6QeOJMYe0kbPP4
mmooBaJHvNlAR7G84BilNdZ1+PA91OdMrkEbYyl9d8e284Q2zfs0xpUdW9mVX1FI
wtLlEksb+mJY79bFCd/dAMLwPYr9SnN73bVeOjORoYVDBqGIMr8kfsuPq0yszgod
JYZTj9AaAepjRswX11doT6QIpUHGe5IyOrVlMcnI5pWwRBRwh40M7PpqeWygX6wa
ScoUWYWsnlE09oQ5/2wsU8RaSKf16lS0+dlV21gHgVRlWFcTUPvfhXOtAOyXXQil
T4/AYB/5o/BnWB+bvO4YNmVJuSKWt2CPh2veqOSqHNFTDAQODTCe8tf1ty8kyfuh
2BeoPhoB+m7ui4EEDdQzsjLMYmvZMwBkcqOSiTGlUnz/lkX+6aBfEOPpTNJ7OCyk
XRQHo7AKgv8Nz5sSS0DpTu4tiXxZwMB9n9i8UuiovIudQFLZy6WOtvunEd9SX31y
F7FK94HYnFL/TuqC7QP6DbVEKUdy9rrpi86OT7L4/JRo15fu5qHXfIw1hT/QuAP9
SIFkQ8ZS5lbAZlRuWnpoxPRnQRE2sV1Ewwfvobxi7ShV7e5CU0Q93FqTqSl/1xUY
kL9cBViztwz5ZjZTnjLkuFbHWAiX442Tv7Rbuz/vHE7apxVj0wo7e9Q9umjtDnTQ
M3B/i8tBSt6Q7fw57c6sCS3CBQNXQ0MYfkAIqOw2XFJxtGEzu0CGmScy1x7x/Pf+
89S0vlGS6/iBR81YTqxWW5GNggou3GXv2sTv9NI4TyHDEcuoQI86pJH6rrnUg0h6
AacRgIw/RagiW2y1w8b0XkXDrEyTYGPoOKJnGwy0NQvbD17oK9Lzyv3GVkIBvRPz
f5pUaG4cZsveBM1Pz/x9qG9Mie7SLQZMcpfkjcJtvFGeH0XdFdEhF1mYIKSbvox0
rTDKDP4cGI2OFKYESR70N1GU1e/B7SM4tpYKM19U4MJVuCCUyll2qH9772AP0bpw
jgpPrPqBB0IhVtKQYiIvWay8VzeQqyZzTQ6iiuB3tzU0FhnS6dSEeKeIZJHBZHbi
g6L6nI0zKYxmRm/ax10cUaOQc32vYBavM8yQCBhdV6inXd6I9321ZpW+xIAUYvST
kNt3eJ2Soq3imvkIeggRM6378fc2whzahmQJrXOCRMR02WzOajrH+X2x7urc6/ab
KH0JM2tT7GLweiVyZwvF7IjW/j1uMR2WSx1xvPMS2xZghZeGDWoM+h5CCXQ1Il6h
7GnhorQfJIuFFgRKpbWPhH4kHa5XrJH6vFvkmxIYk8BukSU0uU0EU3EIsuMk5HjN
easmsKFhlSKrqm/hNISbaqy8tKodNSCWY9K9wRoCegOmSMWWiiss83dDroN7dyKt
4nL3pP/sR+87oxpqf+Qbdi8yJ0ObBwbDD8P2f03zBD5lkXy7vD8iQBMrkCgdhdxV
kYItyqzv6ZAwTBZx0wFLEvedbatqQ5L/Le3rWFF+a85tv6bEYaIQsizLpC8fugt/
9vDfdYB1Lt0ehpOEzTDoUm+eiTVEJ6NHaS1Y8iwQeO2PC2+zo2FqoVil93/mx6jV
sSVZrbl3b5JaN3oLSd5yqYtqH/enm+wNm7lWD8k4AISIzKSJUjO6fivQyZ5ixhrL
ILtNr5mmPD2xKRpo2C9ml+PVPRGcKfx7quoTRuoDwF0bJ9aWQGZ9c1/aVeN6KlBS
udh9PNnErXBjfqX47ws8hDR3jC4S+YmgGKkrp9hjJ1GogaykkvxWZDF4Pa8z/LkE
3dd0EC0lt5PvlpCT/SSx4y6TfU14E0R1+sC9UWkrtrEdmN/neT7xttz+nL77CcXR
ufXSb1aEOZXGWuUQsTJz96MDXQrseKvQpz2hMRJGdfWxrHl4TTteKvOQ5Olt4BL6
ITTm/yNHDYSlsKHuNTEpyu9tN6gdh9UcX3WUDANCV87eFWlpn4cH+0L5YjsAT9YP
zsFwFuc/077K4Rrqaf/KzgptW+xI8IGXK+EuD4M94xgJ+xvrFoOeJUoXzvbHyv8Q
msMTsikcOL8yuVVPjNmrEobfjTJuOSG8I0AIwHJnxDNouVIjk/rUf+zwyjxpUe7j
HCuk6dgAS+mZCL/TquMD7MWwFk+zs7jmVOWJUHtWwohJwFk1O6GeENPBXKgMi1BV
herkMQ/DfbKFtpco4rKRjTxtZGB2UAEjJQq+8awfW7DWyoyvdFBEsVNbuHXIuCl4
TjUcLQFX8cJzc18W0eRvMfUOQuvsTykw1LX4SqY5i0xUmlnnubxu1j/vDwk3PIeo
NeKpmw2e9tcS42c30t0M6DdyJ0mwx2H1X6lacOF95Qc9Glt1+XPXiApgEB9P3SlJ
DqnisjWedFinHbMoTOczJOZuFWWHj9HhwaYsw5j4YhegQijCmvw1HE8visL10Nv6
FND+n7DOXRR9NNRheapr3bUdR1SVgZhpih7bLvwrw6azqXDxq6aNQCEtoEoSpzBR
sSliJqmaNELvqXXo1EAWAF9S4G+cYNuLdWy/NCkPiiA8oiZrDvZMtqZrv0/nhiKU
A5n7lCHYRrU6AEuERKB58d/8uSeGpUGH4DL5ExJVARlEUlqukI/KEJOv1hCL9qYT
lPfenrtbT/g1OqRTWqegq0gW+2RATorC11ZPtSoHPqtpNTAUrYLLzy22IV2atYpA
CTHquP/coL2BhvvtgUU9Flfcm2yYlu7iSFKUW+mMlkOcq6viKrmGYbaKRWTnNFpx
95tC8TQqgGg3DpmKgF7Ksmf60UToaZFgKT4VkzPbiPHynICLAz7rdXIVQinJYZpX
KOAIEQZcOUPXPo6qudB0B5XEmfNq3IOx9BU3Y8W1Sp4Es9NjGZLWC9g5e04zkl/l
tDLpY7HV4QXSkNcsCjOnT/qiBvwgojj2Ejggj0IPl0cN7oyi7k0kSrhZINc3x5L5
ftf70Q7YknzZfUaZvteFuGlYMSpAYskFFBgExO6tsGxC+hrtb47YNNT1mqcCRHXM
HVkVpJ3LHgbOuDNzvGEo0eQe/mD1U4PcevF36N0DE7z2DVNLZz8HYDIDKe3YP21/
7nwfxla87wZ86hxAc1K5gMHt5MsDpkoaXa5X+kicc1n8yHn2sTeCLtY+p7hJlBrp
0zPJrW/LdsJ0pcmd2gkNN6QD63wMAH9gcAgP/4LFQcpklR+qTBPZtPbitX2CEgbf
sBL4dvwv2PXbQ+sw4di6m9Lw72yrnEi0gdfHRDheLYTjw547e6itDuDzzkhY7yQu
/Ne3lwssAUWGFJSaFizVY0bus66sBjSC5xjqe8W3xZ5UNqh9ClRzDgawbVJu2uhj
IHap6Pt+8J1NRXYp1lSESxlyv9KAZ72QVpCQzpIZbSwBJjdN3qBDqS40FlV40X9H
oSVnH9snFwJAykxd+EEs9lWvwWIVjXOJZe+J0xl5nKq57K3PVFfX8Xpimld1gw+v
omh4M0OIAU86xPxASNZSXBLdLbzveTjREQJUv8ZfZ0aT2dKpj5rGN3Tm7zlvwCI4
nT2HNCYBMuOilZZ+XJepO+6X2ureJYXjdBb3DGQp1Gcqk6RUP3nicVlo7h9xf/Tm
JtlZaJA6SiylOhbSEGHNb39R/mSu49Uerpio6dKbhuBGj+ii8L94qcvnJemaYpUl
ExsD3jlBLDVm12UfJANi5/lade3MHljOiRXnh3qrZ5baiN5KGtoz1Vsf2PGhZwND
rOB67JrckjjYSSGpfxDCkRTEQG8eCPjCpb2mwEvQDaRFc0VvjQChAawgwF3SBeJ/
GE8g68yj1SIVAFPYmXg5EpC+iwjfX1zvQvzWvBKKRn/ZWKILaa8t2rg18NFrz0hM
Ic2BUNN/JY0g6Zvh9kSxVpRLMupoopdFUlvNjGwHBB96HWyjMsvtnTdyNHv72eIw
j5UYFsfV3RcxHka7CexDqHtLyAthZ+IUyFRMdsBqMopAi1cmFlJMEWguNZhfQSmS
5E+JYMts0QG1CWBNcAURcfAiUY8CC6THFX2IlPrm2dBe/QrDUVpZUhdkynx5I+v1
fToJRQoQAygcWuPgty2hnhgWmaI1JU/YJVfx5qGN/MFsDPaN41eolfeFxPbnjFxB
1U7nh6dg41DwXrUa4Qf0cjrw+KnVJW3kGUh1lhHpVQn6EohAulE5EXvXg5hSQDyw
MB9DTacH4vH9EUQ4hVXPWTqxR+VLw6Y3sM9xrWbpm2kzzHzUlSipc7fCG181a9vf
VswrVw7o9/IjKET6/ofrQijhhur6jDMhvCq4lFLbBaODZoKEHH0+kQiz7QFfVkpX
mCQXvjjlvSWmykSEN82x6l91E2a+lX2mMcFaaPCK0E7PEpnmRLA3Edyxe+/px/Yb
yC8HgqVBis83rhltodFe9tmb2o43NwfhLfolC1dbLDXGq5Sfuilvls34zxiNodMt
JcDwY7mMMCaTJifLbwRy9/YwqYgJauGLkWPMZ7rBNAjgEdYWx+CTTerJDZtlnNwV
nn2482JYqi/V8etiIm9Ms6hlROmIl7eLkqqV6+YYb1G0eKuwuf22GjPs/gJT3YRN
euGt4ZBMwRzwYVW62wk7W5JKLAaJIuNvEtkYuIeB8zpv+xTDk3n07GJf5Yb8WWtC
cYy9N4q7aUUR9sNxKc2oieQuDCyMnHdKu+evrz/h+nf6g8qDAqM5Ynhw6a5NSlIh
O5zhYzUNV9ZSaBo85vvL0ciJ57Oq85tBLD3j9nBO/JnTtDyBOccwgyYFodSn8xlO
xBFfnaJ6qCn7d2EMHrV4W0/sH/UFtyOyZ9+WnOyYpMJl2qdnpMWycFvNcCcT4GZM
CLjzmTcAssbtns1+wwmM0gyGAEqv6ibnvA7+GIqJRc5wqwDux5hbJedAljG/lkKi
Jf3dnpXnSt/NXX3XKm8cO21471NXktVrLdLeVX8Qj7+RalGUr21dr0WtYQ4sRnlX
2V8Yqy2uCZdIdy+T0bp23JANQDRnTQxZpNcXnNgiieAEzNzXKdzWCMQAXRHkXhYc
ntryzxMkT5sRg8uKhA1/zQPo45PzLu7ygLGk7/Mch9Awrhn3BkzeDh1gk7xhrdxp
xzMBCExA0NfFA9Nx1/20XUIMn8Bpwede6CcqCpbEFNEN1PV43MfoRQbZRzr2ACYg
oJ4wOUNJh6g8VRSUpr8+tUYbrNoXHw3KGsDmmKmbsQWpUzBV698eN/dDSN0P8qIL
xTua98CF1ZjHq5AJ0Ko4wYgSJZxduKZUuSkqTz+gIeNPZVCKWauDd4LBlTfZ+r6A
TTWeaAfuBV7LvjANIARN6VwE9dF8r7ZBCBgfUEPqIQsCGVVqHmMRwqrQNWqnLLxE
UfuT6aUrUQaAGelSvx6fxzqeSiWd0BWbNPjXwGJjlW7UgHlfupQwFyjpraDI6rRh
jKKFdTgmAN6n8j7oNgft+Udqpq4Bo7MkshC1MnxHSFeHWtgPZvipJGFcx+TWvhCT
7ukob8lZv13U97JiacdZ2XidCPopMB2dSAnuQUZvMOXPqJ4lK9WthIejaB7FVu/t
JDXITRigNQu815MfJ3oL09gc/GVBSzo1jbqkzyDVP0nx2Y6fulh0W8++brXaK/QD
jHt+7WNzOuJThYmZd0NTi61XCCs8oVTZmMlEvnsq4HTQ1ekH1S4Wi3/8mjjh/iP7
SQbb1PknDlyVbLZchXbI9q7lpYB6NEOKDzt93dXj/wGh6tKrbtjAF35w7rJczMk6
8pNq4M0V9EAtxMIc/47DK2wqgEQtheRHGzhIDtkWVxR+ByZL84ulER9OX2FG5N6Z
SoqDTiLhvRSpdhFSa3ZX02eQwxFkt4NQ6bTQDY15IsTMGIgrOpSnK7FU5Seavtby
1nnPYXuxnXttUnlGJ8VVALk0CZKdxlR8YUTP2P2NKZFy7nMXjEOipnhcNY/x18Kk
dFc7D0yrvUEGZngsPvUeI+56S//cOvbLrAyqM0SxeT2cx8vcGpPhGhKT+OxU4kHh
G4egvJDGMY/EaTB4qS9p6fhn/FSvz70evEkCm6mDTuRNJfWwI7z1timFpZ13J7q7
RqiN3VSW1HeL/x9X3+zgI9L25iUdWfP3aAllNGmcZAeHLpmtYLKQQYhe7kxeOUWx
CshHWm2oZHrvtSxzKb0mbLkj6Bn2+W7jj4R/k+lTZJRsqfZleKKHKnuskvKXKOKE
RH7gArNK2U8OXBgUO3pgCgDAHyAdHeZeiMEao2/9qylD9C5fbbmwnVeMCCldrOe5
fBUaIH2uBOPQNihlQRN/gayGJ+eaF3bm8LrYwK1VAlTpP/TUzfjD+eW9nK9TU36V
CuxiSGBNDCzAeMyz1ndpiNLEHU/hFdVsdbHe01MUJ8Bqq8aTqhwngA+34bKGq8Vw
enEvCmVik4FpoA4Wc5V9t93fAOmUg4lft7oC3zC9ECVF7YQtoOIfehXdeHit76Nd
gFJTmLH+ZUowqz3Uo9cSgxwhMONzbFI55zQmc9DiKr6FeWq9uU7g5wZfsZ0EIzG/
QcU0jHylwMQFkivSeo9M6z5q8I7Z9eSZOf3gPz8anEHljvKFl4+XB+3tX1vek6DB
h7EIPW4XROgd4vwJ+vIcoqz0INGW8wkZirhirLy81KQ9bAHSO9RvBreTyPeH1aCN
AAFZO5Vd2ZT4ZmeH5tas+koRzzfV+Jv+iwxWFy9Winhk0UomgpaPD76q5+7IRT9I
NbGvmd1tcTa7iaqEGf1jaVbQMPpattAlfp7hffM5p6nZ4fkaCpAQj3mOn/u/ZWMN
I6ORHgnY0sVWCzxtFiZ9H37POf2N8ZZ0lLqKCUZrFK8ywC0YjFfDSe10D4aeKSLm
24TAwHjFeUDXGC2FO35Y9xzC20jKq+Cn9xvryzyOVgna8GefaHXHlxedeDxoQ5u2
w3YBfGxnvxiyQQcQM4ZCw92Gcpf9SZpVO9Qqn9Y65Cj8x/Xt3kEVnfo/z1PX6shL
tmTS540Bgu4zUsXmB1J3vEqvr/O0V9JcAvoa6NRjsF0X9nNIZSyJaB4lOsppXebX
LjnSvb9Md79HsQgbysB8W3AVhVv53Jsqfq1S3ZYKJ73HtKKuzLHFn5QnEBxlq0Fk
F+b90vjtr6ZGHcwCqyd38inzyfBrRspqNR1glK22KxQJOAdILIi/la7+qOBur0lJ
MPlYELiYlBbdRwE0T+ymiYhXJVccSdQl4MKiAQKqJBzRKqFJzuFTWqicZBJr3gge
cmFs+XnDdQ3NbE3mlMUyDAiFp+R4ToMywN2nkgRWuv4xU19T0hxFZ6edYeZwgL4q
4u4y47KxL3RJIzf1QqY7/WRO9pMwykKw4todNLD9HOG4LuqnFyBrwScS5y8RVbXY
1dneee3yzKujW9ik4w1h86+xKAQ60WYwrE6sGzMwd+8/S7PEBXKG8f61CkVgCt64
V08hN88NAX3FYYHWSoUj8Gdu1E7dJx7MqSDQdMkdaro6g7ndmFYBi8R4NYW0yS3a
MPuyfxICrMedfnmGpe+eOILNoPCysIl5IB0u3/Rsa3Q9+Qt7tn5JcVyyAUQz8vOL
478CVR820Ys1c6Sd73Vnw6GK84FV43zPmrtlmqK08Ki2j8IGsmnIlO7pMxa06/Gr
HikPMTB11CPJcTuG9LqZKxALSTZ8QPyyXoTSOaNchbSHMgUsJziY9Mm15vSUn0FU
OmuC4X5P3VwfPfq46YDbRHmXYa+JO/2ovO59nYmPIE+r5PlHkQaRSpcEe3AUDT2/
SOt0F8J3N0zpYlgjEzoY+TGDtF7Q1NBdcgZOYPQw/kMBneQjx3jrgGU+4sRPR/Hh
i3fsto8HIpDLEQbJTbAituMlpU8jpPX6ViY/oL5iCSHHFL9GoirpmlpIB4WVW4p/
kpPJDdn+1BK+P5j8eBcxEoFBeMgvKuiPlC2xsHrUhrHuyoQZXsHh/+X3bwHdra33
5RbD/JcWY4DbWofn//A0HejNEaexgV8T/BdW0gELAnABy1eizDw4PBYu5ZU/x4ha
EUe08Oa9xwO/xeAWgG1xJ0JZoZMe3zvh9KgWAP1Srs9BZX2O7BNOJ7vXv0rvhAx9
GCM+Cy8hu5j7uuPGIV542SYaX2vpQTwJMm13vxYuaZ3tnRTzCMTKQ1W/ecp926hx
+WBXFBx5ODkEIy5A5DBEFMc5DwzfMfiM8Y9Nftx4PZlLPacSqy2BoWs54JSCxUy7
jhWJ9NaYAGFavLkjgj4wuOXjgW0zDg54uvLgZxDpFnYjRWOI2H4yE3MmUEkv5Ris
BZU0Bis8snCscORXcL8lnynfQVoU+8sKpzQSC3mxJCMKFrMJa9/iyQDA8JVGHpkq
/17nmfdDsBSqi9q2jatHaFAWp4lbttKQi/yzrc5a1mvGj3Jzvf1WTHfju3fP/Nnd
+fPpKyo8gMgA9Yi9GDxqVYrKJxCeTqVbUUThf7DtVGj3tFj1FPYqVNM2ZxiJhCeq
FzNgNo//+1OYJGNRLGzs6j4mpuk33NEYrtyoZz+TjgOiS0DKDsP4Fr0hEXLBSBkH
+jbSBRun1Unq6kiCZvO6rOahLPpQJNp3OzkX/x8V2VQvO7Fi7kFiDYV3kdUVAvwc
UeQdkmtfQn+HAHz3SczXjaTyv2MVsFPHur7LK4FQSzhdEwUT9IpbRk7ZdR3qE7XA
vzBGi9UrtBr4rldQXRXfAXpRjuCkOjCCWctY+5mjmBemRf0ILgDFSushJ2UI7rjA
hvWLGanlVnJFBMAtNh5ZaU3L3K2MFyYk3+WhFxZzJxmcxMSw6uc79XZRkfBLTSXp
eXxKgXJ6JQkdL+nFXdSUg5stP27mswYSLIfP1yoY0HuII8/DnJfqPZrneOrxpKnB
hdKC0a0vVk9ucPhFN2iy0HQuPHc7QeSNIv6VgYyAhfR+hQcJlPkcZAeu9/smcJmb
6PPcpN05fU2Fdy222VyYI5X2axNPgdAxaYRRffcAQdya5vfLyDdsrGPUYjMIHKgC
9T+p8CcY2KSY/fNEJBAPDvj2dc3XIIlOtXHeyoP6x8ZJ72fZCHgd63DJUqo4mbKN
QEN4Ls4j6favyt96lmjSDr7X3J+o7P2ceU7xgevArDHym9qjrBF8oYhkkB1ei1Ui
9gu8Ru16e6J1GoPJNjSImvWlimoYU4Qq3rRNejDRA4ej2Z9knBzvDxhZXhG6WsGB
TkkrecXGr+lmsR+Z6ID6cWofBxcaQ8TaIB93H1RE3KGs3Ab3Pg+lx/iKK+YUcLta
YDFA38m6i7BjCiEhDwTdqswXyJl35eYXw3H+kOlWiI8QPV0m/DZoG/njnptVpbm3
/uQky6ET6IVIG+dwWmGb8M5yKfTKUFplrhYzsgBAQiJBnZQwsPOyp/SuDfCsm6wM
Unwfyob82+VMKoBWGaLKzO4AgP9bJsEnuqAa1bzEiFPBYizldndqwD5uUFwPeoGf
eDOEZD4D8jWW6hulX0bsjjAKyUj2GngR+7JMxPYNx0dKA8GucDUmLu/NTClrnoNT
TsmzFI3scnlnD1UAAdOToQ1tEXxPEUf3tC2sxDrYFm9aDTvJ/0+CXzI2WFEZZwWP
EbbVvAQAO74ZJrYCTBC/A8nzJCE+ypVUtgUB/ACXpcKC6WnXWPdUNSS1C1Jrty5p
krw2w80l0JkWFio+FEdyE0s3mXRh1CasypdSpM8sYlqzSCz1X15+Imh+6pxquIzX
VLjtx9H0B/Y6YCMsgTdIN/5Ve1Rimva7fCIYqmmcpdpOJytpnWBRFNsd+Tgs/WnU
Sov7MuRcYzKtPWknA4MeyXx7VTXl4eJ7TIci9ZE6/VXm07ig+Ap2ouUhT3D5Kspt
uUJ1FX+x4c9f9DqA/fs8d0QZEYYiR/N5lg+krpjTf1vsLRsdyuVRqcGfAztYHO4G
xz+86PdUwYQ7LFKFglw1B+6r4Do/s2Duu++2ekx5DtSr48gUT46PaE+dZ5mdQH+C
lfiTVKAcefefttoHovv3c5NS2fXhUABdU9LG9eBtHWq8cphISXkm30K6RlvSeRIt
U7258IfgQ8L7gF0rjg89244Y8f7iuw5x0zaTaw7caEIQNoPiCftUft0fEBAnmwzf
bzfqO1DhLf40Xdm+Y5eIy58pGQoatVfhUcZ+Uer7uNZnb4zZWvmlFHZXRnjNJ+Ow
8275m1YxwdNeQfhQbRhTP4PLMYXHnHB4WoIkCVnfaYYnBt22xlsWwzuFwDVMwFBt
KpPhpuZnM2SSS3Uu9i79pYrczSqfQeBAT0EslGeKwdqD5XqKRfV7XSWe0/a7Qgnk
vdAzQY4aY77ut4d7JSBY1gpwGPRfXtqruFs5Nqh2ZSLoVsVyXh8sgQ4ET4JxUFfA
C/82eIFJXe45ItURUaOZ1myshMMHxI62s6fmDlV+GERfbs8OOHRGYQ6hLkNB/Oum
G0MR9JbzxAN+6PgG/9E7lMMvbLOW+Zh5WcbNS1zL1Ntks+Ch6ONE2aXsYllBr40o
PYXJ83JHQ/a6By7t7KJVN5LAmTgzYlLaC/CRMO0AS2qcheVv1aHD+eP1vQ8kJUGv
34JK648A5QVf+i4yFoXoYnitCafU4Ugc28cb2/yXgzy/wgXfNgkqzLMAxHvr4rQD
vudmEV0qEUAJVH83we4x7uiAdd7H92wXjsEluM0gbONibE1seDOfO6fBqv0loqN0
YUKGNzZ1hxZQs5w7jUZymBVs4B5f7thjV6v/Qz2GxGG0HqdLbaZLw8Dqr1dJX0eb
TaDk7vAKM+dxxnkiih39QjFA0e4MZshb4ej5bMLcwNq/BJd9yrG6/R73PhPI4OwU
X8Ft22bYrP3J+TycNi0hsbFXNuGgg4nsxd/6t5RrVUf7+PhMWi1+KIR2Y5tJZ/ds
uoUSDSWfnupwWQQoDonVs0B+UJjUeRol2KhTtmdBgkvE8ZGPYOMb+VKtK5PKSgFH
toL0nybhM1p/dWC1Bd3r16W1zYlVONqTyPYvMGVFYAtvXFFZKBgeyutZNFfH9PlT
e9DMpg/lFwpf2ow75Dyl0eKyQ6m5JnhK4mME/A7tFym8gj0NHJyIcaKQFDb9wkGc
rxE+PmqfURpX4EyRaCm3nam10RP4C1pALOjzEWZJO8vpoZ5UdRTo+E0GlFPZ+nbK
1SruKpBPYsdG3aSFrvO7NthOdOaO/gV76gEoukN5gOOvnZ7V7RRNXdbdbZ+ihfnB
DrMfX28S5aawHhXJeZP7EFfqQf80sV0E5iySNVBQLSlIMMdRfWz/AdAmKQ+KaYsa
53qpBYSGlPHOPnOcpegqxRnunMSpPvdsyzmZs/Pitg7hr4SqMC3s/EdYLCd690NP
gFOxvGhYx8rQnlofqjOHftNI4M/JbqfxQUHVe0FC/ziyTF6G5Ltf6co7VLLXQ7R1
7xGqImif+GkPiIvJmwm3r0qEK/sGjiKztnJJIHf8WPHH7i9ksHwOyH/jx9MNzDbB
G5jDdVqXtCEqLw1QaycIQCu1DJXkKHLQh2WxIqkpHR6hR7XlhjlyMTCDGcuoYV79
uH/hazVTz3DEOsFRdzGRGIr+h9lO7mXvHBbPwR7AYpeOOhAaSnbOyFO/bSjNCv8X
p7+BibMd5vnFLwcELTnMl1dWqNRU5g93fpMXEzWlTKR2XckW9utV1grN2ysYfyQ7
QY6+ijoTTlDm8lJ3V07mtPeMq2fZbntFEfZrGGc7YzoVN/mtS85EPR/j8kNyG1sw
0c6MT+Gwl+NZfNMFGpAWWdxviBnCsOyOnCGsi9U4M6tP2errI+f5bfNp9fyYw+vR
g5tkwVQHMSvLQkXHtFmiJluEZcRxAlntlTteqKr1zQ5k6keMUr4vM8UMahKOBTiS
/ZZ+F97DxcNdmVBx99PIDY9ce3ek3YBHheRDog1LflQMvy3PmDga3S7PAmlebU6N
t4lMnHXyZESMhquiuNUbuz+svJUBgGRlzgGkN5tmFGr/EsiH62C8/3Hw+o0hV8x6
zpjXewjgVd2A8LsxMFq4dE3DXSDPQsrmKiXyrn+edje1N4T7BkdHfTADYqzt0NFj
exW+OM++P0Id1g0pchk5hMhZsb9mFb2DCf7gkjt43tOSxNGI25s/MO9DYFtsyO7j
M9+3zCzYD44a+ETHE3N8WCbwU3cuh16mddZeYQlgIpYdgUHYHALOci1PELsXNzus
W3qmW0UDVvrqd+YBMu3PLJK1ZPXf1aMbBpmzlel3I38R+umGtPcLLx0Wk0XLbn6r
3itPUJ+eWnCRKDH6ovWJX/EU8H0zLLU1VXcPiDuupweqf1w48KMWq7g42JPL2tW/
YWix9xWIVq2/MxjM0QgJsmZx7Dw5Xgy7yZjwKk/Me+ejoRhLjC28slUA9/6+vzts
JaGGLml4xGhk1+FTWy4R66eagACtg86s5rb+yNH3S/rEyuFrFVrMgD1UsVQuWfj7
kISjhNWa5JqN0IKxsJ7hcns10Aqvg5t5R+rt7AihD8+BAU4JBH2Cxn86tsL/JwIa
HFSyMOTRfpTjAaQJcfsM0DxTDGI+9ioVxDJeMFogTYDNF7RMAfGWL+2bhM/PdFpy
Lc1S8d+Kl9z41g049IUzKa99g6+Z9aPqqX7EVSBvD8t/XBx73PmafMmVo2XT/d4v
nrSQNL2jB2r69D+eibfUJ41Akd3BIgtaF6YnUrPsave+ed8vlV7vZiU29wXcNutj
dAH6cmMfNciTUbNHsBaO79qXAcv7JI4XBC7Hhf6l3TISnV2FR5cfcVj8bjLItRmQ
ildn8nrHp3DGyMOF/NfeZkidqxa/PsTs5kGLDQZDP+cN9pAYGz4/hLx0cdo9hINa
v9p8XWKQDnycOsRYBRaOGwxbGFU2OPrXkV7gSmlQsPDyJQnp2Ho/U4K0JedAqnfH
56qXDjrbrePLSnba2MdEHY44Xw4xsnsjkCwQeDf5S2v68O1Hhs2xMPWPB2hi95tF
UtEOls6dlSBV9SofY9UAeLnwGhQhvfmLcT7ZpqiyJe3UwL5iAEULGUUqjwvVfTdX
foMSkcm1q82DfpU1NLDRU0F7b6sByigT2z5CKwX4b6HmNUT1C3YfjNIVCX85fIS4
sT/9C+VGcHNa8g+Nt7yJltF8SjXK72Dt+TxcGmJJh8W5EdxfDI2ZC9sHfQmDbNGs
C1f4M3oiC0iCk0sOWsGFuMAF7CiDS7AoEiMPrkc2tnaWiUSygFnczVBxq50TiNg1
47VFeBBfJXLheHTWwEz8AqMDoAsD1hsE6qfx5o183cylL6LjH7wFCy/VaYm8JYCm
tL76jYhToFVIWUsuUB2I/kkOMiPDu1oSjtBFps/q7vZZPhBWV/pS8prMbLyWnGwg
2OoCPk4ZUUNXMU/xJWywddcdyg+TWl/5+9RRhLycMhORlIy8K/kzXF95P4W6Tym8
gS5GQr7xlOowRC6c4+mXSiASfUpzW7ACNYaMx7VGSyft7ihxP+ISc2DevoimcPSY
dZN7lm/Asa7BNXRWLBVkF+rUVznYo0lfeE2c/OxWQb5FWMSceRt+KUMJpFunbXVg
QfZ7xR//tOMDlzFIEmPW1zwIjS6x1nnpTTM10ATm39qk839R3bLd0xn7o3ybuBn0
tTZgl9orxvoA2Mvudld1t3t2VO9jvLCkkiGe0N0tYnMUGG0FyUU62yvzm/cHV6o1
J5UNALjgieUx7ibzY+eyc5Ea7bxabd8sRc09WuI8/mkW56TN+Lah1YwP4RO4IMo3
P2AYs+yrYu61hcGHvVL4fo8Iubg9kH0Qnz2d3Lg5v73J4HFHyIsfWobTHFgUqzVd
AU9N4vGwjhqRgd0UaveqINfjgUAtNh4U1fpXiUFFY/cEubGNGNUzr9OkqG0daUnz
r2U0NUb1P9xkTGGZF4MFMMyu1GN2QOK52syHpKKn6aoszNRBrdgaiyB/rpivQatc
eAbV0TVkeKiItgW0lOpv4QxDX4ZRYRliTXLoHSqBV6yuhrjBkhjhHuPeHv331G2b
uShft99umS1c8XTSsEQKQo1Zv63JAZWhVreek56IH5T73dbQINVDyYIbVZKpXbZc
CW9he4NcERhGFB2LhkPaKOPUc+zBL/FmhXx2nm+aQNXJjvXv1Mt9S0JlozggEpWl
2v3cqoD8JsYCH6OlTo2caVUFP6BoV9T7IhPcX7ePiZpN6dYlo5aUeoa6UfTA5DVW
OpLr9Tw8hIdz+ob1dK9iQ6tKUWq0nFke55kjDf7wAQBA3VEGTzO2hUMJaYdfrG2a
VbdEsj4+vhnNIigS0cUjTV2qTC10QJoQUfuHfleTj3yM4hN2dKWztT3f2vhh2VB7
12IfeD+esvnleHdx2ir5v/rWRT9jlTZBreDmOmU4PdUYlEBPrcApe3lka2nu3DTo
qHEf+Xh6b6p/mmvFS3TPvhpSk/d9nXgERENIm89fhWXyYv3b7GTtRo+3goqTfgI2
Wzqvj59zr3DUYk8rEiAsYijn9kghY7VFOqSW+R/3VHuQ/ZYLBB9VNh7XJgFoBncJ
3pOL321dxJvnbE4H0LmA+gqwsxB7KqieE3lv5CbD1lrUpJTElWxrSCk4kSMxGbZm
9GS78JpPDiqHVLQxMaVmx4RZzoOdWiDz2kPxQsXZOBjw+X21BoTJOvZyLYLTZMnT
VGH3PhWPhPF9s3urmECz6ELWdcN8UuiMXETu7MljsEp0xkxs6K+mDoSnprrctd1H
tOC1CK0IVj2e5/viJHLb5GvmKTxMiWto3vWurZe94vKxcmSzvJA2FwipOqpSB22A
Njjz9jtLm8fZR8NGsws12SfZ0KediwXf6x+2kCQW4mHYwhlbtHrGtGj0UPK9Z3be
fsvCbzi3g2THMZxqp+SeDuKfZEE9wuiTOQx9OmpoJlSEzJy2ILIinC/vA02/7MBr
dpUgJmrj2M9mJcQNF09UYpUH4PiGZ6J+oT+TABCVY+qXBtoh4XM3BJp6vW+PXjbo
oA6dTPAWbPWUHOjwdYDWPkeBgdox6qO0nfdGFUPGZJdSkhV/L3OAjf45hz4NR7JD
AxyPynK6ogozWE6oFE29LhlqusNjMFdXwgXynd6S+0ghThK03sT8fGrsDklZxzhp
C/iBk6Up7T158Gtph2Llxrf51cojtYSDDrtHyGPv71jsM3DXS/sNAjNWiagJwh5O
rdwBeUtXO+58eUXNCy17C+9ziDdKw19DcWzAiGgxIq0xOXKkBt67xQVSlhOjPnAj
X5nZq7/qIU2itkuml20Jc3VG+ipTuw4pgXSUc4JS98ecFWrU9g0gKapV9CENEv5y
HgzEuNQucJD8mGF6hr+IynD2NdBi5XxBdDswsj6yJ0304a1K/irFDO7WucXDHp0V
hAGeUjw2lDT0TdI4sjV5W79c7TGwxPgerIisaU1FFoY0frCymfhK8VbsrOm/3upW
kyFvr/QIJehGdPwYOJnaDhpyub9klMEw6zjswEwmQ9Tu99Wy+EqwOg4cT8MPql2U
WbEuN/NFwk1YeR1GRPv5unjBA/0VNCQcSVWlViNFD5mLDjLKvTKPCIr5gxleuYCL
ervc9dLgvlGF4EycTebyj7YTL5iou+14DmkEL5MRIZkHarcfhMnpB+gbmW9sOmbk
lN/f/o4z+qAGMn0DudQVNNhBmVfsen81eYSmD9Y7uobEJcyAkJL5EJ+rS0gxXOOl
1r0X0ebJHQ/I+3aeg94OfusEqDV3Zs06cXFR1ZrMqimsy7UDi6YXap66vXCwiuHQ
iHrUJxpBh4rWIIOJl82P1psvfXPzrhS6kOLuQZFRAPX6YrMnjS9nDegueZE2+uGv
2bOFJ2yNypBmF1qkXKMcdHkbsbhr+Vk6BkovQdxbqF0xn7XxpTZA7nukSozOPqEl
sewhvDIivc77T76bFKC9IJv0T04EXt7Ootma7PoLcUIzB9JlPhWEfz2cEMYRvMKq
3sAIUUZ6L75s80aLFmbmspGtsJdfHi16L/3Gd5YJVw+3+O+JSGOTxfdLiCt+ftWe
6YqL2DH+iBF4Q2EdWn2ev6kx9T2Xep0QWg+MWigevhXEejU6NL27+MJyUWiABy+R
6lM0Fe2yM/4pHzAQYvSDLfQSN3Pmc5V36myU62JpFKurpkPofjfuiT0Z8PxcE1BT
AiuClWlRdLExr4X/Y2+Mw4G+6Ohw7gXVoMszvBEexoqbXulNOufAGQqfQ6ahpkcO
BKFW4hpoFp9U1nFdd67vwS5YE6vNhlFvQuJTrHcLaPGicutRKDM7zSLT+pp8lLj+
i4m36jf61Ya5pbb6zKh/NhfJZ0d/VRuCIqRoRQa8B4qRADy7G1avWbSPsHcggn1L
l5VNPrx7d1BHO+EBnHz47V8+cyulKy2aqLyUNR5gG96nVImJmSUHd6/ROP+qCXq0
OBT7BabtdQ6WpmWXwVv0Z5X/BBTJULsMora/zYpu1pE1MXgoMD9oKUjzLTgVAGxF
a7YosA0JAJnC7JI6M8lty9nZArBohMcW4XQYh4ZFBc4l6PczFWcAvjSvHybARMsn
bjrkdM5V8EMGJZisinuE7AoQ0QPshWu4vyDKSyysoFm1zwFCfFMlrWpRL+j1blcG
ZTja06hYL9POa4sbNjo2sMs0euU8vBLLxKd1wuHF/Olq6CKT3p/iwsIC+BPiK2G8
yTDaflos6AU5lAhdkN2nycAIWRDkFqAq34qHjrL+OhKjURn1Jc5UQW7e7TSLa8xp
svs69RYYO3FriIhhr1+urFGodk6pkKroLa6v96W9N8YP9xNoEUggvENtfhxYFTzY
WhErxn5rnm8CXA9Q5mtKNxANWyQK0DrDmcf9GDxZ84DmEbDspXuYXMehdVLAxss1
h+9PE3rha6+U+Fzj3hK5yWKBIx54yDCUklYuPUYkW1MsGVoB2GI8pc4JZyj7e3IL
x0/GD737z2vWMHCBp7brFu2h0XcTiLSkEdOQgPQDlp6MQXCpAZyZS96ioBQP3V+Y
iQqUblI2VCKddtns10Dwomq6gwkNb1RBazc283VVIR8xtttXmnRk+fg4uE0HCsax
ffX/JLh5gyS+nO4KYc2uLTUyVFpXYWsnKPkJJVC8HuW14iQLP8UmkGHRnMSvi1ya
LH/UtCJS1SYyR6dIQ8rRNWvTYlY1fbJDXNfJstUceGIFh0p/tHAGyBquckgeTNsN
VWRqk8Ojee/xypWlLwkZESgVg5FWNu053Hhi/QAW4ZVO9bYUn7qWAO5mPbY0HXUu
k/1CsuYAhmEQPe2MdIf8pCdS9BxrR5rjxiclheoO8bp6IISBq7gmA4kt6s1JDnr2
gAP3q+nQtp/PczRsFYHyK8OJzX1xIhUuyoPxKSciday8xJbS82vL8ykKeyADsmVt
pyU2tAwPACzVsJ2y0ukyvnmujQ7cvtuse83WliRl/8YxpT0w2b0SUDv0UvYZ8VD2
0VZPaVl6LNWDpEjDhYd5Bkeq6x2iqapdDFxLCpr9GAulIA9++QbgcpHRBcmhFQwX
5Yt5UULZgvcBI2XufO7VObYG3GqQeCrLgxVGeR4km6nsvvZMOIdvzypTdxrIwSBP
cMOWfb8po5JvLsA7/kNR9axkA771edLLamRa3/JfiqjVTiBeddMV4BNcZJ+SDkgV
GHvay477WH05E1IydpVOxZpCqE4eWTYgvwXGTAzVMZW7hyjX7W1+uRhZ8YBos59o
ZjVwlDK9T+aCaCiDa+0SAqlMU698G3qyfJDhGg6odKA7jZluDEq+E/e/dca23RPP
Zu+5Oa8Wqoc2aIcPbAlgnM/GvrBZsOZPxdj2LHsDUKnl/1MINwDQCFHsgAB8WRzS
djm4al7S+wzPaRet3gWWGDutBpi+Jth0rd2ACGCiLWQsy/YOfUvfF1+mgJThHV8R
J3vQiMiEF39/j1tCX2ZD0Zr9CQAj6mtido4enXW/3Fd63eLViKWEav59rtjPLs8f
ZAgC6IFj2NaB4wKsCNAlZCzKDX6B+ftc/e2T3lIHT7eVuSBvgqNB0awPoIc48tMH
fS5d+ongUnzSns7xpO9w4ZeTz81ZDRVtXtkt1ymkounm5ANyxl0fxO4ZNbwLoUhy
IAcbrrsVPXGsXqEzIpSPjB8s6hVxChlMaZQludw0/hbDLbPR5oXoWPgnEJ7w8Jik
oRamUqe+G47ihL9aiylU5+X+cE9N4rXARoqjdQiYNxMTtY4HYlnfzfBsbJz+ezsI
SBJ5SvNW+m2ICPBnrRhWhDotRSG2zSv3zqOs606xJy7wAswiuQXFaXcPlhYew51Q
jlYnQQFuzL32BPlBFsDnSdovx+pkle9HCUPRvasmKWH3CQze1Q12dzihClC7vdFq
i/NwszZ3ZTT4lT+0ys/7ScCChEqHxXbZhdu23XujKVuLGwi25VzZ9/oszelLLPnB
OIRzLTRXiNy51VR9S/tUhBU93WAVm87vfcSTwxKXPzFQHPqmTbHF+irDrDzjYSkZ
CfKyW42obRgC0KkjX69noKJ54r6Em+hSZ3u3f4fpfI9EijOUndVrHgO5bJXVSv8H
MjvHr2ekSCobzibycYXf8LxnmwqgCE93l5YPq5tZ1CHBSAWcYwGb7GWSH3gzBFre
WKr5WxhQNbgMIFT5SAv3ddr21IaMqQ5/4n8DW+jE7RJjY6azv5xNfKe0B+Em1WbY
O8h2fWTHcW+QHvGpV87DuUg9WISA+qX9o730YowwTFlEIhazEgCVUAdQmznaLfUk
TglH0fBlcaDB3w9uVUDA+IMRYV7d+H8OQQ7KxuZEWS+nNexSy7trXsq8x8lPL2aK
jkUKvaVGEStUEnaLGFSJjIX5U3jtpXgqKDr9N+VNoe5Q+tOxGfnDDdcFLiUYsUTe
5z55aA8DMpLZcymnhz/LYWeD/2toBFqYkc24fwUDqnTTLZQ7EhTO5Cx1ZwJGZq6/
W8sHE40bEhg/vYzxx1jPuTXcx/PZgRzP00Vquz/dkqkr6o7bOzBkuOG+0HrroFZS
fiFW1aviLhD7rwj807m+HaZWWugOwkEtqybjOSxfdcg6TKzb7PBe6kvzBxPV9AjL
cDoTmRaRnt615k6c8UzhkUX5ClxCJi/tAalg0l2lX+RQaw/DHEUpaL0y/AdF3nxp
Qy5FPTACcuE/0n1OU7Cm8fHsJBIS0T0yxhYsGQ81gKSPvzHrg93D01zpHOw/n8ti
9hPsqSHIILnoSsYxXGD4Ioki7rYaddqnl6h3fSaS+B0oaXsw/q97Ov1j9PBkMkcc
jEGIW2113c5lPC1dbSeAucvFkemakfw/D/6wVTICYS0SGdQ0pXYn6NcZ4U+kZzet
d6H69ix7edhS8cw2el7PAASSIbMVvihpmlp5r5xWHqH5ZRo/fgz8VMSz9b0Tul3o
UGQWoEIoX5Mdd+defyUhvodAWFgq6+e+wW5ymJ6ysC0qHis6WP+5nU7diMrIdi3z
v2+bhPl8HGNupqAgkXywBu8M75FfaU4kOtRlEFLs7ctPtKR9NcfIT8wwuwqYrFof
EQOA8Z51lE4yehqZ6Ho05If+MZpabFoxb6qZlcBxKrYkHuvEzKjftzBKsB0B261S
+NvevLzTOxfX5ep3ctQjBgJz0R0PduDLTAnysDrfnSMVOvlHy0TkNwhAR5z/XqZL
DZyFJ779rDD542q51C1+qkuJ+ZgQYFhzUSMFNUtOPm72KKo9zyOAsQavJ/sCJVbs
prWDleJeQLrw5ohGvYI71XvUdYezEI/cO3BbSn8ReJucXVChKo+3Puw9QtOZ9bNL
TLVBhzhJWajNIpAFV6EDgSGICqbKzxm8Qo0Mt4o58zEy/Vg+/CPnCippx8NlI0Y2
zjTPml8nNU4erW7UD0P8bdmqlufRCblBTjgp+ubVO57BaE0B1iKZna8F/RtXqCs2
BKOmkZKKxJJGzrvFFdL347NTizRSz2/1Pbf4aqlDx3OYf5y5aMh9uSHq06M4YLs+
UpHldso9CdXFlEBaKiqZYQuC4yhr3d+YpDRrrjOQAsxGO8uf1ecNc9TAYAeX7W3q
IF4c0a/7ZyfYLOdQULq3Rj/k3iT/eMy2PDJuBLHP3NzqXtcECDqjGcUa9PB4zd/Y
x5EAMAwvphomK3qeXih6uMv0IEOIquWuogKwRbHNDimng11K6DuqalJrW9TC3i+n
xNnvs+fjVTkdIvuFKWqhs+duYEUEW0Kh5rHp/uaMQ4Tn52E68AuwAwttO3gD92lF
zlsjEJbwD6ePt8BVMnoBKJsOvryvguPggFrwjpkPPhArVLjf3DsyyLOw+/spGCLS
NbDB2+f9zbEA7fkMlib7GTLHnoYZk7cGbvZMhT//wtAKK2oH690eC5QhwoUVScnQ
A5ZXPkCDbB/N5YAToPyUC/vRhP/abiHv86e0B29ZGiAYNlMTUBgGdjezw++OOIuz
ya2NMcsWop63F5xzZigze4VQSosQWbziwex6s5jGjKo8a7Y2Yn3SliI4RRuS2gTW
j2GmEWeXgdbISzhDftPC9D0yRbyjYdtnvhufchHgWGweV4rDgHFHgUEs5PJhWYJF
kPlPJsY1QBSIDmnhT4wLwjN6uQiijuuurzvuHOboLnW3tzx2Sk0aySmxSkRnG+tU
PeYkOyWren71pMZ3QQswtSlQcFG4eCdeJQqoLeV+Xn/P8swjmwoH50vBRD+iwYCA
8tzeb4xFi7F0ymgh/16WhBUACqOGxruHES7Sa92V1een92SyX+8cKtizWNjylnXd
JDCRDDfhgaA787DtyUdZcduzf9Zm1wQ3xPFZoM4F0R9Mj+efHN+pFJkQ2sXJCI9x
dkMT4/nVGL9nm1EXoJ3/IAYTsQ+TbAJoqV4NJHM6HEleCxSaKjUvUPn6ONk+7rmb
jo3NcxqQfToC+zIOXz6nPQMhuZ5fgFGAShuQZB0yxnw846vNDqKvNIi2U/CPF4VY
OjmMzKiL0jdZifYctv5AbTVjoApoqeCV1FvouKaKYVLoW0pH9du+JEEBJlCVtmeH
9ytxrPiZDL0UL7b2wgryhzH/1AQ8L5C/gvnGoFe9jt+30mRaCfLCR0ZvtxaM25rt
RPS4Aj+aW6PkdxAQk8RBA3yCdSz2Nr6odfiHiP5OehkdjUcXSpVDzD2ShNLEILTo
cR7ubRIwTa66Ni2M1/ioIhCTFM6P/FJXcFtnt0x9vsJ+1pr+DawjPckBuV0ELu6d
JJkL9wGVYl1zbdhoiGuFoQJ12gt5N6/47X6UQ5D2IpYb7pWmtRqs8R99Wed5ofaY
2LlhZhbeWxV1nKhjF81oZrrJGTKKLyOWR2qZy088I9pu3mGe6DZZALaTevqYfgNb
2N1RxTM24bkkegtOhHjKhmgqWl7rMXbEm9S3Il8zgRQ+QiXRArHoU3173P82PP+s
kp3QBiB21rS7lTPKpWvnLH3p4VT1uPOT2NWvMtG8aKyXXwhd9veI6NMzSDLB1/mm
1JxdFexG/fxJW5WS1qepykCTJxv2bzg9Mrex5WL44y1Xuo7mXZw5bysgNN4zqmQi
IN7ixpFl9egxnpFz4N1BDOxPLTwZOyDW1ZmjIC0wYo/L5NdE7ZUeDphzA0mh6nmO
Rw9UHjip/ky4wwBFpZEt4xfqvN0sW4robK1RANVwl6IgLyRYFZytIaSYAWIYIN6Z
vEOqFpNOj2Dr3NpMBgEgFNgdvkzBb8Audv1GUohfdJkX+neMuGaAMfRa7Fdv4Cjp
pT6D02kqFvMqGpicZaJHZSaBbKEIL8TSA0QhXIPuI5OFi5KTZrHEpaa5Un92vL4w
0O7EaIEdoksbsFC7arxPz2Gj0e4VHBG5/+stDQjOA05Sf78T0CFwLalw5hj+1F/Y
EHk6w3iIyTX8Q2bIhMexD5NpftvDRTaa3kPwfMFEhQyACXntf9a281go4sKhFpOl
oOfXx/BELSx4dHJ0Ne2ORQqmR8/MtQKpStMtIWvVLIbxbuelxrOKf9z6B5frQ5Af
1ANM4Kc0LKzb0MBCVCExkcgAaIPGbOipjJCirkwBKlyH2tuXTrJec9m+0cUWto7A
d7NHniZsxKskj+1CG+0NTnH6nPo85ERTus+kTNzKyCJvtwuaisIoHiijo+fExHZw
NUHV4A/qodwtwn9bhILMhjvGrbnBwQaOoRUPCccAYgF8R6O7I23+T0xJBfLD5qPh
Xc7I464YnX9MfjeARx54dTcaVzr3Ig+QzEwWTw99BqbKFOJXOjPJrFj4k4JfqXSY
N6y5m4jqRJVhtrGuNC0WkKoPnWkVj6GbHnaFsgz6cFlmEyPVBmcGSbZNpt+yYwL3
5kHPWrYxzSYP/1scb9SSuCNurPbF6D6Id6cZPj2CPNmbZilc9Qm2vEZz4hCjjfwF
s11un/l9iazXpl2vLYOXxVkv5dfEH1ffXclNkPtOEziRYRQQ1cgXOnYygOp2jdRT
KoUY0bTCVsZckBRmWwtclS3kZmQVnYM8yHnqEtY9/3a6VeaPJqWLdBxCBEmSVYM7
Av5u8JWajyC//0gaXhqhRm0U91eK+GVeeKdmiFOLGDRNypRInzsvkzelTEWy8ctr
4b4p8QOVulZzH1sMl3G40BBTZ5hOBsgflGZEU0yt20wHw2pZqS1bcvK+tuOmg+VI
I1wXG+S74L74MTSa6U3yAKXc5+VXTxsU337es+tKsFFPwtsMin80poyC0qYjXY8N
QqTNNNWdebZn8dbDRQ/YxEopZjK18utO9iBmIkxG0VCsuH8mteKr2aO+9dEtG8TA
sx9QlxHVI1uysT10W2eLIjQai/hPUVW1ap2WRQtHKLpt9R5rJ1nw1MvrgCiZHQY8
4Az9CZZC5k6aW9fcxRw194Y1njmjXO3Keo5xk96cMgey3QctU989wjTN56Wzodn7
+PUNaZaiXq5vuJrqDG+bHG04Uvr4l6lDNYq+qpBObj4a7hIfDXTxs8prMYExEPcA
G8dhFomuyQ0E0eXupT2E4WpPLO3w6oIP68U2nsdrg71pbXS7S7u94GNKbGzz2VKx
EYkh7EEFbsov0myVuvLDwNh7Ef/VyqXnhQPmm7/gF6q9kn5XQJ4owewCzT3xO/+M
1615SFWtMJxmxsyrCi+Xg9g0ULHlRmLRN1x4/2M0Ccn0+OHFoPpunEzW1t25M4XD
BqePJnPAzJLx9giyP1l7BU83fIocX/UUd395ybyxX+9lFiVysoEqfm761TM79Wfn
SNWunHwZZE2yywaBKvV6Z0dknN1hW1tnEZtTsAACBBHDFPtyswC1I4bQxlb1symu
RZrNVykYcUyCUlAmHHZLw+fbzJYdovjx7+IVyohpMc4b8RnX9CdElHo2NSlUg7vw
ivjLsQUDuw3UOO4OONgpNwQbi1S7AhQS7k0AaJN6vM+FVTlFrF0a7MtTIucOplpz
DJeTARXwH95HguCEwGBA799QQOb6z12uyMszbuKrby6ZTHvpeUSbuxATooZhgI+m
EtzMaxBFC6N33SHGu29H650LPwK/FKSnYd8wVNR0f8OmWFHVM2fkJ5P16qENf3TD
zSTOkMwSGYyn+VmnmKDhvGvYGuxeZkPCt+7tH24OhkxpAQ2uKQ7Ki4UG41xkwGYl
FrzPKmJq7UEESjKK8LS31MHdRTOnUW6cgIVSWi1KOzdjb0VBDMMsDL8HvRtzmvI9
E8TjSJ6p/pfY8ULTJEm14j3q2TmI7QdrhUsl1BFTiIy17jEI8BQgCUpYiJECrGXz
OgyO15LpDlZKn+J3ZMbXujRjKGvAy/xet0IpPLLitBumxefMGdxOQlAQsoteW3+i
zEVK9gxsDKannO5+aDPMm0JfI9kny7jC6U34JlRVsiS4J5CODXY4AMpmAokkfzOD
FP0g7x+n5cIIeKU5fMWrbPr0NM9bayFl0xnuziLLCbl2wHx9+8b9m7dw/tl0cp24
dbqhrUftUi7bMGxBDqKzhiD4yjP1kJs7A8tkUezteS7AQrUD0wuiDSzEbMcGjrOO
xTgZyl/nZJo27x8+jhH3Inq6pGLQ/eK06Jq8v3/hw3bpdTmxJ9/VXRms38wst3QY
/2zyY13IhIO+IetVLAedWo/Hw/VvmAksWhG6hCuadk2SWRoAGI+J1zZidKDZiE/f
qLXntBBig9cGI6PRIri4SLiDxiflib4Aj/6wa7QJ9hSAfIFDdxyWTGz7tJTJZVq6
WWTjhoWscBsbDB3KlGvwC8rA9tRQmiapSFcxGCUxbNLxkUN6/YU+0jhF+uZWKmPi
edrfO8ztBoCA7BQrEXwEMpYAkyCGZVxfAYa3nYcD5lSKFTB8dkQLQJiGkEXbo5nq
t+xLqzoud0Cyn3v0AsJNrNtlCqL1T0RFrUPjD2TV3Rms7ZgXXelEvagvIyS3/csA
BQOAM2tfeAE6jtRIhJaG4HzdIUfPscefwv85/EDORy+KIGdO1ucGQERTmWDl+oxf
VuceRclaRz2B/KP83zoOT/YunFnmyKMoAO522wTmPXw5L/2ws0MMFSFrC0vbxA0l
M1iRWHJczkzrG47TCUgxX6zL37p2IHr5vJT76VulM5EuywKM2G3PDeq8AyZNYLR4
j3H1d+L+KYwtBZInlp++Enoquc5AzU4ybvoPMVw7IqkBpq+iu9jMwQPGv0mDi2hQ
hFFNdex4t9kVP2eKqzyd1RZM0exVLUPJVUMTwqAbom1VDFy7taXNF6DpEIkrR4yA
NO2hD3kLsqOmTkhymooxOHHxaMuhWKGr4JBX2oEMjtGqnb5yz74CRHOrxKtnmNen
KVKn5aE/K2i1Npuea2kKX8SJk98lEgEVF/pa86vvwgOMYl+3iFqqfMLgoCkzI92R
v+jyKuUrS/ghYx5NrJ3w1gZrGCci1w7JIAmB5zn4StrmX87Dg6+/J5vAS9YLNHY7
h3pNQ3j6V6KZk4SJgEbfHYjkHY2vz+AsF7chgqtIkzCMrRRcw+mNxclXdgSdnYVF
i2YCeHhMdmIG7HQ12u/HkXObZ28yrJBdH/SNKwLxvZiO8ZZ7GdJngPshzEc3dZ2a
MYX83FkmWHsc4+YJfnEEZRKqf0toQZQTA5Xolt9xAfEDYbEwmbLA6bowUdo4BrW0
q8sP2if6I09HFs3S/gsju5vDVr3W52W2Gt0u/gfE+x4B97jhSt+ejzrNoVJsH9/Z
CIV9AqHKfb0U52j4sA2yHYMAZ1YINXEAP7ZsJcMWU6kwf0JWhgNK+Ib8lNIC63wt
ijk1lo9HIoDm4ariMpIvF7mBD9WdxOF0T+i4N4/OwhhMYymW31Dg8NbtUtCHU4P3
74LJjute7An/1+Vx1PgDuCzxu/WxR4yQQE7LQ8b1gQPv0NBN4j2VR41zbIjLem0x
CDXIlLtWXgni6/soH0fpIOlQRpaiRI57OteshVaYZWbBttXpweLOOwnZwZeitPaE
Q//i+6MfL3TTsMolp2RS/G7LUhTtr8oWimuykrt/QqhYdoas0geoEiPWduXylTUC
LrmT1hvGx5PHltBi7rWVuqnQ4VBqDtv2AfjJxHNWxZKWoh7J2DmisZCPKRbHJ4Wz
7Ca48dNDNWF02HJyIMaRBRXAXEqoEAtIOXLoWItil0yXM/byE56MqIfHaIaLxwQx
bG7xpEba+chsgWCQ2xuMHhdE4qXj81hI+iTQgIJnvp1EojUEC6IOVyACjriWvaig
wcDIpv1d8Lo/7amQPyGZARMMnSftU3ZIm+UmEO968ln2DgBqjI496gRwRNYys190
sKoHcA1eFKyEwTJm+2vEmVLOTTZNwpZ6Jq/qBpYso82zOR2XZtuUT9TLDsrMaKal
q5cTmtC781rRhyGitoYeMf7SRQXc2xqqdhkwDB2/huzE7XKKNp8redUZKJ8gP+6T
iNosV9ZhAFouUdHWFc9LfreS2SdFwjOi8Tso+ShuCRjT6a7QbY2hIr/tWATToSv0
4OQ/2nCxlfiw1s9TEcSu+tt0rGl+cp3pOhrEPQf7ftPqCqmd1XI54OoBcAt5wk2U
hX8D/KhtIW0wOOQRjRRqfmIFk6wff8zpJ8IV0xweR+bEqtaYWbmYQqdGVlzel6Fa
UZCI1bb6LKbALbhlNUQes6H0anTI5bH/BCq5tjht2Ru1hiMGgcDUjIgCSs2GA2Js
V51OcJ0HAomhuRcbhDKNqwAWk2t0JuFEDNb3naLYCIpD8wv9CPuTsjYi5zWVJhWx
auqYabKWwNfagRgwtRM8UUTDFpRly0tFP+LYVdv5+TXXuyCSqyMpOSGq6DOC6BSn
XqCjxYRgjODNucHL3kPekCnQwyer63y+kcYi8aDjoFkHlRD6i9g4dBBUIFYHs7yc
/NznTpXSa81kYvmsfh2myMoo1cp4jngpUwau+hVOJ6gRCBu8Mm4u/Zq5OKwZ8Iwl
FQJwfA1poeQYhWZwmdMOUCJI4UmrfZSMK+P4jI5d6SK70DifrIejDa/M4pP7Jc8L
ZrjiYcQ2Z8KINSAvfOc1Y33n9OfENy992Ajk8XNMf2qdxaJMPZ9J4hHEwKFwd/Rs
/GmNe3i7tYP/saSlL4N7JRwobprJzkSqPgAelR53P3cS5U4kmeM1u2OWx86mDDlF
KicuO2CPKKXCSch07jSYE4EKunV20/FisE4Yli8rfiEsLxMuJAVp4nlzfZMBBDYC
6OVVEvKV9A79RlBG5uezAQHb/cbbjGoUVT2yJuo7UP/S4rTOffp4VSXMAyPscwr2
DCxBupDM8susu7Qb9L9dkpDe5PNdYyhtCYB8Z/iH4FUnvMttAvbAIQtD/An1Zm6n
wYFWejwZH0d4hQL8PIhziF4hB1QuAw0dhLOf8hJjRZILCNvG9h2WIV300sOJaj/s
Wsv/5kHP6GKigRUL55lc3UeuED43O+mYe6az51A+37E9DQB5Rg4I/Qq1sbN7m19I
2Tw7U2bJsF0wItzLlokH4S9gnAbSuklIR/Jxtg0wawqbTIS+nqBt6O4d9458CMKn
c6hv56iRhJONRMvaPRdNFvNqyAjAA05qc+D8cy2VnEEA9wag015Kka1oIx0Ayp5p
llA+ch9uB8St7iTKfvbj6bw6L2NHUsLNyELR8LhS7rnwMN0wNx3fgzZDKHRh0wc7
xh7r5od27maA7enAVI/7y7ZuzAMkg/LQkstEIV3OCrnIy3OqObAIbrr2UNLCxICM
ERU/p5y4c1JNi39cwJEzwz1QIOfS1HBcQAxhifpygt/qcQsWGD94nj6kQ+AGk3If
a9CtZAG6ZZxFoGuouKYh6JwBlY2eVJWo8BqJ66g0YlQrOTAzQZYgiD6jxz/tQUWW
SHVk3i4p60ymQgf6TrNdAo4z/CW0Uef7qLZrV8hEzJtCTgPxqAq2SwvKCUBDf1CG
NTPWRUehva43n3bi/uvfgI/7ho6UA6UhazBYfmjcQpgQTPja797ptKr7Er5WH5AS
iqBjIMpb35YPN7lEm0/uHXUdkJ72GquYFEYLZBnnkYInXHx/4j/JY4wydvSEYVmO
gk12/2IqJIdgs4dw9pA1+lItpRTvrlSVh9aCHK3wPIIc5YTLJVkpyMpjtG+r6opp
B4zDPKKir+ZRcnnxXx3jW5dp+wV+SkGCYPKi+70jZ0EtZX2pHk6IgQtAkXKtMpZ4
9YH3mYDzcHQYtv80BmoSzBmjl1BLw7isttMXkOCR15a5hVH9WTwCc3+rpfKN0WRE
DP29ION4yaw+DkrewdyXGpLrTnIWsgAhYjvqIe5IyLPygUnAvSAHCmQiebf3dRYC
sTSbccLZJwWiIphbeeLvW8IZ+fbnrEdGU1H05HZGofWEFXi6MPgCuduj/J/8Uziq
wXQzUXVpnvwEsHOWb3mlVWqwZgs4GQPGxJTS3/U3wDmWXfg9WBazqgukouDsF8u3
EtO937BsarP4FzGJBRavEgCM/HJDhZzL2r6vc3xhslGIB76XQus26m40Qvf3ARCT
T0+PUTO6OnXgqm1+Clpj+Z7CabWjb+5nDx9b7GpI7Kj91TbzPxRMaEr3ZPo3zmT4
NjZq4sqy+m+VIA8mMN7p+mwK7MrZr84eKMl6jShLmmgXmZoPtpkWsZ4fHu242qUv
6f5SBzFCBhj0ZqJKo+szW+7qhFsHYJ/yHqVDjmuriycxizz/5Wren6cT+8NyhpKt
3DOrWpc0gvGnNeVt3Xm2cSMkPlXDnSyFzjGPgSnwUqP5S9MeOVXy8R+1nUnWyBYr
D+RDBHKrabP3x87IqrJey7m4qrW42xP/E7bpTyCT09QM9HnofyKUQrkZ+yJLCWrB
kTtaLYZy2NmeI+gPaNd1SZZ94bsQOUpEZYxjLVHFaDRUaXZDjEmSERDuJIUrFIQG
7VxEsVhf68ItQBNPrzI/QNnwbrtX6y8vhxH1f1Gu7T/fZF5o9/mZOjcLO1MZWycE
nzsqGK89is6hIqotpoQfOSjlCvZnGmrJDiNh0DC/79YTBfRcFSJi973/Wuf4YZR5
AOYqfDbsWrTVoC1Ps+i+NGLPNyI8qEDw6feJt75AuSq1j6WzQ4GrTfrLB4kDBga/
ZwaAK0mUPAW4M27UVPtxhOguh/Bbh9oEhqK7L6y78GlnWL8Bfw4JucQib3kxdliQ
mnuKCJHVryHT6UQrhrMHI2xCM3Y//m1cDK6Bvxg9bVh9dAPJ4tMu+y9izh0MuP5X
KVb+4WojX9h4sTn4GW4faUwfcrUb0WJqPV0LQqIdQrE6auGP51WaQPOBZt0oBdKH
Zr0waoSu/BxUkrZkLe1kRdVBRkvePFb7Hn+E5Quy0fSqb8Pvvz99O+qCa9xLL+wD
8xLeqdZL83p0M1Lbx51+AuFsFyS0u4WTy8rvtr7tK/RuTkl79DHwHU0J8MCVgjdD
KrureKCXncsrgqiRuvaX4LZcWS8Kww6crAX6GndjDdooXvDituAF/G0CxqwkBu3K
M1pm6UIdSDUl0xht8RuWJFJ2FGg33BIANnFWisSA6J4WRNgiePxf4d9VVK9z4t8Q
egU6n+EsYtWW2bMKa7a05k7ul5DuMs1QCkAWketf8fWrJQwWiPYaV1b/wpIyNB8F
gl+RAenC1/hdQMdXCX0bpSRMHtV9Ovw+2w4lGMgYdOXiNLwXmyYG5IBgE2DUYOxg
x9ybqVsBwsG4eR+4fqdTgpQz9SGb7IQrBHeOjSYZGhcQXyEkOYRpX/vLGj81yENO
bsGnTzx90ofDZh7dOdReKTFBAUsfpzl9jk1UonfOq7qE/72UmbBpPD1/bAE0Ewom
f/z6MXOXpEis8lMpvG71TwzyqoRCl90qiXIChlYhVUcLi96bVdyQPio0IhaVhBhv
YVxbwzv7GRenWKiUoDxICiS22DW0xDE5HEwtBmdrTWO4D7/CeGdlqfb8WzaCQP8z
Dne1odAlGjTTxNMuYoDjw58Grnh/p1Md4UxdW00DhYQ4nDl6Jm9yFms76Id8h/Dp
bmGLYgbO10H2QBZ53Co7AwxjFv3Z2LkxTyPKx6sgTIgnKhT8tAPCxn//ETlzsrAX
kFJ3iJq/3GwPAfjAYyk5p2W1SqKXqbQvlpnzEVdVzYujbNhnCYDwM4Dvcx2q+7+O
UBFXMYD0pIF1F0Y8hkTVfk7fgRBdyn1HU/vKh9CzkCRFPxP5Awd+OrsGJRyVoIzp
yMLUPL5YkckgkmOxpJSaJ07/jXO15OW8aQoqy3wfeY1dMZajYIsB1AjX9RdGQfFD
ihVFBH+oL/fiu/VxiwcYzVvZA37LLEgBoabZg5L7EjbncylF+aVAFEik2G2/Oo5M
+tg9VrqKPJDoN6g00Avr13Dpdzd5fTe3+3X+xcRGjZ/0tGjxNA4roXDpAKE3+1oD
GgulQYXe/8IdgAcgsGzS0uI68Way9blWdqvlD7Lcod4KS42PVKIs2JzuLvcXJ/tM
PNvYPJf12pjSWfz6yQ9vNiKagcCZG77bAqT8tTlwD5xhdPucdU9eLfyR7+eKhoIM
Y2hnmLiGiD/FmU81f5/fprUAZhg45q9Q2IwMKfvkavz86fgWul4mFoRLmziUpkU0
z0Zr/H+eUApuDq0n7kcR+59UrNf1AKU61f2nU6kWa7sLPyBQa1xwxm4aWUPkDLmN
eJT5iJRdHh1A73cd1EgfLXuvPCe7UVfCjIxwM/COI1ul6ALFaWOD4zZKPRUhB/zR
k+lw5HqYWG4jI1jdmw9MTmhu1UGkqPw5RjVIWkKg+tCr5q3z4ibIkzc8PfzWEH9V
QYYfE4d6ltX5HniDN1e3J8OnK0yElgNtrl0G/owiOCXtMY8gFgtZxHyIGbhotzPW
Di94UeOwBKRwfqoJJkT7mKAF1DuYybxFrNG/XyQ24dGV+zQs4Jw1ppBtnNBGN0Xj
mLJYQC0CTyrkFU9v/ar1vZDKOHkhwCbaaQmB/SWBIOngDVpNNdj0xZ7oafU353Dg
kRrOnM8OB1LRV1HcvfrCl2lim24A1p3rvVijsQiet8riFO+ifjldOP/FkG0wU+w/
BwXOOlzFbj61JlOM8yNGXH3tMp7OCya20LbscVp3c4SsE+7eLN6ZwTA7Bb2jzl2M
QW6gMnpeIunqwSFhLtU9TQ58l/jew6lzcLIvWoSDKXZbEZi3Nk/MxhNYhgX0xMGA
7pBmafEIIc2nLwkpTgX8yt/Y2nCoKCVmOkIW+01SuZF3XNhpbovhzbXVxmswJ2x9
rU6jArwHBSluNFv3GmS1shUCfB36W5b2YrvTgpfG51/Kj/l8DnMFzvMj629/jjAO
b/9D6KOatRvTyhNAN0Xk6HPOX6b41xA2yR7cKt7sTyJdd8dGVk0vxeDJ/oZMbWV/
4qlqa1ozQw/olCY6KsmctaNURzf9VfRRhRdDX8J8I+uIPaLhGwMJMiGtX+IUVgZ8
YzhFTsLYulUjIFWNyThtF9z9niQLXAWf/rR3MTDBza6KSRnPFIQce3AluLne8YkC
iYviqmd6YhJstwTAtd23TRiV4U+/RzNo5GkU8j61mPUn2OPIuupS2+zsF+7dGtAF
UJvXsEAzzl8xgrufz4xf7GDzz8qpUeD9FpxYr5+FR/9R94lJxOXnMoLwc/ogtikF
Ytf0TZXDbc+c7chBci3R3eJPX5LHvrzH3JTMShdiby45qGcd/li3knEC6QnbVONn
NvcnrdIm2JoNFfVK7bBRrWS4dfoUNAsdTMO6AxxabZwXPwpupGTwWAjA9okGWsXT
MFWhw/gQwTlAYme49pt10qiRrA77vp9ltp1gdYs2k+2uFkrkQ4eK1h+pQ77ASsnS
nYJRXEZA3q40PNY47bVs4kGTdB4BnbwgGix28ObcNtfousSJLKVn8rTEjNGpgEOM
9lyicsNFGyUrAsMpXqqwZm6UKkXxm0Vx/mnyGPB02zK6nhpIChVoIpTSJyi8cJEX
/s1Gi/+6lBQQHGwKviReidm29ldxNp8KwyeCTkj8vHvQ1s1BzlLzXOE3FmEQlR/J
Wn2GtqzNwQXHZdFNQ7nETw8NuDNJYjQdf9ev1Sn2uVRAomFFPDXuCnKUZ5Cv+1W/
M3/S6WuuQsBxb/GUhGRhVQgpvfUK2S0uG11exy4U9YvyVdcf8MfEDbIMk1FfLx8a
5HVm5EpSeM7g7VCBq2vmZucPKKwgNKN4QLc4CaZeiR4YrZvoN3PG8HCtASa51MxM
aNqR+ICGsC6ztblW3KIb3D5blfP2T3Mzid6+bFPZZlsRovl+NVmhxto0xpXxcSnp
D5XgisSfc9jKn5NZWnabNhTKl8qJ/MqAWcXfO46cMy/9XPJE9MpQPqmNYgpnz/DW
qkRROQG29zB0CFo2yC7pAcQ24cOUbzqjR6KuCjYIFCMpRgqBYY0mdvVmW6B1P7pM
BpbWrNaIqsAnMducWAx1Lzjm/PD9O5VWiky1lyvLAQJpyxOZWNCWvT3FEQ5AV4iY
5hD5UaCks6+EMLgzSfc96UkEEd40DeX9TywJG0qEQdVTodQkCybZ1nLA/KqaZ991
6bs7Y3b3gIBkf+xtcr1Jufr+0KPNX7spSqwB66MejHX3H/1B54BCG6vx7pH4yZVr
LUzWUNQNIMRlmXdnrvD60N51Ia0E1eHkE7LKmptaa2TvjVkZBSFObNrKZWFpNoz0
Nryv065hHyu4uU5Zp1B/Eq7nqf0EBaaRxLaIQH6H+72Iy5YOqa3vsFrxgnXOyfwH
xgiRzEaTJMc+6NeodKkARLNLAFGM0zIVgFvaZXNUeiSlS6QYs/cGKWuK9Fb1ILVb
4KoOd48J9bK7Ri7/tz8gZioBPcVbgFh3/dqkwyvnPK4cXRagIZEs4DvJn3n2Px2t
hD/5aWhYK816me5f/pnJGgaECTPbDnR94H7qfRFam1dkeAvtKJ0KxesoWvuS2kWW
T2VCQjbHAZY1llFBC0MrIiPN8+uiMXPgU+zSIu3jFFV5I6polKHWQslMkw66BkMn
O+6uT3jG5nLu37drfiYDkCH5sqIVAoECIsmnSGqHEwjUjFnGC5hUWabDuk0ovW/0
0UrCAkzkerzgn/fZ5r78fwUvFYoakZ7UlU0+a2e6UPUPhtMKGfcA6/0E+P+sX9I4
Nu9vrdCFpOEPoj9tEsTqKqrNH117YkrA3TA6WmAmWTxXHm5NPSuhWGLfeOo9BIs+
gqXcGdhe6VGk20Wipm7+T1XqqFA8uknW02+P3Qiistn+ExgPTxTtWkhplTnFuJYf
XVkaXVbvwKNqgYakZ8Xsw02qLCVIDp8mAqHM9aYX5dmUCl1biMBTJMW3JMLTIYWj
Crgh9P+Ch5RaRicefAquxgvQZ9fn3bh+AVBSBtZoBa9zvMT5DiggEAhd4winidHO
uZIj/qX5F1E+VNhtzTtZkdPL/Pw8uOdMhoSvmylP4d/qa4c5Rx3JqW3nDibbTV08
NcqeL0rO0xl/wI2mUHQibYeB2lYtJHa8h9LUMCoytJbCjMRN//HnpgwHF1BBYvwr
e52wmqTICAMimJprLl+HROkVX/v4d1tRpyrnSW5pqmi0hSij663LW9jKw9/wk11f
NNAr/fuGmDTveCMr2vj2jUIth3g5kFQrghrpaK1KVozkNZgsgcmWIuZM3us4AUEh
Fmx4IGpmJB48s5KW7Dw4oCiqe5ba8MJKchOvB8rdH9pPiV9rkycmdYKHSaga2Jmt
JnvRGLhUgdw/kwinqIPChD73SuwmlazYvlxkHLh4fcxDehWNVJghDtFHKRkxTXkD
BtQvfZBNY8+EdFue4qcNtkxnvhtX39Rz1cHqIsVPdvo27izBNbyYy4ENpEMunaiP
4C4MkgMisWs4tzefgfpCdNpDkGB9PmxkPViKtE88Ud1qVQL585a4oNoKoAG2q+k7
AO48EhvvPyr/S/VcatbmikqItH/WtPk7YVM0JQrkaHIjUkV55VfggSvuBvtoM3Md
G5mDRtG1mHDWOtDuXhPrpFml9sBd9UQ+V6aSreORd5F7uQ+tgTyNHbrsngi0bcuV
GHBWPtlRgmGV8WhKEc2F7IctErdzWZuOBk0PzyPL2eTu7kxLDjBbCJ87THLOwicH
bNtQt10ItnXJpU1RlO+KrVivWdXojYf6BzWSvJhd4wTV8hTW3L4cr+a6af6HB+tA
xr52m+jY/PoVBoQw+9Q3jmsolW7+cGMiMMWpJdZ/m3PWAIG8sOILAuQjEXq+a6pa
lUC+gnXE8GsVYpgdtc8x8A7pSs04w8lWLiXx/QPZpZlWRiXCpHwCAMRHdrOFzkRL
/f8MGx3gwY2BIfZ4rCIfEYbSlAyRCGXlnV5ordm1tWB8maB0AtQX59bIeV+YPzi6
QZWDfskrN07qqMunoQn9vMVIVi066jjOJ3yTokZAT29o6SgTL72/3+SJsTphMwbg
YvmaRu+zhyCMrIDU2yrlLdfCvcH7Y5oAd64HV5tDCYb4rr0qwpy0WLkz65knXTZ4
lYUai+rPkugiKp1pBcUpptNTiUpf6OoqDWbaRKbTkKGuBnNfwlcPGtReqDuABWYN
PK2GRR4KddKWXzISidD2DYJLanXPk3QgrWsYhduZ7FChijgDXuwD8mWSX3WhCMnO
k0aS1CHCWeaiBRrpbVUqyWLaWVXNSz/w8TYsiZsEq0pim0PkW/2B0jDtZIJwkmoV
JybPuVbq3BcTjLvtKXUJB2XtiUxmtMkioJ3Aj89K/ed4D3DW5mHxl2z+cA9Xm+uH
RfxaMZEEpGAuyO6N+6BXIzAqmG1cgBL2OunIC6Al70xbZ+OMxToiiq1/vnlzFkxQ
YwfRuCLKJVmntZxlHAL8ocWso9E3GnlQjZXBZhcoKjjGX662h5hh9rz1xWo0ARfJ
RjdGtCRiRHDTmEg7/ncpEYR2SIdl/opfj4Iq7HiBdugxDFUw8BXREhe3+7VouRQp
XI2zGdCfxSb2zNCEZDdjhxM6usRwUR+eJO78IH5V9HiHUNe6zjhHF8qn/ZtHOEt6
jesMT0VXukhlUz2/xSRiFE0tcvW4igURztJwFeLR9s1bDrPhir1bdgx9WoNHvJ4W
H28B0F2PhYomwrWWo7j3wJgnqktO5R0lo/N2QGNsnPjX0JAuv/DMnJMN4UWqjhdI
lXpV+U0Y7RdTdZCaJfj8LwdygkTQiTH0XVTvZJp88o0SZqL9+S6BrMPc0LTDr+C2
YM5JsIrSXVITjI0g5NG3Hl3gax8qRX0BR5Ksw0BVim7gFALxQo05YT7grManok5K
Wbi1je1Ut/jhkQsmItNh5s99eXZCkpnwTCE9GUEdhjWRUo97x7kLjGehE0DvYJea
1Mmrdpwcg4JtFNgxHQrzfxifNOV+7w9Na5DMTRS/synoeqjQcrERQfexNOGQXIfZ
49x89j0mgw/pCbMiaMsz9pqT2WR4Rt6WoVyE+zjjUw6b4QyzLATK35Sw1r1gVXwZ
svRADec18um3iotsVtouPBrI7/10piexMFH2cgX9olGNbMHS2bXP/umWYDtDtlDo
5/vfe7CJhypyO4Ylf/93Cp7lV2CYq6eoi+KqwCvvzCtABBP5SBghcF68p2TUGlSX
Hj272L9c707aac4NEZx/e8cTc2tySyA8KU/KXSBlfeJspwSqa/28xyyLBoH1DRFB
3ZUeb2K/8Ns2OV9PXdJsRdh1zC/jv3jrzngyj9ZeSgnZ7xHVHrVW2okhRNaS17pl
5gZZ0bCsvP/b6egJKwLsy57VQAB+OE9eCqsmzMHBVDFPuqAOoydPWirAxndK0hxm
DA3RXtYeI7EaAdiFO8mwIURxgbM5iKCg9DcfA2nkZL2dR4vvx0b1n9iBNA2dn90N
AGdP4YImxF0JlD6qjVcZV+0Dl33pZEifEdoOz4JqaPnMdmRTKLA70/9+3fBBqq05
h/iaaJhz9zFOb/Kc9HGYyqWo0eE83pqWdN42YCGoERkhYPi/O8hkpifqnnbJqqJ4
rVT9ipM7X7/AyQ1+jbROxdrQobSzJHcpO2+W8FZLsQfV6XdXFb6MoCn95fk38PN8
YIDWx+aGKarbA2phmCMwYlcEp5kyob6ArSwN1WQSHGsZl2EDt7AJpWqr3tMuvY5r
3nm1dZBDa5gUn5hznfHY+p/s/uLIxMEKJ8ZuHOYT4QWTClLFjaBKDDAjMhkvAU+/
339Xzs+DqJwzP/+sW5eI5em/XgzGHmCb43QbUF0IfOeqog+WBq2eVTCK0sZJMHRe
Hej/cc2Usjk8sbjcSvgZTCnq6+FL+qF50iJLNg4UO9BPIvbtSxPDNlaijYfJHHuZ
qrmrFRCzHL1pJXQ9RVhtoDohjD0me3jAeRZ3nFjuImRTLxnPyFy42gc2fXl0jSFr
VKqZJNNfUwltuTMvsOTsMLP37Xcs7W9E86b/PHg02Ta1LW2vAx7Yv/IVVkbrQxNw
OZ/ml+92l8D0e/ZiqTFvNdEwzq5eEkpXcLSZAtvS4eGqnBpH4Qs5dcDiTOh2uBcU
fYHvmOEWQsDNkvkwrUk8u3EonxFAKoU02on06h8fGvIW8Lv5RpHSni3GzxBl4aUF
aOU8zw58IP+JTg380R4YQP0dN4bic/R8wSMNY1aaev+8MXwqV8YWx5PaRRjhCiMk
BmS71MV4wb+b6ObGLVOIDObg9gsqJdWycC6xEqSI6d9VwROzSE8Uluy6ASxj3Y/e
EXZBYJlT3Q6eV3X9fvy5rpqgHthJFsbCpm/+tyOIK+X5Q/zxnwdpdDgGqZbhkRmN
vtmaucskRT8CfSpQeRI6JEqinHmmEJiDaFlkX154YOpZ4W4ogvUjhwrS/4btPhIo
W42CI1weA4qMixr+N0LxpW5WBesNmgSzYO3lUhhhWX93T3/a47fC6WXS28qcNb6u
Kx9Eq0n1TRTbYTOm4LOUb3cka61SvRP3Z1nr76SPa3ybOLSPE1N0R0i+cwn9F7Cm
QDzPN1FXbDE3AWBRjr/JHWgEVfeBgWCtp6tY4ihOwrUjKqJRptaG9S32OAcpTzu4
+679F7pniEIBGeuDVJT+VbY/0U50246gSNpd4Ln6SLijTYx8wwixGodA2SGHbprp
IebEGokDozYeG9SxVPJCuNnxaJ69d1iYjZkmvDew5yw7i2qQ1N19V557TkLky7mr
+1nAxyr//JoLAeZB/VcGmGGorB29V5puwrC+Oy4IPF5GEc7tKVphi7xiGe5AOO84
bTGY9Xq2SAMb7hilTJ1M6eA5FUNVbqPUPSFtyuF9EifLR+WeNd7DCcQ8Icly3UO4
kGbVLIDMTJBimF8q/K6uHZNQMkCsCnieYUk1coG+/UVkSbBjyVCvJACTbI7uX8wc
gWS0d4+mBXk5PArj1P2oaBK/jFK9i4D/hZktHqwN+xPzF4ATYn+FvJ1NxbBMijIh
PNYckk7EEXPcF5pPnt6sfu2MiSMVD7nmRw+GsZXdipXbeJZDjPN2gJLrZiG+euEB
5mzTtyFidXzZFP58EDVa3hsiSAneUReaqXgMpTNCf/gOg2LFGrt8uqou2G/wE+q8
FtHunp/TcaU0bLSY1DBpeQuK7E6Okbzt0KBMeDt/bidcm57Wx/XhUeI1y6kkh/Dx
o7SYFiSf8ah1Uip4ShguzT6fFAQXcOy2N/HsH9B8SJSYynjaL5SiVbhQOrLmcD0Z
fyr6Q8KuiOpDNZDZ3RPRH7jiOROxNgO3tN+I13DYi/BDBWlbXuD1ERfHGUdIQ7BW
KYFhOpFyxuO2CcT68aNhgvJlvzZpRJkR8DpKu/z09pvLxVjXDqb3AM8CH6d47zI/
n67DobIJSFxlVoJPa0MITgLGDyz12axkzYMgwuDd7Bf2IZt7D1BQpDewOJXzpNFg
R6MZOi449woosw2KxN6QKjZ7vd8bbhal6/Nm09WhLBgL+aXpHGLms+Sz+YqxnmkI
D8NL7CJwomMixp+XpPClVdaQPTPgxga5ZCTu9XQpesTk0TTibAC9TfFeMLkRpDkU
vSWO4Ki1c2VhopmHm+0j+s0hPltkzbH2sJNn/LRfvmjWD6Ub791f51Hif/rfSHpr
cYjcosJ6jKOnLGjj2H+BpYT5oMuzEstwObVfyPqqnwsXyoh+BX6cSmO9qTlVDo2x
pANCvB3fMudbuwdgbhGQ6kYTDLB5nIE72FAKWjflXe5tfuBIaDO2HB1IpajRn+6T
lntR1TgOdos2h+BPFbAWKv54U7JUvjLHXuHyu6PkCgDkGeFSnMFB7R/mkn0VjIeD
XsZcDte+idvABxm7SDo/ajVyz0hEcnvSYSRrPOWaPJ5Sq1YxNyMa2JgnN+wHr+4j
IzkGkX+k5rNP8hnGNl6ZjVKJUXoXt5FP6gjvk3ot4gPYMAq0iRoAOjsgq6eFo7oZ
j9rNz8dHl+73kWbz8FrhdBH7lMHUUQ8AfkJM4+22qFAarBkV1t+hS8uYDQESBZ1W
ZghD4UNIaU32qTA6hWcT8mNyzYHP5FTkfPQd4sW6tocbctm2rlPJoXPKL3B7sgJr
Wu8R7+03DZmjVIhNmHQqcRB+rvlrfQYiJYoCp9Z6cHzGCLN2wnULLNIuu+0uP3CC
YY17Lz+OFXZ15Ts7skfWcWsSB8jrsawpLlgZMy+feW1YjFePI4JZN+i3nySfrehr
sqer/tkGkTWKBQq7JFcsudwtP9ufIe5QbvTg2Ni+9dOkzC189xRsX+8+ASGl6vZd
d4a4/Ne0NES6lIX0wwrx7e+cVqZRmjXEtrFfcTmt/dOoRXRke3GTOkBdNwUjKVQ5
2p2KiuJ9UuMHdf44Ukqc9MSXkFqPK3RAu07c4IqbX/+mcuGi5Ow4ek65oxiWW8ZN
rSV/InLrr8sRWoAd7fDvHvhUhimkP7573e+k0rRy1vb3GdLcoOL5p8TS2bVOBXls
TDBirJGY4rsOSe/52GavIQPw5+1TsyODdSBnBoElPtubYAiUlPd87gQs/teKlGqh
MNG/KtirFuTzXYWOgV/pO2oGhm/9pkRmNVADOWA3ldcAmKmZ62nMQCu1nJZtEfeM
AXuU/kqZyaBUJtv0he6uu/JgjE+kKeQjI9HSbRNIHXzqDH8cyM2L++gUlzgykcEG
SL0YpNwtdcBn0l/iBaq+LyP08fyXRCgIMQ2iJXJm/f0Bd7MkH5uK09WiYlZOowbW
nboSoAsvzILeimxzsyVu3c4UOWo3g0chlvhTvwgGiB52RRxp2a6U22L6A3ZUEOAM
yueRA4lK5kQy7Cl7LkdwR/5nmhU63C+XMFpUzlc6pj7TAVKlyt5moUkv0pK5r6bc
uQEW3yah5GsQe1cU/uddPE/KTw2MNa8+syNIeiug89PGPBDhUFb/xmCpRVjzve4g
K3AgHfS5r48Jc82vbgfCrJcqEa0ifjZjqTj0sk3Z7+L+c8PoRAge1WdNj/AgSODt
J6hgfD3+JKUeksj5wRVy6flfbKbRxeqlOJKEskwEiA+99GGUokFt+rzka+9lv/gb
+Y+YCt26wgyC6WntV0Sb1AaErPE1WuAsX3FH571G30XrTYd2WMFX2YjxSH4OYecS
PdTd7Cf422xxRfoBrSVFVVlHCQRtwY4Bj1OLQmvSShh9qbo0VAFipsuAQtbNkmUW
LI4jcifE8PJPBIczkIb9Dii+fDMeOVGuZYfkTjSIa+0yy7NNYd8LxQoagilvmT0o
0YcCVDRKQOObCjyKhu6HqVp46SMTgrY6eVsYPvoz+MHR8DFubyYANFaYea32wCMH
C17teZbDDNDXGxOzCN7yc1WtigqZhIURAwSIlZjCFFrXwtCvSdLbnyZ6lvXx6f+t
jtfcMEpnoMCI6dvt6cWJAnmgYX9DKt2C1exgKeR3q8YGhYs4FxtP+FMLBvxfIKVj
9DbRfYl4lFW/nJes97DGGvC2FTpXKGlGH5ef7H5Y3tzKOg36Ey9iLc0gMLqdtEv9
PzeXy1lt95IiLYoEg+1Ihv9omj4GoY1mxM2FZYVyu3BIibaIAmmT4h8ngWSf+w+L
IOgGXjOnCp0WlKEL8D1MPs2gYxoRTZco0u0dex/GKT9iVIssuyYjREvjX1nTjHJs
JQv3x3rGnZN01Cybh/CUDidyWHEYM8YJHtpkQKO1qL3T15U7J66Ma98fst31ozyw
0AXlHEMrV62NDfjQliJ2dJwGXf0i/fJtEvU8OsKjsyhQLl1JyQYglIC93ffLAqbG
2/LlvmozDJ4zHf5urqgK5impVoZjPxUccrI0Os5fLbUvegPIzO3wl7aHP6/m9eYO
adUbmh6E57UdtBFYG7aQv37Id95z/UJ8Z4xL5VKO/F0T8umuanFCgOrJ7Y55O4tl
dqZVpK9XbEVyT5pMaCZvNUsK0KFA7iOa5llzJbg2yfgzeEMHYRR0Bdni0W1NbAX4
QDu5gNYeXQWoQqHlNw/K/2cq5TBWXZHZX++d3WA0WheFdZd0WJv3h8vzuqoyEMWr
S2m7XJqPeCwKw77MMORZQbyS1ZO9a1e8ISwfXmyq8XamvPcvYUfqLWnR5vk3YTsf
snabIV/ym+LBXDOHd8op1m7PG3zddgSjUt7uF9FBwNhHFBJxn5IiIYZLfynGOEiy
fUwUAusTzvpMJkq1Hg/iVjihDnUpJo4n1W7ngtclymfPElfKUrcuIoRxNaw5zngt
GQZEjERAvMn2uNIrKHB7oXlW95dho7tO6/IrTAAC8KPmSO+/pC5aTX4a9T4ntn99
sDPaC1s3hitdRvcxdxMhdP8yzqnQDweCX9dT4cMltgq6jF1KYM15YIpXqrV8Znw1
rAs8pMZ7UlC+nImapt8iX3RChWRCA4Jcj1YfbJyNG/lje+CnuIOeA+CQJHnV2n0m
RkCYsZuqCILzVreLtgcXCoe2BAgc9CnBsG5AISLQJY2kc9/BMNeH9tM6w2Aiat6z
BQb4Og10ORFAZ5dZ+TMGjSpJTauw/m3TZ1wVZkuO2AqhqGv3aQkF4lpg+J3PIf7C
6AUs5RZ5XI7PD9LLpyDs/3oRYghuogA+H8sliZuY2qSTiuWCmbPtNAtdlFPhjl4z
NbyZdKXHvMb9qGspNkM3qyh7fNwxyq2G6rVsrGA0Nd3p4RO/HbCRljbVDMZNHqDP
Wjoe39sxPgaX3YtUcn4H6WHb1YANUlwDtYdJuR09nzJqdT3Gr62sos9U5ri8CZGg
/1beqU18ybZMeAOh6u0m+n0npxKOVt2OcVGHpHprZenuXrHdkb3sUlaQ2QlvyhmB
PA1vqKzzsC7fnRRx7QfndhiXd1xD5rWnJeLl+wn6lQzBf2QTAihX6fG1lYZju/nt
wiijAY8mcZLIBWbGhNce2z3v0V67XpVW5ma7WMNlQ4uHyJm9M8VlTMPig0NEp8nI
I3nwImv9hOgZoTVdorV8w082FARLUoGyMWd++gTbVGXvztOMIAEicGMTN8go7MnZ
cHz5Ke+bHUobFPNEYcViBZUXdr5jsI7tJvW95R5B4ovbLtb+VO96lecFSCCXzKE5
C8uuf4QCnlIQ2yynHnUzsop1b7LnkM96gKmo6REaxzjAeAwVYJ8J98rZwuzbuTwS
73SF59kvPzfc8JPy0/e20bMNWn0jZ09ppGIw9SkkoV5dh0rFe8GZ5+lo7dSvl2Fa
3kIeRknvXtfbdWimDsf0hFb1H/JgTl346xssnBuAKt2BU01+qYcJjBIXy6tiyWLu
U3FB0LGprLKTiQjbu1roLZeNzZKaMRUcV1CcMQnQyFjnbjtjJc0S80Q8yqJmFI1x
NZj+9l/dIcuomPdtkku1SaxQQ47SZafp+qraEvpnPEiJ/R2rw9ZoOXRepYbtYMiH
PzN+auVKwGZXh7dl7PnJJi9b2Tej+RMUhxfDuns54KU52vi3puQhz4N+WS3Njpfe
xOShsuAGlk+AdEcaUraWPknqgXNdsRTRV9QGLhEsOesLvQ0h8NNnzR1WJvgcMZZS
PXB9TRMnZVrU43cqlkRcZql5pz1IlE7wVTKfEG+YcdMDwdMMMxytDAS3Czhvgqvk
0J62nUs8HPVVaijcrMehaFDr92OzmBwJjOwyehByW16eue/uLVeKRQ/aJ8s+2Smr
+bEOQzE0PV9t8Nm9fAQcTkp0xwl87g/GlXSU4SLvm7za/T5PVhCyI8SPDzjYrMd1
FK2JOnfxKaTb6BYBOpdgZiQQmDumWsJ4hJ+XcpDJ0llDUPhu4Gn9LRsFTCIu3+Rp
8LvI8ED7xPpoL/1S0/JEXTOB5A/jIgZetc4kqnRmh1wBTQHHApHLdF7CqG2A9GrA
5FrOZRu7/+q7k+Bhi+ocvVXEFKgvCz7JTYDQ5NLs6iGOdhgEFyWMklIIlMAyaWmV
gVBfc7blwiR/NN6iJw3AqZATr/zQr5hFg3Wn6JRJUyrrPCSahbpEukvzTA6MW+T4
VB2S/oxR1yXHF3qwJXcmaojNuo3odToeAzYhWzwcIgSUzKbuv9WSvwIAspVPq1qd
y1PjAzsT5s1rjaX9kP6W1kCGYhtxGb3fmce67CNLaR4xhBqHLP/1ky2bbgFTcruL
3RvbCFD+M6XpIHU8VqSmhuXqjh2a2/ZIAarBJKA1orpNOVbgQWkZh9yWRwo86V2o
/WCEEkRBbX+s1HjCjep+he2dqIOfRQhRGg2+Zx0yBqwKNQpKo0qt2TatjR2v1nAN
KcUWpy0kxmYB35rZ9kTeGW92+DP/9lD8z8tQmWgesARp17I6n8DnXrTPbdyF7dIy
fvMVUrm7tks+mkz3iETtPiR0nhE2i6U2IyjKPUXjkrP6hDSu0uPXZ6dB5ATVoTTw
QdOEkTtJmAjoquN0azwsYonW0xBx/bkmds5V4V8awfA2bDx7vMOQPsm+81SDpndK
fpXGBdOQVtjJ6D7QSSN7D2jdequBLHPp2WkOAAzTGvmFStpQc3xYryPokHKWSmNu
ao0O/+TqFPP4a2qctOFs7i9eGx3/BJaskCSL5pFjmsslNPnC3FNNZH1yUDUDZrMm
tmNu4QDeOz/kYYhiP/SDgoE7ZTt8grRDgqjAseTfV7YewtO2YD/GnnRs0W94Sv1p
M8my6tmztSACUUj/sFq9EIY1jaNGF3wPEXLsRTnk1jskNnYZ+YBlX6zOY56AqTpH
dfNLfe2MFITshiVDyH452jQ5bDvqZgs3A351Tv5nYV78izrUw7YJPRDUoY5KbXx+
ML+RPVHsi2PDUEvvsQfGWpVAaf31pSlRTzjVKXjrLt7MfSY7Amlzfg9eNjWjEEwg
TQD/qZ6ywbrJcr3g9fFSYo++TtKkXvXgGELKco/ol34k60ovs26amGzF+FOLwgmX
dVzf4j9q3JJWkO1b29TDTLV3XAQRhagVWRgH3fbQhiXFdh23pq8KFxUMM3JeH9Ve
9LCYPmejbJGwWuXd9tXapSnZG0C1iZdhof7j1L705jglCC7gUfBKsrcdWcXoCJjc
9HKRJtGNJjpdvXb9uGKWUZgpaowP3ubRqpQNvjeHQvy9WOn0cN0lBuiVMZhgZLD0
D52AvXNd050YINh3I+BP5RFK+T8i9nZvbrwbzMuOfCI8zXdfPXdc8gBj/iCudGc7
+ISkga/KE6QlMTv76ZQZjjyJaMa5gWeJWXYlfUweFdjR/tRNMo2pGorP84/NQvqm
3GvCrOYMQ8n30J/FITEqrwX8O3kn/6w1GkDyYalpa1/pb8HMCESTI6cZnkbvmGmL
INFQ1PrWqSSGAkZlnQ9xDJ+DOTUlegvy9wc3CtZxHaBHXcKYeb2Y+Q+i8Y1H3Trv
z/Ph1j+x6yZUjezFj1Krs4Ir+Yq9lKLiXuo94NMDSR4JZBlOyN2HL19t1IB33JGC
xuc923j3abeikA5+De5psjuNBqd/KNxpdCFJSflTTRrnAj4L0jxByF1HwiZJtQ8O
W51w6o3DZF2W2ujyL4eyCAl23t8uTK4w9aUrD4jkfIGv0g7AhuL7e+4LV72nsswe
9XfzsGWw1R6GMR9SmmkNyswJjtInZJabDGPHp7ZhIxBKgm2Z+4bN4oiCnBq3YC4q
gpIJSgU8PYe+cT6ZDdsK2f7ouqbZYYjJ3mtNJAiqL7y8gYP13j/acVv8G2lAROMQ
6naatShNx2F2UGI5p44M06HzXI3mZ4u1ZMOe+VkD+xcx08jBEMzg+isXx/Zy+f+B
g+gGV4iOTfR3AYhsi5NXW89UpcQ1LNwXe6kJrZ6gDWj0ejKHoVn3W9F6ab+9PD92
YWuI7R+0R3PGzaCTQSQRMAjRGBptemxG7nMrj+GU0bHO0gYuGySzA8vhYk6fXLwI
yQmM2U755pohcxVD3jnyqD9+UNR14Ku6N6NduC90Ud+tabm/KbU/z+JXKei8SHVq
MPsoLlko8jiXbmmgg0JtOe7+pyTpEltzYfOHcsP7tis+Vq84OuTB1qzW60dtlNNE
+luhnM05X77W2p3ntxFLtMffOuuMQxCwBQfIufYzSneRZ7V0VoSa5MNRI5CJgiyQ
V/HGIVCmkGMtWSo/NuBF5Y1YPYGHX4ByexA1GD2Dns6PEV6nIJOus0H7PEBwmirc
McOmR3Ht9ROmUFA0nwlipry9P/vqm1AP+3H3T/vZsEA1FjctAuk95a0K5WVrVtHP
AzjeVWFjHYeOR/EwC2sKBDPrXLd6g5zUNL4+2tk9LzMfNvAdwLBOAfOTnpW/S/Tm
NSL7WiGID6P0oYytc+/XuoXTNYixFDEHpbV50F8p5Q5l8NGkV9NhZwqKkqolmKsF
+9A9tqTea8HJ4xX27jgtIaG6wF3XlzNpoW6DKcFPbRxv3bdV+NkAZ/HATsnM+5Jd
I3Qcbi4e0z/cft8bKyCGYXSswRfrsS78VHUYkeILbBK7i8PQqy/mZZ3d3POK3P9K
PnykE0UnmxCXGGoDdcTwIFPuZSwiNxnRGO+nXXl5r0+NNmT2QwRHRiBNJnYP5hGw
HKvIDeG9YNfSWHyGHuc12RHTCFIxoRtYmnPhBumyvNm5RKLyZzsx+oGeG58CmkKD
q0TrdiiBJ/6LTWtTy5BR+XbUQ2J6jUOok7SoDaxcgVnI/DlueEOQo/0vGBF0tor0
ryE8tGzdzBDbLDUUJHPTY5dKSGorzX/VPCDWWJ/RLFlLzRUKkZa5sn9MHJaoPbVA
KOJe7LPrC5UOFfu0obFtwpfbPyppgDBenFyS1+gjHoenSDV8YceOgZ+YJNcnq/on
Hu33ziJL5gj7U1ibb+7LmVSdDHcrXs9zVC5EfoXsXGGfCXDmJHhgyZKlfcEvqODU
ffxURJ9u/GGEsH/Xf4SoQJQHqprVRKJRHQIrF8FaHmiqh9j4OjeFNDOuJU2KG0Vy
L6MV2JIttdGF+ibMjfWc128Kn0gpgMKNaSbGsvJ9pCoQwqYjrFBs957rOuQILB0E
ZEQvro5EIlUjEqVgLBL++Zz0+TlM+GmsV+Ew5K37zPem2OcaIykW5aLIbke4gIRb
8pddB2py7kSxmgHJlvwhxmXqG2Ct30lsCa4yF1WRMq3se8VNGIezOKia6ro3LNWT
6bx1gKO8n7yaoKmSPtgAldTpCBOLO1/yLL3LZaGBhKjGAb5fHb4rF82Rl+Ni+80r
x5OAsLniLAC4ptCqW5FvKHyhqbKG2DWn9G+9t1dmzs8iST7yzEoC3NzfsmikBtA1
wM1dqXVsi4hM8RSgQ97E8OA9jkP+3tCzLQ1Um0Z88RrJL1cIloy/Mw815evYkNDe
uopNDfojdmVI47yDX70Lvd4cFf8PGkVmNex0qp/87OCNay3y3L5omb6qa1tmClmH
kGBsy3VSno8g/08oZXfeeWOzdB3xawX2Psna3WUQKmRtWZK57l7MQb7CxRsxnCik
4kROQNqTu/DBA6HimjyHZz40oE92B9782JFmK4eH8DdeHgDpiAvf9zA1o2xSNQVb
nAciEWR2n73xlOYX9GP977LAzOA5SB2hVLj2Pus1euHNwtc8kZjNvKWavqCp89wg
Iccxmcu06pjDgdD9Kzf1Q1dkl0YnggxScurZZ6WxEPcoAsd4OgUuEju1HsVeoF+0
QS1z7/B8pXVfkpVjSJxSCqgc69iQN+fnc5+nqfM7A3ScsxTVWlq5swQPIqMEMidB
2vE2x6t5JTXau2TB5QaXXSTv/reM9xRP5gMTl5Dzikwz63RQUkkSxlKo1AtBZDFm
BrFeh2id8yTuvxzQKPecyGnz56bQtEA8SyYOh+gwUhyWROiWx4Dbys2dADe+Vr5X
X2V5O5UCdcjy4zGITwEeuQo9L6NCqXq+YrP8zBm37qBKLVI98So8zRDBxr0Nu55g
doo4O3TYm40VUsQGUMXjlAng1v38uIwiifYxr7mQEwmqbFfa+WGogwQkiHasEeuz
DzydI4vpXvYa2afWTm5bsvqgY9UlaPDRo0TT/QOEkd3G36JJauRVJxU2ab47HaQH
5lQ61nW18uWPXdg5mgFDjvO6FmSjQ9u+Cx/FX2wVwmsG8wruP15FvfgEAO1fuovz
3z/Ek9owdJKy7nUdkWHB2+6/uowUtr7dlvr4LGlDbx4P+7l9n3GHwDNiTeODnp2E
y7LQwYEGDp/3hV25jcctRe/TD9OCCI9Bk9zzdZFVcancxlEWvGc6Zb6SfXG72U/M
vAckxYkrpukJl4BSDwTNegYpuhUsbNB10Hvk8bFist4DPZscTHp/z0BGVKojOeGa
ya8GdqQB3yt6kKNcWfm7E2ktpBOnUJjyZH6uF12PxA7AoGw3MCl8OGr7huU2eNow
y7J5xg10lNJ2d9KxGsbXD5sZ8tNYJ8cu3sGffceCmMYGt+/QD5EkDSOs3L42Dmx/
G1QvYtg1BzVmcv4K7Jka4Ouxz56UVjgkhNycRG4ZMcjBQf0Aq1soBccsDBsVDBq/
o0pGvlzwnV5TSI1LLHA3q4h5bfcCCQ2M+Rzecfnhb2yLcJqDKcZIXG8XWVipqX8I
Lm9+sgMtT/+sFsP7yxU23gnKKwnkH4scBgxIlSu8Df49SfKOWITWWC0bkAOF1vYB
ko67WG8WpegtTH4qGfxX5lTrAvZyQ89KdWcC2J8TUNZy3mmGNwQSGQw8P/IvI3CQ
G2SEAJwQ/llV0VfDfujKa8d+fHsN5ZYOwE0YHek8mHV2LGpMVXnQ2XFXj+fIGsKs
qXKQx12xAr9LTpXW/b5cbUUUTZTIPc7OZtOz02BbY52Xh9/L5DdXHInxOdN7q8yb
HpiMojNn4pEJSHbJ1tXGovSiCrOTxQEQJBH79MWnGC039rtRZiSyDMs5XxyEF5+m
4fmr1val2+Z/XEsBQCxPdosFLVtmwAwWmL7TWvEypMI5w+WuNZTXCJ/GGpi+66fn
ud6drxU/kTTWY2BFtpXbjxqMqquHEJsmRuon4eAzBTe/xIS98qh8NuIkzsMWVjMh
qFU7Jm+Lxf917F2FpdIRWnqBwfymNEhZzw4iGvmla8442GQGe9QYm490IIFRE0QB
AOMeO5r0LUhkPlwDDnm3HqEIFJqUXZ5/mhjSdC6yTDo0aRG2PtMng/eT0og7lzRL
hH+XrdOLtcb2Rti/pD689FwYFBKcSuQhYPD6BhnbaEc/NXO+dTu3q3Cx9zXIo0w9
9IhWWgNoO8gSRR6Gtw2ZeVlTQKlEbPKwnMLj+3Ygf8cEps8cgdkbcebIASYZzUa2
TCabZOK7yUftb+uk3JICmCuK9L4H758U8AliRloZrU/9j4HCJTKKq8tLdpD/hTjd
N6Y2uT6EQSGqKJej4XShOPrJpI5AUE9sH/KlDhyJlGkycvyYPTunfPs7Gt1ueMBV
id7onmHUT2cGUY5wB7z33FC3FoZPkfN7VJSnMcb4I92t3PoyMy5fCvM5qaV77ODM
5SjsD2MFlGoTQ3rXoMBZ0ckitVQbo99KDQtCXjWNfsJlLz2rhYdABVmUFRlJTQIx
o8ddP2LakP23JhOSu8WaAPtP8AoIAdrTarPYNJdtaoQfQ3crjXDPvdx4grXyufwj
Yh36ennvqsOYcretScLcJINgxgcMnPx4/QIirlk46uJYOEYBUnxrK/+TqSLeYsMc
aX2yt7ue0HatY8pAjw5PcjniNyyLtumtHA0ygGkyiUif8EeaIm0smm1STs3krmzO
XOReE0RgN7mBHrCurJ7Jd1sq5/6drMQcpvFcARcRlRC8wFQWL9E1DxmEVnNb5vGI
CAAnZJ2FAefQ7ZaoBT1gxQK5itwnO/E6TgruB79LNRX/am2IG+ZoZ1eLhvTkxd84
76q8rxucwzlQ/i5sC+wsTZS9mr0nqs5kaxlsWX6sMcxhJJyPDU7Cm1WxbATDscL1
4ZrxpRrBTVK3jNlWI0Q5Ik+UJP9ihm4yUCBxtd+flIgsxh0Wc/Sdn4a/Mi/Y/Xb3
ql4WMU5LrVULlhTLZsIFPchxfKvTh8eXvW9QBK8L3E210yD5Ynz4eEc2/yOv+Yzc
W0NOLlLg87i7tUdfqkb5TWkdmMcwUOTMyeG35mWv/c1fjl2VRrEWkeIptRS4Or7d
dr2VMlL3CY8fWDVsYW/eafZm5qSU1CJmj68HDzpFEU5B49D6zZ+80f24OkVCebXM
rLAhcyAyjk4xQ2wRGlF/E7BAmLfMbw+41HaOitGErGlWmAT1zTWXfdETpmx+YyXa
0swMCb4KES/aXxDKqdZnSAugmIP7Uv7+1w2M16yj6kA3IW1w0Kh7XIXoHhdWoxEm
3FM8z5Ai1T+lmfZXsOj++08JhgY6h+C6myyrl7XeWswhZaR0aGAkEkZDeucYJr2i
WyZ7/inzdlB/NNRMsmjAwEZueU9Dk2U825QoDDD8CRkeOKLHAg4LiWub8WoDW9ar
7aCWlpbfuznNpXHOTsDYOTyKPTo8PCo+rmkel9lzdGtY3KDdt8uBKKLV5zBJ8grX
SnE7l+scVLJH4BADlj0rNCgdPF9kEUHNyDTOy5YTSRGsoCAwkJee68b/Wd9cF7ua
q5YUX4uc3SYY3z1W5eHxID2CTVmppBYiF+3A0AleIkZadgZ7sBIaiiX+Wh5xkTPm
1GbyoU7m/CfpVRjEny8irgCWnTadLo9iA1W7Rmsx9rdlDo+SHsZeHTjqhlNdgAQF
mYQTEQDuRxCt2yXiuwZiOS9gTnP+Dwf0OEu9Y++zqdLFQK3yyKSo4/tNSXTvcRX/
VduYENZQlxy58hKE9cd30VvK8tw2VERCfMOuBEQU8a99ZY6x0tmp/GUWGl6PKSKF
jjonpoczYvCzx1YmjnFYvtUgsempbqObg+ykFcb0iLPRd0HwL11RqUpio5jLuEUn
YkW2kKeFu9yYRgE4NT8ddttUc+PwEUqYp21RYzh45HXZNFhsqoNL4azDzQ3L78RT
N5zf+4X7Tw+uVqLUbymHU1Ys/BRgLEQb/lbtbQqml1hhYQOWOZzWXvjoVP/PHco5
YlG14/HZVjmJCfWsutTUqxpy/6KM2m+4Kdtnr+sH7Xn9JrIEKEPRoaliwUq46VgZ
UxAR/rtPaEgLEMCKhqLjoPcYzi51iXIgObCeTekoLFKnQAPH7D/afdTyn3T02oDe
5hxanaeAT/rG0QIyuOlLBh5jmEiHBke1KjTGckTwkT8yVdRty/BMlpqwU6+8kb4p
FiTPejidoIY6iJ04TGPVElhcDW4BJYDtjM3c1x9Bw061YcpqFU4XqpXGNd12HXjC
NHsjd//OyiFeolW1g0TeJeF9z+b3tXvkH1658DbqQwzQhmKwkSdq0KddTMCqyIRc
oZp+1ROWkzziEqnWbi3WCswhsZLyp1AGSN4Yx3qECJ+1864mMC3t85x4D11PPZOZ
5z0O+kXmCvTMKpks4A9tyS3vuzsfkB5OPMDqbgB4CebHjWSWkXjgNJY0K6YIb+pN
SyvIPI55shTqiUXQ0IDxpFM/LVJ+0NENWpvs9NkmQIHX0ZtkgsjeQdfPlUNawXUo
Os4CgujNNzo4BsdBEmUvrwt4vR9I9wDhuWEOgNh0cZhNw1XZH6kQSs3n2Hx5HQ+J
vGxztsfYjOq6CXYLqd1FGwVH3aAyYiMR/4mim5Km/4921GqeQGd8lqpZRw90Gfvl
n8zOn9vNpM9BtpgLe520MG/hi8JZ91hbF+lUs2MibHO58b7z0Ax5G1FfiQFgtk6K
XX3VeSajP8O21amcybtKi8RLKOjCZsWJMnD1mpbDh7xACo8G2WFOVffnt74uwgW8
sfTiXImkNO8s0T+VCHDa/lsx4bK6FIhY7S5y1RxOSLAGmikdGd8oHb/su2i1b0Ao
vprchK/pMm++YWh21eemDSrtHnPlz0YuWTcX4ijhzT34EMEz1WqHrIbxJoFQTKwZ
9wU1gHYh9r5KHsiNhDxrfSb6LzgcVpUGmgH9aH7X1DQpbZFcJN1+gBFt2dPDAryI
8VooY2XDD8InKQjV+ZQPLOSKAVi6CnROwUq5Cohd2A+S5sv84CIVoORh6TJJx5je
zXl6b2SUkMNP4Lr1/igbmm1WFQWDSzkTOozRJA+Ea13IkaiTjkDqK3ZR+nmzZ3Od
d0wlb9D2BwqjHaLGJWEr2p0QrlB9bYtpaUZfyjOnDeIMMlrxpxJGKDlSlJoDyOPg
+3Rf1GF+lUjKRsrSi+VtqFEWiOYTT+xr5Zerwn393BRrzcADpSM8W8njAIVEDBbw
VOe5X2qs7qLwpwBVC6GmFvqocymiM6Kcm8AkpFsWsL2Fj7Tf0xlEH6VHThJh72Vj
9BVQV2RBTq2YQpyROGTdDHdq/2urjqy0fUT/IXfe3g1J4u1Jk5Cc7XrQ2Rf7A7sR
jH53lyNUyAq7eQ02yBN8QzlhiLIIrx6Sf45beudSLhvOodwGw0PcLkrdLBiaOs+T
z2x+wgHcYbnVigiq9Qhh1B1vMGUSDBOVGbFB2BZI0goLI15CaF9DVexWrO7r3jrK
7XpTwy6OiEEBIuH/BcH8LCgH5N8M6om7B7+JnlGZShMIgSV62sy06Q8Gg9hDrm4R
hg9fyO6/FVMA2ypafsN7v4POkehUeoWQjcIx4eqqfvz/Acw527ZV6tpo2ntzQmb6
62xgS+t/M9Xou7V9GLhw7sQZFEMvQDmfO2iM7W++2HKgvZJ1WYy9yZQWewcisiBx
29ziP5QySXcfE9aRlaPx4GMYAx7RHaOAKxJdRYxumrY5vmFc4nLaTwsHr/q18D5w
0n+sxHT0KMrQnQozRjoS6HcatOdw65Rj+SNAtMZhW2SFNuytv4n7h0BsBHVFmhDI
Dg2XtCvKzY4RBKGz5OsWQq4gN8uEszfgDESB7iNiGx9gCCGYYafbKvLN6FZcPzuy
myE6khiIdEbONjBFbsuHp46Hm5GAk/XpYBIJVqQIUQm4ymvqPZag/PHQAgnkhZUn
xZlMUThf78BzwHnFCJTm/sz+l520olvAyUoKsnUhebs8sw+dsDIwWGx92LYWgHoq
DumMD5uoIA+ICPvNhgd/qLWJWX5uY2MoNy1G2wDE5Ar8g4yg5LGxHcEID1Og/leC
fex7j6zFpdzBNTqTr1/kQnxcQEyXFOI3q+gppKjuur+NhmFN6cqSd23UNUx603Np
NMl46pqM0f62o8Y6oAXIJd3jCun1U8MVcm+mjaM6/YMDOvWRhRWrRctiFkhSyY7N
tqW/VANpWlMVoCXWs1KdRWjtPszgzhvxXutUE5ZwITQkt8EI7N97vLBp9hvsHAMb
/FCEf8TalQIYzqA8S/XCvcKhlmy+p1nG4jFUVmabsDVIiU/Nl2PWOgU4oOYVpURC
7ApkBzCBCbdnvzxH7IpX26/FJ6shoo91igxa95IclCWZ5AJLMlNPB1bSeLsdGx5Y
luKJMUEEOEcHyLuvvKi0frOD3/jTa8cjeicVWuVdl0eEdOV97E/1hV0zzin28+1V
MxFzpgEiAMecROgRLqNmmRwycJRdW+1n/Ptm4fR3U5r4JI3kyePvPsanKyr2t+q5
iplOGlP+AgALfLwr5+CYj0e9COO5TupJIoPMz38CubsO0mJrvtSfjXMKC7hq75+k
4U7+t2aEL5PAKoWGMeviEKdg5cmIaT0Lv2fC6b0vbJ6RXFyE6CynaJukeJg2nYRI
/v8V2moiPANKFONcEO1NlgpJVlFuBK0wxD2mnEFJtbYhA03M5sYjWTUab9mcvcWf
Fd5eOTdky4zYyw9EvRk5UlTVmzeQqkmSIm3zE2L1N1Km0bI3Ily7qgw9f1ASbXJ5
9NwbZuQvNukZaHIwVy+wFPvM1exF8GWbAuugJk8TGQvu+fx6VpiPQumIGzWYW9gc
ziIKSveuwF7yBbE7DvobGUYX05vvRe6QL8xdgmEhqAWJWfRpDOF3egKxc8KpMsrq
cCivXzYtPCKkU76dPcQiH2mVZKr6ABvMFvmipKl/SXORGTklQGOUKk48kapYcUCR
HpSqMV9Lyufh+SFMeuK+qc+4YFPnrOhz/iNrKV9njcLCFnvmeTgJzyUpzdkaU2Nj
uyInbPKBwVBz4x+dSE8+L0DAENsH3xYVuUGn+ilG6mrIpQWJcanJZJ68qepAt6dP
HOvOLI9QLu2/0lCsCzDCPa5fMiwWs9uDk355b/KGuZcIY844URogSBPjtWhdVCHV
iI8N6koy+mXd8vjFZMm52XVq8C/Y1fOootywofoCDquDuVFQqwzt5me17p2Jq6bG
BWND6BX4nAbSn7z1Eth3JjRi1ukOrZ0nmD5FJP8+xNVjHHHNL3np+oKf34w9+APy
+ylW7bIFungVHXdx8Td4YwVKLv+bNBaE8zADiFC4dvxhCi3/Z5o5aeMFhISYfljE
cOhpOxc8AqzkaKzbkx6/7rGIrHKqRqvqsPJyc/IO4C9gdY19n689d/RO5SRZOAvr
JA2J2034JW/wmFiQ2rFcOahA4xsKWlz7bOKAyuQTbmEaiLw6lfyACTIiS+3M0tb2
6FKcxliUoY5GKqCoZFIo52R3nGdEH3gQdbqbN97v4WVuNvq96jgTDVJZBgXvDQ3i
PCEYsrMzuruKJms5q0QEya3Ddjl9fDF9IdT8n1BmYjSRwwkmFXMfq/RjntrNN08Q
kqQjf/RXcREeouYs5z9qDU7cL19kwU59pUe4V9NA9T0KOTbQeQYg4ouWg8nu88jp
kxrNKDs4GuuhJK22IxIneOybCXAwHojtNLDLEkbzJQl+TN2UXSKeG3qTe5otNY6L
j8qAYqMuUiWxYcRuRUTnStPIMLal+o7/NSFXw7vP4ZBTRfxsLv0dXm5qL7rVwtPK
YGr0Uk+kSIIHjbdgKUuAL71DmpEjuMKRztkUan6Ny95cB+E4I2Exnhu9BVMwlbSZ
tNLKOenoVLi6N+GcY5pbXJQaPk82rcfrol25HLuQlaamJuSTSR1wT1WO0aCx1ipk
oKEeVYPb2HBBJD6pyM+1Ah9chqlAZfgOfL66Wz1KAN46S/6w6Rv8yeiA9mGjs4nS
wY1FUt5U3bGe43sWnwMUq0egd0s1gCHs1qCnoQwEPto61zE2dA5+9HYlUfzngIGU
CT5GD2Ui4cdQEkq7eBHAeyC3iEBclaOUkF3rFjdzUo5STMbONaKs7fPM5mOODgQV
jIJ396ujN0wfyRKexqF7HwBCXdOYTG2i8ahaElyQAELuEFWgS06EQ3z7fiC0E1AP
vBouuEGAxECs5rYq6ZuTk2ETCHkN0WnW5m7IbTsKR9xt0HzaHx7DY09h9VyvQZrx
AKvxlcc6uQ3q5erikxtVZG5/fObkLGTKeQnsehwt/WydTBld02PbUpPbEKKYCkPm
10+ZrNPHwA1XW0hRJxxqpp8Isp6jmPxaptFAFRa9iXUqV4BY6moPvKGjmnDPT3op
Msfx8oIizHhLMG8d6H3tKm/bE26NabBIzlWVLFQ049U5KTEcc/XBS/CwbAypCkuL
XBBG+ZAhl8ImTh19Bv+qDbSDdlsWUygLZ+F4MfpdSr1jdnY3bFYy5sLYhzfua62g
E/R1i3sL+mosDmWbiyEtPlbl/YwzQkc5dwaN0Vsc7xNHHZyAuT1jfTY+houihmWZ
hw1wUDg/EI23hEAdK5fN85fUBlgRluG4Gcfc2wvnSRCxhp5OS2BwbLjJsO4OozTo
fGN7zPCsjslISAleH0GgrKhFviNW8SqRKtDte4TuqVspc5naI/CQ5rLJ9ZuhBQkl
zFofaKEoOoG7q0UuyCpOFic2eT+Nvg7r55jE5YhGhz0GJtoGP7CXsqlS6+uB7Fqp
g9oyKf+NmMRq2kwTRLXcc3Tx3UyfcpQC28LIXlscHEzD6vJ8ULOaGkLWUVWokv1h
NDQ1rAHZD/L8iJ4UH4kICuXte2LQBwMr3/YFWaYu547CR0L3SdkwpZQ3eoW7kIdT
hKl75KvTHl7PP5VqxPGMiCnshoiG8+V3C7sl2yfMznjrmp5nO5m0OSFGttCmG0Ju
DsKEjWY4UxZbNIw4QvHBpHNs8qACRBEuToub6QqBow/Xtsa6a+XFK/l5gQ+tPjPp
MbBqVDG6fkT9xC6OO7ShoDIDG6EcQMZ7LPRVBwRE8+ii4YQOMONhkIhsk/8W8QyO
eaY7vkMtdF1MQdTxDp35+xa8BIbDhotMnSspSJ/d1Z4tMh/l8eWHBfwDyN1J8yJ7
r6BsM8Z7ldxldtgKxNZOQaI+J/FXTPtOEqAgC1dSY2MeXcbl4wxV9Zr8dff6jXMo
tExuB7aC7U01LZMxlp+7m3bg4krMoORLHS4Q5iCZ6Z2PpkREZw3p+VTetuemxBNG
92I6mTQr294oT7xzHD6Do5WYyRp7vGSNjW+eqj7TvP24ghjcdmjgbkVu4SPcIdCG
jdDJEHqve4j4SKxWxx/eiXLdpqZGoMnvEXLHHl7OVLVyoyffKdj4LDF24j6vv7tz
OyoxQeRwPIcUNq6x/qPr6iIuNj4qbSq2YxMcVn4hF04DxpFHB+Ey5jdm27tEbk//
nPxIrBJUs21RaX/dohAk71RX3Q7GBQhaaSVtL8dkS64QXQXipKRXvCYhzNAxSKEm
ZPAesRAVECNFqeXCI6pOe2NSwoIkzHWn43KiiGhqJlhUB+SbuAgr7jbTV+ErDh1L
WQGhcXugqRnPFw/qDE81+ZXSJtri0rrPK5eaLsMvDerjetGffTP+wYsSACu+KRgO
TnRZ2MuJmeTB4pNIBPcpZQ9ow+sB3ikmFOh+Rr55zT+Ld+ULIBj5Yr/8a5lHvRhr
v336yAQ6eEhsdI7H2pOLHUrOtg+f8131xO+dStSm8VNLAGJosEa1Qj0GvqnV5JGD
B48nPKmvsRFSeE1UaMVyhWgE/EJXO9n3kkg/J9gDGS8PV5YgJfZLr2n780VzSWaD
3p3/eBuARWPIxuH83OopO97/k7k/SUpW+j8/l3UuTfg89cyHkslKMpBDPwHAgvkA
2gnp6BPLP+OdO1rI4OoUyCTu2lSaj0wM3Kr7fyMiTVyu9U0TvdTJZ1MOEpgyETld
VrrA24H+ekkXj1fK+eVSBi88d9OnBAxBp1dQ58OAht2IocF41xyxqOTBlqaOQrsc
Qpn0pD+FPGmFb4kVmocTzt13ZXW80vARCFZawpnVW0AtfjWl90mSNH5HhhAj8NC1
L6L2uFvS1/BXHMOviio3ddjQjqihTQv6rCPaLLZBhXVdyLP1M+XpeNddcwReEWtZ
nc6ALkf/Z1L9xdwZZY4EmE6YVssqZC8tn/MwsOt3LDqGQHqU7RYLpbz+oF5bNHKQ
5wFXn5Q32K74MwlWuEVAXEf8s3rA9aHJQv3+Iva6dUWAxkrrO0sL45tC2+0LVWVw
9q0dai4IzogQCv7hhjhcba3H8FmLM78CH6KIMLfq9hG8ISdOhAak9cZ8J8Z2+lL7
yP5BjjcD/PU9BJoN65ZzUvDIUquMs2rEKcCOZac/9wHgHl7AC0/rsJdKEt32/xY4
2awvgGgo3OxZ88izwHzOqdjB0owAOWSVD6enO9SC5UXc+yw7J10IiuQ06XmX0k5Y
nBeq5jQAq4teZSwARSnHsA3HGQ4B8Uuo0l6FmvIqnULjl6WTlxU+PjcOm4oN4lna
DDsar30JNAnZHJsrblw/oHlxgbIX1NTL1m6DMtgs8s7ozlrBY3VeS+/2pojz1fOE
q9DWVUtY2KN8XA5wNgkf8RFWvLvBZJ5GnsqFiMt7mw00LboxeVs1HgvUxpy+v8dp
Se1FVK32HH8g61EUwDrs61dYFmmS5yNNW6IAmN8tDqev7fQN5VkfNqguCHmJXIWH
VAPdqa35UtvzB28eG5+R3nT41utWHZk3+hFR8i2mwDgfytZ3RtNsoNTmqT/aozgH
Vg9kWm4E0mKeJAaX1ApHr2CU0fcNVGxVxSgORh6Jxb6DLEx6fRwZ4y6Cu48gLU3c
DUj7x9ZTLFP0qLEVlnzpr024pjrcBMPh2S9pMYxvi1Mw4epSjHC6jh5CXN8qymfv
w7ObzdGmvulDgGvGT+LXwj4EXnKhIb9nEkRrFv7m46FsMI9uSjPBJfIdTK2uLFd0
udF7vpg0LZfD2DxDfVPrmNqQzYL+dQO9HMTtzjrcVB0IbM4nDY8TUK3z1gvq+7uC
QIaWHSEAtgFs/q0oOdSK8Uvsh6jDylpLIgP21eJ1l47N7cPLBgkRQvzL8uVELwsH
vJK9ickY1zMkJ8Tlr7DhEKS1R9dagMSjfBHjMpTyogMrOSl57cDuKOHiZ21CLbXC
6dW9WtDLh8vHmgQPAVEhYZn1r1BFJxiVxhbEZj9zLMxeX77xlaTmD7a8nAHLCvUG
bCLCLv7N7dChekoAXU5/7wSXZqsUmMwvzb09aSzmVz1pg5xMpazEsC2yBDTx6Dfh
iZy0/SvgDcKvhRGaHrtZ7jJMRw02TYUwEgj7zaW+xnPvAKA/oHka7AdD3woSslzx
XT97OM9xW+Wc5zFmv5Fql9w+fL0HZcyHEYRER/ip8we2+nn9/55d4jcMLwXtjgSz
XeOp/9eUY7hQMl+x/H6hjXpSE7YZLbGd4rToNm1obHAxnoqpCzH/m6xIfHHWom44
7CHo7Sv5TL0ZFr7CmziPgC5nr8YBJbbv58dzy0Nj7QFVTYNEfvukNghreJ01UpuX
mxo5OoS3dRt11pZhCfD3kjqGizXTJwVlIfvZoCbtHuHIlqdd8ALzcLup85VdiSd0
6aBHcWulwpgX3+EZalZhDh5JEgCufxnQU/HEj8aw0sZ/e/a242aBqLOBy4f9AxR6
Pheh9WjttgZRHHwIh3ceQi/jo/KDbLCwthfm4//MZxuRglre072E17WUv2vRCzox
Ez0SX2yommj6AkJOwGR0nStc23eBBPDYuogI0D/XQgdwaORIQKZ2kCaGKa2xNqH8
XeV2YtJDPxudqVUpf9YDOnOvwlF2yra2n8RUokechi7D1Ou9hclAkS7NPu6cNXtE
DIQoyIU2x2xhQj4atRI9+MVtHTfPqyKUBbInFAI5gPekOTZGLvV2hEjN2agddh9o
Jw+chKlofTYro1zczoP6FBOQx9d4wa76Gx3uNYA68R8Nni4xogsRGtU0Lo//RzCY
jsJKZMMBuVDrR+loUh7h9BHUcmm2fj374eX2GY0qz4AUTwUkom1gibkijuxTf4qh
z9o/6dC26WKoPlf+T4qkDFlnhtYyVNEjdFCpTdtj/PHk39LrbtfQBo71PTPb37gN
A8zna0BndQp3Pk07DYMy9fA46YWCvgEtu50GeKsOJATN0PNPNTe6J9N1HdHlkQCM
kv4DPS9ggScjb7OpNSJpZwhz1QyfsOK5ThBKet2IWvnl54DwbbDUpSjicEsMEWn4
QLe/eAdQT/8V7a2fRt2ZNPk7HQxEDQJ5owmgPDEY4CPphTxb85l1MiuWlQFYzYu+
XMsanQOCvDwGKxVzc+VcufNH8Sa2biOQ4D/r6X8hX9WJ7RkiuDE2sh8PxWkSW6We
pAn1cibd8gohqdtXe8R/eRo2qBZCVRkJmwlZ3Ciww4fNdn9CPt09T5kfxVU+5sBm
IuWl9NHQpWFoDakqx5kdndrrD6jFBn0YZ+f8RUx1t9ZTNGYd50767uBgWUA9Hz6b
mQmPJunsCg1dzODa7V9Eurl2ZmL7weolhrXN7aT5+RC/5d+3/YLhuDrQto0mjuve
pxWvh0YQ9a7gqZRzkYvaSBMBlrFfI/jCJcV4XjmK/PvIGipurMnnDgtScgJfr4L0
wIdcP/lDl07dokSTEdiMmdkoxQYdEX3N9qBZysyZbK/L9l+bLBdLj7aIp24G0PB1
Zvw8Oa4NFMml+kVFyzJeO1DAxWPMpWwMBg9PsFOW0z7xu68I3Zc1ua+/3DuFDVyK
1cH+Z5z2t75Y8HuZhA7nKm0GiOC45Y4qpdo1khAk8ulvHEPpsX+u+AOo80p7XC8f
VSOhr+x29/CUu1lpJpGaAjCbq8gG93CyP4LnMF9uug9PWW+Xu5NMP7ZXwMfyXxc2
Ynxan9YmADxy39Le7t1r/WAHQpxDWKWvt8U7iSRuBCYYS6n5mlGVYl0rfznCjLfF
eXDl5wC8ytE9ZWy2B1N1mNjcIBwa8HExUSQfR54N+hmuHYbi/DUCrquvoJ6OVdpk
xnEGn/QALVW6+9Mzlu4i63yw7LyUZTMvdBCVCA3G9RrpVxg2BkYNVfzlDISAyVTm
tB9flEwiYK9lUCYISxmkBHa4pjxqskkLTJ7dZy3QJUTC261rrBr1s6PmjTL/+QXG
kdPRyTbvLJZrscWyFhExmtWJSbnu/5gm5Axo3il5MeraeoENAgsfp/TPTDvtAMf1
Tv2ZuRcssZIvxvc3x4vL7k9yjEXsYGM+WlPehOGDjYzcC+e2hL76HlvvciYr474t
R8aoO4gbAPz1gggI2BKNx7j3HZNy1t1+JCGLAT6qdOA2pNceLYi8joRBmtYYBvb+
7z4m0oBz5toEo6nP7tZhYktAkf9KCUeKrF+NVY1llA/nlBkTs5pBoGLGpcujL7FC
G2UHNspgpiIBdn3F0JadO2U9mdnDwjBQoI1Zo3yiSyOU+noU4IM7K+AMFePEbZOw
8NgHXlXyGHlYDWh+CoTB/I3hvvStoAHKSwVF8R2y7jbEhWZ5j6O5DYGhLdrl1Jdv
P0iptx2JmaaH1LETQEczGG8+1ZGDw/ZpqOJYS0+LTPwWw/dzasefdHFCP75JrBiQ
rq0yc/B+rc+DRq05DZau4r2B3RQ+PKWDOyaw2P8Q4OYXsDXbYZAg+ls3jA/Rawrz
6WQ6F/YkY7h8wsIu7h/nVNLzIbdsIx+JxiCI9nQIx5/+6XLk8tz0EtuRYj65OSSX
Mbzp8GoCMVH8qU6h6riRtFFRnB/H3SFjQUdmWY+J4egpkswE9RXQpjjogH3K726Q
KNhlkdu73UHMOhk94Ato92otval11a/k04Z2IIuwbG3wiJGmuTh9DuRSlnWVBfX2
2YL7rVrgjT/RpOh3/b6BD4CrpWJdkVA+18IckJgEWxuizYe1vIFFe8VqNr7Nhpuh
0KLE3v1LJfTaswh7fDS7uIcwSihi5rc6NjtZja03yZscM/KGaaZk4t8eT2pF46mI
FG2EOeybKbwJ7/PQ5AAG3CuxXBRKoWYAVp+JIKoESq2dsrXi15NIgtA+72Uk8N2i
7HQAxXbXJeSl4V6vo2+0gkEsxDPpsd4vxd0U1rUTtgoSZqrSKfOKD5NR0fHxaa8l
Tm5zLMorFlh1EoKQCvlFY/JZsgJsk+yy9M0yThC9CMMpYPYo4gG4Ode+ys3k0Ubg
84qy0tV83TRNOel9rS2Bt4+vVtZ9t4NpMrtYDJsQNQkmcfHHoDwMShOQBxktGEYc
9U87kz35YVv7HgEQ4td/wVJmSPrD5vXqM3tWuGpS+XYtnbdkAMI8oTYbVwGIq2nN
mB1LgkqNcPJTLxxNljeZ4/va1HQeSLLSZG7ZhciM+gmUOjXiAn2kMIavOroQdzLx
JoNTTYtsNFaBwiaKerajsncXDH9u1ePFYAxWxSFgUuSuwG/MpbuIsDn6Zk+6kHsS
eiNfLDKKBkFDqT/U5GEo29ZXppx6BnWF3aHG6QN122XX8twSEpjpJx2jsPNzrCOs
Nr1gC8pzWxUWjHxT7uVxik4WpioeRy0S/MFgfaShfSdr1WqylIyjAf5V6EkptWCg
1TiR6oxMHifJ/ubsb/vJyRoSM/YPY7WRElsUXor2Xpz4KkpmM/b0hppLh6yX0GOH
p15wTJ5oMzhOpU5TGKfystXd3dFPFYoHyFgAlKnS4DLAohkR5mxnjJQJ6r9PW4GS
47delr6DCinX2HS8vDvr7iLGCHccA1aw3sm1YaKvTsDiO0tQWRBwOkG4BMV6zs86
PFsqru+9sJ45AsBbOKqH1s+NuArjz2ibFu6+wkd3zK4BHdOYhzP8i2fC1AndRPOC
bto2UcHdHfWUDWmq+cw600t+SrtjSbBKrCWsLBRP+mPAw2YHMmNgLTY231sr6I5H
AL0muk7I3AdYthyVIw5h4qS/0yFQRwhmniJomQ/h9h4UJZ8qdzy5RA4/1mSa2hER
CdpVb9YoBZ/D74aKWS7mgOSUvXujwbsPDsjFF3mm7QNC4L/ZtKTopZRUq4UOn90z
CMmIwDViW7n42iIEG6nEh9bNCkReDQ/GHgIks3Y+2AdYbojkBxEs80CdjlSiA5KH
s9X0YB3A/n9Ksln007qU8qnC/XoqfcRrrlk6VlhAc1ALWF0WP6gHd8jLQbXtUUS+
gHogrT8ajUxVXYmNGI7BMNGKl/dGxK3CnVS3J6jmiWiii7VhxNJvIl3Xev502AfD
qyGMGXRQSrfzU+YXN4Sh5d/ra/7ga8f5W67C7VHL7AFBo7eqBckCGzpDaBddltqI
jI79AuJAwSkZBmobhS7hEbSV4oRkoan+g6yzIWAdOpTaw7ZdqV/g/NOaJM2MEjYm
FRjxMvMdjmFdgszjSr4FTmnjwhbSaKrXYoY53PD05U7hHtKkWZLC1YFYt9ugXGKD
rz8bNetsua9tLe0hyFwDVUW5nqLPeg3eo1F1Ym93Lhbv9Mv3zxcHQODtMne9sk3K
S1Xi/Bq8VfmoyAV8ZVLm+Pn24aqNhZj/qzN8aTRBiC9dSBvliJiIMog5l2L+tuGC
tTwROG2hO3u3h3+rO98nlViN36t21Jzk4JhfBai0/rFpdJQy9Fu49ulo5xp+9gfA
Vln6YDdOOn+8rsfT+YVUE9JOYnaeNCX/frPHGMiRmmwHZE+7KcjcbC6/6/eM7rV6
3qvRsLE04y0OJG5N8HJ09dAI9psSrzMOeXJ6NH1B2SzCjbLrx81rHKXHqmEPJIpO
/w6KrVtGEYzlKLWJ2QSq50gyG1SVQSZkM6w4YTQgMfIPqXHRUFEsWgHlCOMjv/uD
UyVQDbPaUTJA1lDZFJyb9qA4oiWx7xw4WRuSXnrhQw0U4Gr+hNDFGwFJDBJBIshw
HHva82s5A7t807bsccin+2FcnOMlo7aC2R1l9R9585nF3BpwcUcRifMiHQvx8IIk
6LNqWRtuLsPUEiqE0c+tSr71RlOiIMjwHqC0wsfX/d61IctPO0q43tdMtxsH6gq4
7VlNegU9TWJ8b04NXoiG/ocTG2s2MgUome0y903F+SXYaI/C2Ew8NC/BnZwuCpkC
U2oqrwjqRp2n6dthCdOVJDF6Met+X+Mickfx6PWUE2qKbZcFLmPMH1kl2EcM67xk
PG95z1UknaXclwUBm4wC5UL+MZWFbKFwuOKPsqWUx5iNn0w9SruwtgOye1oI+XmS
S8S0MoLSYVBVQ60W8j264m730INYDH4m2YNwYPv5BqYdnL6Ur2797PP1595lV0Wz
6t4hmJhf21UyecS7sekahbz9HFqOYxw8bX8IlnvIDiXFYnpIDzVo7HcVHu/NLS0S
YOdYvX+jzoDMrXIi7W9EBEHDvqW7giWRPPsCfcrLjj3lp6H/+zH5vZGdjKHTT9e/
FjS8Ad64XfQqmziUOpbmqo4KFb692rVgronstPiFB0JKDOuamfsOF9FiLETFOZBY
4UjQmY0m2Y+5y007+sdfAMn0jfnnG2q6xa+fGLyjZ7jzwAQ4kwbfaNv/29VlD5wc
Cq9MVVGJpYXZdolzLvM8W9YGKP03X33oGqX9u3pGTqWeiO2BjCex/QrvuQtc+FIR
VDJEiV+O3bd6ZW0ffbrLW8PFCV6huUgseRgglokl3ibHI5weAx/K9MPLRTc9fsnl
M6by/wPXVmubE+aDZV0jpCBixWyOa45eV7m1bBf0WMtvR9SrOkKcRty+oksZv4yi
qYs14lL9IakQfvylsFtiN57y2iAzf0z7p+HX7WWJCs99xME3fpOcMm2XiQVRk74X
K6r4aB098cXPKJAtNTcaCDp3Z+AhGVse+uDK34Cxt/x+N75s+3etSNCFV366kaSv
eBUwKguHxyGV87Zx071YJ38POUKKvSclJWN7/PJAa0tQ4+6/AGEIRIEAxZG2+fnv
4/a376G3PhZeBQ5NtEOsJ44NJ2D6LSCUEagdzbD0l4WvMVesHfWaCjBaczl2pSXT
ZMOLO2+m73gWLFgO95JmZ+8QoTQjQ4BPu79NNBzyWqFWSQ5+dKeRbYX8R/L2l4SB
2DbLPuRo07kGul4EoEmzkBLPf0nRp/QYPA+JCwsWSkQ3TB4n2uqV1o8CpHxq3sA1
e87ob6vZkyqUIFjzfoCj6KI3ulJDrYbwyr7oVve1kgOn8L7kcvDMK19mowPnlIva
gsUBTTd1Jigoda5h1sPA373fsydcJDPqGTKJu5vwkFRMvorMrDBG5L8odTdYbd9z
RmSlwg2cnWG84pH3boc7iqv8m/0I0oUJ/4mRDkkV9zgfpnifdkZExO38rxvvp8vr
yuEsVfB1gSWnWFxbzIDdu0YP0PFe9F8fxA6MO7w1b4I3ije3nJChAnx18MuPZpgi
mSWPysDIobbqeqPAWme+A+HEEVEg6IRz6Bo4qVpMVAiF/G4oTCCAzO/EKGNwr0NW
eqDo7JEvjSKclePy1HH2KXpU1DZKyKRVXGlJFW1RjCnYmi2N5K9fQ9AcHyKOuPty
393yA3EsAqjXbbrHiBgahPmTx2+KJQtMZFB2EaOdPXdARc3DVTf1XLP9dCZ1P2+X
FYpyvdBQ2Kqwoor+Mbpj3dgMz8L4lJVNSDLQ8/wmUpcMwV1ad/sxai0qaceSrSmA
j2ar5d4VypC8ecS8FLb0eSVipmRaRdDTH3YEspjZahRORO+VHr9ydKvBL6DYZQPH
QaLf6B8yOqYULeX9SxxFYD7dv2jCLIRB3CWBQS0zpnIm62WniNUUNUv7qI5Zja8N
MTYn5JBzP5VLu96BRUpEXE7I6xrf/FXFRY4502SS8rFGpSwHe+GjH3UAuXdAvkGU
1HOmqBMwraLp2e7+P4wLnIcfIZBcBkHz4OGHD+l/gI6xFTRVzRc3ljJUEnB1rfsg
r6AWLKM+XRpoHI6hB2WFEMF+0olKHIp6g1RDLgjUMD/NQDKiVQfYQ00CTDmXAKl0
mNLkMpZVS5LcbW4qLbEKFpZJx1upi653apbEo1V2DrNnn0zWwVZ1QFw0VUwB6Xol
UbxgzAF7SydEf8rPC+7Mbz/KgxTvtupJJgxcIVaxYcDFd1/adwGY2U4y4F6KR1zH
3Yr0hFoEHplCz2wZ4PWwK784XVUugmJc9yhO3/ZER1tZsQzpkFayC9oVi+GDmqIH
z87OFD1gi3ih1pEe66y3/jxt0tfuz7AeNgV0p7AtnFZibadljHHlY9wGjdoLopsK
tbjBMqda2H1fmcHgVYouSGqLWP8G6VXXF0d8ClspNKzkDI02O6Btj7877KCsHRf5
C1+Xim2toh0EUBardx55w4ljq//W3U3ayH7EmX+bKzrxJvtAghan17LfW3d7VAbA
NWgtJpkZKa/SvyIV9cg2dYKFif/SuqD62Ym2fJOHlGbhzms7M3c29H80b+Hab7n6
MQTPqy54MWCUWZt/wVFXmLo9HvnOFJ4Fy56aGJ9fzyGa3mv35GgzkePWXGj/iUFs
PfSOIoljAaFUv9qSoRwbN79msfw04FrJRgmyiYPucTxWeYKQVo4OuhPcDY8jxrlM
YAcqQdNo80xkM+wfBiUBfB2TKhb9r2pe3vfiRrLZWc8lWemLoQ2FCsIwZlAjvvMU
wo9XzgLshbEawOF9wf6eFOhvzOFEyY2YD4fhmd4KCRbzVo4AFmEANZU+IwMcvtZ4
7N6q1UH1M5gmI64antH4432bIRNSsOh/DD+a0Up492AVwlpvq9p/MmkZ0IpVd3O4
6IeGDwWOGkRicwfBvfrz7XcnsgoSXSjAEJynWuzMe2giHHb8ZawM629iwqR1ACTF
RzgDijX+ENScQwgM6XO9LltyhVj1pXuyt5nRp2LMAINUs3XRO+N+JxPcSOU27msN
Tu7MCw6lFNY3wNNjCheKvqWa6SIV2X5qVbCxc14YCvXWYDEp2m8h52TNrKzUDdm3
mnZ7CerWT4CDqoNF5rqhuB0dCNNi+z2QYZkltrvlZatXl4VBHko5QR+8WWHfO7t2
B39L6rG6Hg0vnqkv9JYuDp8euoqWiHZB2jULFEBlZ9eiGMF/S6PQFgEYpt/1Qs7F
WPntRnzTOqK3KMRi3xl0EQ5eOFb6Q8jjwJtFBHC1OXUHdnb+7J/M9oOgXCrJbKCq
aZuvjhb6/ngAlbYV6JIren2VKw7vE9vDPOndex9zvk0u3QJRQePJ7kj8zldgHi1O
NvhBC5IUP+Almxo/GItJzMqyCPCseMHESTZqLBREn2FTnqSG9Z+VKOFgGbrs1d3k
9sklLd8SMlhalEddNaltiQ+JqwVdhnMV8D78ZwWnCTRrsS4fo5TvhVvjScvnucZR
M/DgE/rt8lzxPyETJqqnjq8CtCaD1tcVQ5PNKsFKFtzuOrDn7uBTM5C2uAVq7kh/
4Wm19sMzN0aMXJ4x/dKnrxU18m3OeYIZm6MT2gDHME3ER7qmapn+H+OSwM5XkAM2
jzQYCkyKcRI3vKwZo+/XQoG20w/dljQ4zxD6aO5uGl1rHI3XvN83IEaSaTzW6nJZ
PriCV9kaDzLXbccp1EYBj65wYXyKsfBypA5HuJ7DF+5zMBjFL2HHBYzxlI7JU2Bq
AxkxkRv5uxFGSj9ChujlO5d9yh+viWlqxk2v3BZIqaZgYi0f95u9OeoocBPxzNnI
s6iFvLtbCtWkYTHwsr3gMDJVfIsCfLCFWgSQgm9IaHHECUUY3+OvmIs4ecbG3/PF
y5gQ+KM6nHEjc01XQedbEf5ztHEZheXPA8/hILNt+GR8oFV6XiZzrMKZeCEaxQGS
B6dO+iR/n2xuM/6KM6HVhSyC+wgUUjNW3u6FQUX1yekhHqznBuU7o1slJ8dOcB7L
gb0CFniSEKGRt19U7amHRm1pFu63oluACcjnPHGi+Wy5g0xsMAp8XZa5RbHehSst
5STq3OW/Q8gwuDhJr42maLpiu8r1RyxL2a3KwUI9JzoTNzrgY1H3KSlSPaHRSaN8
wBAJ2/0LVgBsYb5ApaWBV7hU1gpXFoYq/1ucSGB2mmcXkyBuBRfoNZK5u0gHIs3P
uvMwCfTQo0HzMWTGl5dN26CRqdSyYjIkZLzzu131ybyhN6JMWFgyn5s4vh1mHcCZ
q9e9zcC3b1uE48fI0b94NKijsS3rJtijYAq9vR/QQ/xlkYWHOLZVhYCaePmun5rT
8umd4FIdpuL1KTtHossVjGtOVkDy8/xH3FWE92jTckaBfOMmMsX7ZhKhGT/YDqEN
o6owXCwW2+MRWRODe6GGFnTaQnWPrdH6F1G+sQIY452kA6YJ4q7N3o0ImbxPyRJu
c5joTYJWyA448WtUNZIMcG2ed6o2ONW8TM/2W35wUqoO/6yCLcR5ThiSvZ2PKuTG
WTBPeWTBEQWAS3WpVdo491xY5SOiOdWEM8km0Fl3293bO0JrUkV/qXnvGuZI0WEw
f/RlpcnClVzhngHdtV8qsKKy1/ULrV3N5dtJTLYlKlh99pHCby0O9VsqsLM8jNVq
+O41Eo1PxjDlOi425mlFc6tlSDrZ1TmTYOC/uAeLEpTx0GadPz/OCTUeqJgc0ngj
c/s3S5pQjuAfxwefvHDNiFKxta6VXNjbeGyct1kqe+09M9/uFZqRuvclW04tLBvj
aiKQhWfHPI+e5l507CWS8H8I4AePXRfRRT/flF4EHRMKZ6WVb88R+XmfTjlGzJVr
uk/sMnasMYaa7RunCRCyxWJ7kgo7qEZxZnSNCOnxV2H4y2zt1L1yKwv6uC75b5Bm
MxtPd+mlsf/g963DhX0ULuA5hgvMsboKwGsVX88yRQo0kbRpqcrl3pYhg4H3FEWE
Zwmj15v4/gMts5dPIkAHjyWHCes9HxLf/7zq0jGL7LRsgXYo6ZYS80kkdeHRrvPP
ks/94nmJYBF7KQIOG4XleFtVAYRY6N/toCEXjad08fo7pAcvnsuEwJdIwZy+GgDf
jkvTLzc3331PCGFeBCpYQRAOrIm9H8Fj8/fjy2VE/jHhNcdNtslFA263Q/PMW5hn
EMOKW1saj5VwnLx6a4mux5oUG8gIFJylXMgq1GjX8uhm8gihF34oFkay2vFHhMis
fEmPH30qn1dMnPQ4gI3NBiReg0DvRj9B4KXmw1YQyGaJ9jqe/6KXVeI3h29OAj/m
kTer7FRuAnc2WGL2W99Oe+9EttzqJaNg4g83X2WPMpDAikgw/n6BxV7pW+GyrOm9
TvaMR6xJIiZOPYmatGFStEujkNezzjGcIcHGdpq+ZEuBTLSLIznzQUxpS0brKrAl
ztsNJal7DIJeYwXjMqRfj7Vfdjn/4y2D9MQor4dJiFVBkZQBYKgjKoDGb24l0MH4
Xqih3IasOMUYiO1ZZcZWuWtK5xt4f4cJrjQFKlvIY37TzB9sBIr3LNef2Z1zHbU3
QxeDBuk86i/VxOyZrFlTXKlay95NzvMbeG9BRnr2J+sEqilAgiQVW6xq93xKTeax
6PCzppRrSwhOCLZ7UZG+rrADWeddc7n+MXFoL9gyxD2HfXp6yvOLft5IdJBCH0ta
uK1lXoxBHmkdOpb4P5kMUEqMg7wASYb/LZT+o1Cv8n4MKGPTG/RyZjmrQhIzxm8a
2L+oi1uqLRKN9jOCkelJWI1Swb2d0HzLVloisKLRZWqzca8r3zhXkrDXX39gtTBv
AcQ3Q/se028UutExdxrDI1ik4iNWy6p7+qB9/6vVyRO8/6AUxLjFYApqCZwAo2nC
QNOuv9GBD3Hj0FV+vZGw6eCwGIclyjXuC8i39n+DUjHCYxA7UTAQhj7VM49NFhVA
0Q500JaFPMcqY7NH8nKLh/Nd263NCZmtDmy92ExKjzZZyeWIcRid20JwFRZyAS6b
hqNd9ISbF07CJatKAdL1rtp0Q4+tc5ziToW3l02XC6xBvQXo7F4JkK3tuuti4ae1
CJKAL68rzyTyyLbAUdRvy09vvEqc8fHS/9QSn5cAXpcJB44VfZ7a4C5cXu/VP1rd
Jrcmi4r5oxd/edk/zcfDJFz39xO1fc6B+VQyeIs3zdY6ZM56TYnN4I+hUYgtIw+H
RXic7pKgESTGTOoG4mTU+KOEalLSwKcPDgB6rF1w5DycAjvMX19L98M92XUSF6TS
Btr2dwARW3YHK90zz3zhgTSRXV6wevTt+FRMlZPJYnVJQ7rn4znQxScnmvzVMfiV
0brkaC7EEhU2FO0ngI/nB+BHxdQ3ucHL0sCUvPm2/tP9SGMPPIJ25Py/HGQVUfJw
NAjr0cVYIKjunlxSCpv6wBmX1TzEWQuknCh79/3a1QKiNkE/+bd/IigHqMdw8VVh
2kKzE6c6u6Gmp6H65KIacDORo7CUZpWjiw0bMPfQTc+WlRCoZAfYS+z/W2EpnsAV
i0GJd5M+FIzXP1TYXHOgD7YpV4yUw2kfuUeWYfcyhOdXL+jY7EzmpHjRDRJcDVp1
SIfCtebUKnekp0Sp8gvtO7MEYnh6aMoHE9sLVIyQjFOhdasu3PIEaL0lvlqk6iXn
qlkcJg0iJ4EPjVAwGvXSjTSSpZyXrTcx9Kd5EQ/oTS9GlSLFW84/cgRtvoYjlHMc
qXV/YJDHMi6roMcGJVvsdnlV2v5u68FKYqfib9Yec9451cEVzQ8wYba8yi2PEXKc
VN+lEisII6E3O1cSyTt+20zCrZkpcBQps8r8HCFdGW6l7tJYunbtm/xXf1154QZY
w74jZ6oharPTs8YMmFXjru/Ghn493cmucBFQfD8zSmWBTrK8FjDode3YLlGD3c5b
IN3JAnYjpUQJFsOrMIy3chPItx/C/AMgwZDd4OxEd6KACwWhmcUKkTTln8n/IMNd
Fp3Y+5wxeq+C7I/L4KtzKkQQQ8a4yZlr9dw3p3hpkFDL2O4Pa3m/TSxV1hsEySEx
zogVf4StoPtw/wSBZrD6AqS4ihWv5qfsUlAq+SqXfFxcfitHSAyuoOpTJ6Msi4rM
Bztw3ofhHxSemt5kidA3Zlv0L7vAnRDPjh0Le+DbcaZkIZ2ANIudERUuBHi8ALJk
QN4MnmYNs/g8o0RBvws2fRHxuJjgGdAyO8Z6QjyPoj3KDRyaHgKV38pWQSTEdtsx
x55fPtTOF9wWCK3qN0FkevB7rO0zET45431BQ358UH3HzKru0genVWf7qTaKD+EB
waCMEghEV5FbWuStG6SeP8lHvl8zCvEgdRQOvuE5ncirhtJkDfPDTrju2l66u13f
QcsJONEzqDYsVaoy5+RpHTkK2D7YhqnkLCmGMzNo1ASKd8lvTXsT5tVIidQdlsWO
5WG5jOU+2F6SRSIkvNDy4ROxycVd/Xo9LQYaeMwXE7D/Ttc/GSSF1FvkwlLc8z4W
TbZhmqT0Lc4V8iE1RZcKufEVvtaL8EtXo6CZB758uc+RVsyGzmQnovQjosVAjWzx
WyqEAKRuouWoc5eHm/fETGULX7H5Tk5ysi9IjoZf1Uk7BXrPoosUXAhVQm03zjfM
B939xO09SvUKcDljnyty+CIKJ1kcUutxCb6mO2GnGfqRmc4CyKCEtznauzUetJGx
+372PrrdBjCnsnndKK4cge790w0xBp1x/Wzc107YDuCxqewsPdZ297LE6ee1so/e
LRyJEyzw9sjmDokpAHZvapj5OP9D4qzXdjWx67m9B8YLxnEoBVTAyvusdKu+WMZ2
meeTmQeTJfLxzTXTEyHNF7b1MLXwfsr4+Q+nkGQFOoMNK25OPt9NVp+jlHvnbRl2
ItGqf8TW5FPV/DQX9K1b/p1EJkeohgtWuFttrrkqcYUgpgO7c+ddVIY3y6LnrdMX
AIUqEEoMxAwNjvOHG5uo/VAB2Fpxv+WuHgWMKrc81eeU0LEE/fonVPDY2WcheByI
kN4CLlTnnfG1sd54XVdRv/kfq5wJCYlAlIG9NON+aVxWx5uI649E8ScH3Y8MjNgo
svI3iD3+sbaid54HDhtUyoz2kFa1wvufeYT0y3F1w1zqBghshHzZjBstMV/A1Ieq
3vdvqDkD86YTKq+hbmlm45hhkYYBMHgwRQ2J/eaH80tAq/xNaNvOwa2VETufQ7+G
b+k1mel8qEZsElXb77oWbaA2JB5STipx/XtfJoYrGnkzfapUm1oVKWZdmLB9POKs
Nn9eH+Oo+mmbeAly/k3jCJETbPGQNv7C0FaDcKzmYxxuC6tpBgbK0dqhqABzcdkA
rj6la/K0kG+AMSGtAYmv3BHqmUr8920YPFrtFjrovxECxf+B+BXZFviqkoEpteET
8lo8LBryPybeGSgkWisliNZ1TNxLzb/rsq2vEuPzLp2i3uB0TOffEAoVOkrd3mY+
JUA2GG7cH81jsg37Ada7kF2ZkaaSPB/sQAoOlzVhC+aM4/uDlq4C6+tSZ7cYxECo
iqAuWLmldq9uW1N8buV1FSyP0A44QlPh9z1hlOF+IoCjwGqPpUAjXCLbsP/21378
7ixrQE1hyDXzlYd8R1whPBM53gNU931ofrMsmOV5L8+/qIjBOvRssIUsOwDFoqS0
oKcaXcYXUXELrJVOf/cNL2U1CZVpR5jfyNSCJ3FJ+/ZUEveKrHMxEG6m4jWTH6dh
3nnEqh5TGnAeBW/DpIwDVUFH7pgjJ+QsTnMKQLsdyHw0YWOrkvq35MIeDGjVDGUy
l7ndkdshcKKNAZFonc17Co0Il825Ps1u1QuZqF5gLGaxCNViDHqn2h7P0o2oZLjy
1JJJgD2cy8Se3k/FjgG45qSHoqhIecIUHa24PM9Zlx2Zq5Os7xCpROKGCqIIMLF6
pS52TMeARxiW2KcLhzURRKKk7JszDjIl6kflumrsCPpUCEWH6u03jA+GM/4HgzG4
pOgtqBkDY5J8eZAhKkDzi9MWFGCGydKz+7WcqV0mYX6G6r22H1X5U0v4e2TDFldw
meRl6KVGtAERFX9SNnCSuk5csPP+9Zjx0nhIdQL0moYSM0TY/Zn0ximvfnmRVo6F
KaLu33LgR7YV6O7c3GYgK4p+Zdj46/lOy7ld1l9JUZEkol42jkeagYaq6nltyLzl
dN7rpoQCc5EV51kCQjwd8ELWwHXWRp8bR2AP0BimXT+4Fk/4/ViOJKXLbtnN/Z6c
QXOzw5GqdMowxfj8Gvmgoxlzq3S3lB7ZuPT5ioHTRQulZvmj3CjyvVWxEbNmoW7j
bLPsdmGL2dF4mhUMuOiLVJYHBDCfyHtwNpP+hZmuv2c8fC14mTgLS+TeIsJ4/H29
VuwbOPqECjg8jymmffVBkqv7qtuLJH6rkqkqxpuPdCSjK+lYU39Ew/I6UKTBxiLm
eOAR2LV80+WyLJ8Qf+myb696NOnO78NMI5rffUBWZMwj7B8uNmJxkMOqJLsmm5lI
7UpcNfxmvUKlCWYAnkG+yoGF2K+nVVqXRGTCWpgm0qnAzcsNxicIw6HuQSfYC0P3
r/Qgxit3hKNeaEYd6TZxGj5LlV1ApHmdoHhpejqOyCoAYDmReRJYj/uePW4m4z0N
1jv5C/imqIdR9Q8yhdY9g7KeO0DovuaPGqVT7Plj/jelToKhsHwwXxMNv2Vc59zV
2SUXM6nCwRji6JGIzAENf9G4X0LqMK2W9RMNPeVqa6BlfMFsyNV5n55sMfQzlJmB
oRpCvpoYLpgN9ZwlFbs4TRyNBLk9+5JuvWkpuX0HFRpgNNKb10ZkhtD6+C64Poc6
LlXCjm4dI4UsUnt92EacV9fiKw/Ztb0YIwZd6pS6J5eXb+wCFnlLB/CsLkbtemhx
j3SEQFz9DzL9usEL67imXJy2Q5e7RbaPnkfld3uGQ0JvZxNpXzQdlorUoMFO9dZw
GQUVA/iNRKzE5H5YYj0pMk9ilQ3yfNSlgN/fYqnSXXbJTyBqVtvhVEsGGKKCT8tX
lZdlDBa0IWhOTbsOLa9sgbH/7Nf75RXJ1A6iJTMJejrF4Svma3w8PTI3VZcycduz
LgVzQOffyjupQUWnz5i0GxMCAJZdMUZ1kcQ9iS3X1wO6qLvIb5nXVGVxO4z3hrmV
RsS+Xsf/wIhyPW2P0BxqhMQ76lsdEgz6WjppNzs0Z2RwKidFOe7eMUfgyIKJqrUO
+cVN4SeXq3a8SR7lTQV+do6qCRMHPGitots7J0PCW/lNQAUZ/iEWyqCsR5uwfFhf
52G0PD9yj0hxk8F354fSb6MKQ7pncgdceQkhecHCFCheJVrTTS29huo0ApYnzny5
UDhSYaV2LuvJ8OzU937dTxkEZPmjLYF3FgUs3v2L1NYNy5cBtkN6CXcEWXID5DJE
aN/GlZn+Y8X14sMHSGJ/tjZm5ZWfpMD/av56ADrtJZqWQg0Te3Rc2aSWjJblwOPC
RCBSQ7IIBO2QYTQPApC5Yz7UTdhxV3br5FoFiJBYTcG+VtehiRIOdBbkPKBZaP5j
iGkZqrfMPm//cZOqfa571YDoFlzkt9zSI3HP+ftpvkU1g5HFo2PH/byNeFEmaRNq
6WTLSAVr+3iMNvTGlSLQmDGHQomrgqUNf1/GeViwLDLYBSxtEHIl9C/l/B424AsC
ALl2w+lVxzcspqGP1GH+3HZfm5z5pJ83TVNzvC5Agkj3dnB/q/bFLH2ZzRDWy+BT
rAGzIupza5iNFw8O+YGc6okcEErvqwJKWdu8gKKaNk+uw59lD/NJdQX7BAyTdR1N
EyiJHuJEEBZqCA46wOB2l5H0mEfDY+rum6Qk8uEtTfLDjKDgZB6diW1MOqC1rL2X
343Fqrw6N19YkqzSe1VnUAZI7vMJZtBadup/t/i5e0mX009wgSvjGVZqcylA1Dpo
I3aULq940yh0XCXuNvLALgJXJMTX3rSSCjNZK1v7LXO3DUyHgN2uUF2aLxQo2a9s
+bGeNPrf1poqDIcIM1DuyOWYZ6Mp57DrSsaYTd9DWHO1SPfSuSyNNMXQjFZF5icy
94NjN16yd8NBsRWHpFj8CWERL0VcjlebYYz7ibXmEYd1Z1wiDKZ+/ZVDEmMsH4Ko
NITnj34zrx3g6ZBW4tcdWCs7tNWVzha0GrCsTR4VNxxgEXwP53+qC506+HAYq03a
uFdzStJYUaYoGEzTXRQ3/iAv+Yi6s4T9u11BZc1ooHRvMkBxDaIENDTXAkIQHwby
HsaiX+gWX1SoIPMDhTGmHM4QIYVDJd2HnXU4kEJ+fCv2j/1PvjLislq+L98RVW2W
OmPdj/A/nuX3JAHboP6mzGunNeTD68iJXenHaFmLr5UFivXymnTpCHGfjCpg3oxO
BczBcPNdUDlc/c2Oo2PsY6fydmUwo1AXd6JAUQ2uEHx5VPRkSoihHfx1CkuSf8TK
9tBiv8Y1JU8208Iihq1NkR9IHhDl2mgITgJ0Dd4ItjlfP2KY0iFgD8D6F9EBrhb5
Ksj7rfo/v4PtqSajsqgLpgu+sHs/H1JHxxtscnPoinBUD8VbKAlAH6v6ekmfcIrr
ZvLT5LpXMHar85AqPNZV/XqjKDd3oWDpOxPtc2ZAmkGPXNzfXV3Rqsem82xj566o
Un/zKbdr7wI/zKIY9UnNkqpA/2+mLTQXKVTLXcilxh2qcI/MFD55qX+v9qcImbSz
SWkP8s6W3CZit1Ja+bqPSf4ZFuhc5iqjUqIweQWnQVQ1VrIvcKf+BU2KbcZewVVg
n+AQS+LsGBLEzzhqbqo5fjMQk23ZDi0YdN9TdI4PngeXUX53/2Zkeab356OH79ny
WhgFnGLAeyRIsHmrODpi43iLJQvqQPUCDLaOWvVI9dQfql+Y/9sxNTtQm/9latu8
0+w7J9Vkf2nb/OETgckuLePHpEo7yNgUEOyqnIBqJCF7oEEP9etZNBKzVFTqIYvH
l5jejZBRoZQ0Eo+JmhgtrgGEDtV1yKV1YPlO5XtFBQMdhHumdfkht+JmFxKaZc04
ni25Ol0iZMD0hcRJ+djter59q1azZypGbh19dO+frbu2/q2UUJbogxae8NuPM/F/
i7edHkMAQY1jZhHMhn7PcFQ60BQ0oPQ7kYZnoabgpwDePgPq2YyNUPc3on3gQXdj
jXhl+goWBTefpp9AnXzx19Y57lT2o4/LcIwGMwtOsJ/YbNk9DGtvDnv+Xh0GDPm6
Z11iDKnUJnZrHkGAQhK9StGRxDVVuK5z6tqVuSR+p9rD7otlZD25L6uVjg6i9xqS
mfkZ6ALlUesijvpfjpQhmjeY/fR/fDg51blCq8qeJvdKFPd7FRCmSFbRGv1Uzk5P
zZ6ehWc9vhK8+fZlYO5acMx96hu06RL24osaV+CNHGO5DHBaYkKPeVUDA3ayicgC
HgnzqWR/LWPs4UZVMZZuJLAKIVgSfFIVsN9P80FyB8Y6hMTmr2SwMTjA93CXxMP7
NycLqX4BPBk1eisisAg5SDnvEIpiodAqtC8gQ7IBRCk4S73iPaV4NfTGxAbyM4gT
If7q3Olkg7yJObDh3elxDkN1yRENBJngjRIaj/TndsKFoM2lhok0/cTz2Mxm2zF9
544oVevawdDw4gtH1QQFRcpWAl7bYZrHwgOL9NhwcKf/5FfHx1kecWMyI4IZR3qc
d2huocIT+VdM1zKLn2JuEEvPf7n9V6shgSA2w+LFIPQ+0APTFNc/vcnK36TuwRnM
qWfblW/b6O7Q9Sn2f8Hu/4Kl+GmhdVvayd3SRiI34OqZNlMlNReYtjX7AwLp5tSZ
jfTGdYtU25i/BBoy/BCd82VfUVAH5iLmYsgbWl4tuDPL9Ez61OcoLkSFURgRqdVY
En19zlvHccGqEmnL0ZIduHDX1oslF7UYHZVucN4AfERlbXdmk5vE+lz/CB2BiJKw
EePdwZHdZefCa66blzWvdpRuXNms4lEK9fYCFN+gI1HX1JCh4ZaGVCbaoBSi1PiB
/E/zEJhkH2dKl5htHtju8gmsn37An9xRyDi42n+Q+44t4ZFAdCirQh0arhG4BEOi
Ef/eUfDc60UIl9W19xcPSn2+X6uMGcmRZUdvPI71SyrLPEPr1S17bvNiSj1e2oWm
hlrK5VESVyOCkn7RmJTWd2MQLfCRAIKN+WWhWgo6tPx9ekSWE2+iSfvX+ya3xoHz
+ett4mWufTOsEg17eeR7JTqKvxY0j7Cb5erlNrNXrhXAfYbYBa8cTjaqmLX3Seoz
/rXjwynBkBW3OpAe5bkOAkEGELaYs0y5Q20FMSWlzpT80uZdN+4Mt6+t4xgCQFxm
8DhUAvfMkUwlSx7allxSUh+OD6J3e8FFwQ+b1pfWz+zaqTIUIL4OIdRNnyEpY8cV
GeHb5UWYrffDKWREL8GdDogPoYtfLRN0AVRxsScUYSpWC3MbYJNf2LPWAAJJtCTU
4ueIVu88opVSxTKwXGgceIf9kLT7/D1oO+w/GbEQN9wxEGj4JYSqFOgh9G2ZZa2H
3Vjh1IHDbl/hRnJHhHqolsxH250BlpaPZ0Xg81bDlYCdRyrQqyUghUlJh2knwGb1
ko4RgKNWZ8lk1278hQr4/QEKem3+7VfAoA98GYUhYnzOdpF5ynstmcp1yf202Vl+
cRVHhMvb9WeXsrMnnVyrewdjg7nKqe84H+k9Vnr21OBp2A3BlaMnGdmQ7ncgs1bd
NTbJRYBZIR5+CE8+8hscIZDMD5TX8lAimv0dphnjBOAbxDAqPBjRaZ50F9u1ciON
KMTyOHuBUQBqiB4LY7KqIusA0vSn/Z84xBY42k/6F513H9RYoo8HVH8EaD0Tjrus
IbRtFJC8t3HWMkwECO3jW+QXVtGZ7US/heUCZSRUiyXx3cWF4f2cgaifjxMdIph8
8TYDGlNJ7ipMibdHjhWns0YHbemvEY489GTi1N8Smle/VQV64V5VuYewxw/O/Chh
zD1uvsJcUhnTgXloAluOv/Fpe47PgIhUjQmg3eWhuwZOXxjEpoTFRF6fV2vaWs11
lqt6R0Gt7mWuuD8aG3jamnH5teLiNr8cn9319TB1UEEeCjza6qkMzbkiLLkG7GSQ
Ljb8XJQuAXjny1VPkJeiEXzqI/sVkvIjFw6sycOoSEDTlZS1KyaKO+OBDSFL6vrx
khG+5hKalUQiI7b3ifZ0M/8XAnSutREHzt+K2XyT8wrNxJpqTXsIl6xnjfTwRH7B
1h3J542kWnscQQX0sohA8Wk0eOt2COiAOO4Ha3H/JTp69JuKS9Mb98YqG9XfY2Ft
Rng+LuNRn21fEB6Q5hnz1wVwCEHZTJ/9BPz9hzI4ttc37QfpAAueMZ8LA9yJiSBk
mO4fdoEiXAEJyHFCHMr/eHfwG2VYfJ19tRuNzkYW+NRBGca+9RrlwdpB5Wd4NY7Y
JOARfrO+P2heJ/puHHS7G2IoR49mNq5kTybMTSv8+Bel8gWelK3HpjtHtsqdCmDv
Mvod6tXAvWBzK35GCuliwjbsho6dsAFfv9JbRxQDNfkCFKym9Ox+dC+TzQstRBtc
g5ilOmkSXvYDH9Uhl74vWiMeTTPcc5B9DfroA0+hH6zFuE1dJ+ZSwwKZnaiDzvs5
9u9iwehYSixGHbaEA/n8lMfWgcqq+6u6jv/IblMOzdVB028OeNbsI6yByWCXZn7K
eK2JJ0075icUh/PDXpGGWWEM7vcsNPT7U87XNFN/sLS1UHTvHKac65Vmt7/LKXf7
7BGhE2WZrO5g6/ZQOgCXwooDPZhyDzRWwxT3Z/qqdAJ4ha/u7WjaE5VoiDDXvg5H
ER0PJFEyA5tVwRwLwzGUfqOBSGUQFQ4fJSEpnRY+IQSqzRcyaZZq44HqUPD5u4xz
TiZT7tqiLFa/9F9mdBuraEZOlp0fQrDiB9N4E/lgf9X5Slxxd3mrQXzFDd+zXcgm
IQUaXVytldfjejSguOxq/OfM3k80aWAKJB420IyBTM2wm1KgubErtu5whYcsV37r
wn4rxDJcLChOKuvqJaVHq1chG0id4GXk/SdeQ7zdHItlxN+QjeNYQM9NGNX5vklx
B0ootg0NTWD1WFtXBxRngW8G8xtPSU2UxHUd9sGybxMg07eXLBt4R3SQqynJS4SM
8Cl2dS+5rakOkuZrX6ZT4rPjVe7JeFwYoeBzml0+BfoDs2fsYMedy78FhSbE1qHl
tqjPNiB9vTnkPqndavH4kptRWkQYBCWrPS/yDi2rycblkyHk2JHtspsCH7yKmP9w
7xiVerSSellBfsNHBye7f7IIBbFTP1n3i0C6uvCR0AeZp/nEzsl2jUCP8D7n86zK
Qw4nqFbgMzb1CPaozl2YLX9YVB4jSf25N7G1RCrI+GfvWpRxJoNIPnBQYAToTWOh
RNNKhPjoVKhzNXkzZOmI+wWL7r/giKdtP9iL4z5LTp0z5irrJ9ksG9nsaofKt6og
1o94pTVPrx5ZiKzxtwKjDVUibIyQHR+XVTT1gsvqbrDdTbU4Xf+yfhc87dwz5a5P
ZlSMWOanpPt9lghA1Lg/jUrlgTn5xkHoBwqozA+kI457zR+Pd34y0jiQbobJGRRh
ziWJwKZF1Iaaf+GyuSLdaephDr+EqBSJT852xHDMe2AmRs47EEUfCmG5meLnkLyd
YFbDYAILE1Ao5YaTZnNcM95bvtUlun0VgB8TJWZOpJ56jqYobPylwG0ahSMHxlUv
i3oTbGIqJnH88u8sRuwkv2gGpHpwb4XM24W6UroLdVBkhz0W8hgX6tsoMbLH1sHo
yqvXM8pJbQoKwYMcUi0sFxiI1D8y+p1TiYE1qsCPYbcSlFnqhu337WjS5HMRI0N3
9CemrBsThWuldVJ+0JWTo+EOCzi055jnAqseOo+Oznf2F6F1sKTghxqbOIHv1YNF
nicYs2nzej4b2ebd4LzJii5GzW87p+bHmblRxeeSpR5W5+QUBvgNgTo0YC8W30Cl
ry4SIkxVGOYynGbDOaGl9cvLyYkCgMbgkadnP/aRkWZKZSVPNvtZmTtT6Nl9RXNQ
QmZ9g5J+/Feb+bNElAH978fRznUcfDp8Ny5vLYqYtdpM+1lz+uGcWyvZrhLvgYy5
KhKrUGpA0qa1MoPVsn2rbF6e2TU253Ay5LCxekMMx0KONUJo3c7kR7E6jhKo6riu
cuqOgj0fTpgTYJxCyEwshho83OsEPxGTFMNcYRvSJDx+fbCb/XZRQD6FPPzpEUy2
4yqRdUAZelMWKHQgYL4cWkjzZgSr4FULTE3jnkTOIbcx7ZJjD5CJLetKi2v2/PaZ
uUx0cKrB1VJsv/OlYH8sC2jLVckgKcptjkuQ0Fs3OR3tDsgpIrwzAxLxhW/s+YC3
wF0e3irZ5ltn76M5GYWF39KSWsea/RCJbgZP3Gr4ckLKSa5ljkd1cPbdwQbea5Ij
1CZ66SlWGJvssDqAD3otSb13fY4ODPe8wyHjpeKembI/kmgP+WWO9vaN2gLkFvPu
mYQdO6tHHqu6MDfWAVxG8cK4NLveMt6TCGrNcCO9ZWjh+0NCzm+qbav5+K+i8Tm7
8RScBlltPEzav9p4Zn8TvBhConMZjhuDgTbjcVwIpL71EEirGHNzDMxylndqlD2q
wu6/DrxIEViT2n6i0kKYfs1sHsCjfk5Trcp/98NTzEmCHYF0XOrZSUUB/U02Q/69
8Gv6q7Yb03jOK8+5saJs1LdHmMxArAMG4tU9fL3nzhQErm1eYa9bifTezBXuf+mo
LjXHIZZQNnjC8E0pyvBQVGPiZ/npr2a88toFBAbhjO6nei5p08ucTP0NMXruQkiC
gXYxxZuF8mdwJ6a8i07HnC91yUPlCON94aGnnADhPYfD1HXibCo/eWNi3hvA9kbM
dv5hFliOWoCAzZdPuktXaPlcIqmEiNWTktRkXKqOSyie2l+XrC6ovO6N4tN0R092
UARFCyQ8XYmRKDrhZelOMh+dmPYOJd+xSUIRlJi6169KT93yKghW53aZtlw14YXk
+UhqXPvx8TV/Y91/iQ2e0zelJziiPw6neN9nkR+nGU69m34WhpQC0BAWovnnbg9h
0N60ZeK0r3QDtSMeuRsYW8TA0QZafUPgyczG+ty7YDi6jQa7CAjl5HcbTnpYOzQE
Ol/av8DFSSDwR63OQ7/SEDQ2ArCm1VpEPLRHdBZThC9XsEzuF6TpNqRaknOpPz9g
2y92FA2Kn/npvKhxYFutmXomARGCqRUC6Ex0XT2qficpU49U2I6Alk0258FBa71D
JYkp1CKKG//TD2s4LjVQ2VNBMATYwMricMSCifOanCz7GrCz3+uD67+FnXqyb/DT
KWo4p3WrEfxa2JHpJXeQ7yXFi48qiRuTBuUjYbdM0OwFqQ2FPDIs+kLCHmLsqaUm
ZQdDBeIeq0GeOmIbf66fQ3wEx/sBMbhyzTLlOhd4Ab8Xt898G+LF0/rPNuSq5DI+
N6v4kixzzqlg8AaUO0a+BUdG+j7ID6SFDbNgGjWPiy6CdnBLks2hlUegrMWEvp54
1ZZjsikb/TXZOueKWn9NCSLCdEu2ubqH3mgDiRO/9XIuJw3R9yqvBP2B0GoNhiX3
6/h74OAoJAALyq9rXmDJ7RfZtqHQin/EcOvwzQ0cV4lx401V0sT2w7xnY8NJwXIo
1tmiUmO5F0fLsdiTKJ51crhkFq1fDoQxjGzSD7oRNZBIeQPTxotJkbx2Q7s1uCnF
bUW8D572voiC3iwHRiPpxQwQL6l2/DmLbnlb0ebAjoTFZmTn9TTgiTqmrWrT0Gnl
kbcKEgH9aRW0s5eH5WejO10dOo/8pFO/c/abRiGWzm3z26rbPrBmOO61dFJb86ov
QVkYqcynmKYUe3LtG/8e1Vxw9DQ/+LCdAWOG57ij0H+h7MHlLJoDU1JEWdJx7/fw
jXaB8t4HhoO0ohCDN4hgjdeLA7/Ec8uHeDywvrnXd5H68a15c4JhLXfG1w73fhoO
Nl+M9VV5eTPpfYAaZsrYNWoothKB49EyU8H+G9amX8sC/s6WioEc2e0qDhmqAs37
+G5T9okphCt4xMevQ/oNvw2xFL8HZIpQ2lw8kqZ9HUjZgTFO1mKBeCiCZqGeQXIW
YYrw582n2y5cV3cjCX4ddHn1q0D4iGHjB1wM6Bu8oAebVosQKjyXuzUdVG9+vsOq
yRc7PPfAcrkLEgHc1FQrqzuY6K1E+MusZrBZ3vHr+wGtcmrYtUoUBhGrrb8gZOeG
zKAsUOP8BA7BV6fUNTilahMe1ztS46GqDVmW/HBISsFn75rOGz/zmReJL8ugSdQq
+7KcZzmB7HxlDM/FezSQ5GXGR+MQhIyYflRjixtByGZ15gkVv9oK0OLiyznx/Het
Mq0Dksh5Ao5Hin2qVHy4jDNlU2Vzl/EX0gWC1vy0xIOMahAV7bcS1UMvSBQ2WPi2
9aNPK8AeRVUh4JGPnDu/GNxFODrqincP1DBJn/bK7gsUyoPyHAi6JsFOnbm9iWuu
DZm8s32yLgC8GSyvL0JSMvAJ3o90nFPQVSJ5xruw3aNYkvKY3cT3aZJhN03gA57K
uOw4XTSPr3hS4kmNKCfvA/0ie7itYZAfxhW2Y+LqBz3xnkWFMtC3qpgqIwXP+/+I
+afGnMRpZgshTwn4SxcrZwa1f3INXtGj1BfZF9hJzHo23UCB6SKCsjNkwE7uq4Ii
M1JK2P/kaARKotkxLLitSvBFFRK68geQ5JTJaCJhEJr/FY7ylKF9/hWlk7upDXRW
UdBFTT/SW6s+pqS15XEyEoLpNhpHOEe1Jp2FwRl3G54AbYwYOHQNsiA1waW2wQCR
3vxgpyt6PFGtSNaVWzptHJwnMz6u/BzSncBmsQLxF+S+gyynSlTufVf/foG6h6qr
gxxSq35xSEHlzyrlY3/6J1uIIOKI6trtO1FgZNlgH7NzGDbwnhJWyOZU4DJZFCyB
dVH4oBLRrvEWBcC19lcpr6KHpEkbqxEufGDrDizqZoouy9//Nb5dTMGPWHq7RoUJ
NYL43eQSaJROpKDuXxg8Moir0TiEwHs+1z4dbl2h/QCDQl7OVBaTZcKZWcy9EygQ
JCth4Je54Chxug08LR96JuP4SdhWugSpcYgaHLA/Ikd6k6EGgpdDJx9osuQeAzxB
j7j2YbKqA3Iea/o8GMCTwkKZf5M6kPKNNH+yvXARUtkiQi4g/zuHX9gZwwEfekUp
cvQYHGfsLdG7QT6zQ8EmCqwVqZOTR4ajbmWNDtLG/AjJ0dmrMj1FEOrqPskf7Nzk
OpHkSv2B7PgTnWDpPdqYb6KWvvo4waszyvhhFGkakEEYZ9g4r+4UV//wH/2SJT1d
QlsybpTrVZNVFiWj+jAsZ5YGIWUQCJF7QJiG12Vyrxw73EFjoOtknbFSaecUpZ2C
ED412QP6CwIhYgQnA/PMj9hk5JE3fIL6jazHivP8zeLwPa9IV9Ll793R3y3UwQpI
2n7m1AUhcQK1S7XTtxCg+W4BrSAoTACkDAFsE0I/4bHMFhljbP3eJZ2eRmpx78B9
6e6Mdp8Kj0Q8tdRozmgy8nyZsBgQ0fsafUe95UoYr5ZBMtxOeU5u2AhltabBuZ5l
jpD48VYBomRVDJK5oh2tM8MnXIFJO223ggFDV/0xEPexHvufv75O7U4VU0skSt7B
uXW/AKFIrlOVlynqNCazeuA6l9XvVFNmEe4LouXljV8X1tcz+Fnw4CaJleACY0PI
TWZCuDkSj8BJyVYsPf3OfSicu3WrqcWSDx6ELyvo+50C+k6S43ebUjSb5ZkrlMaX
MbG7yMtOtduo6Ra3gGuUzD3Y5TBkMCAt2AwCZI1XJtvWqUJt6Jb5H9Xg8VPqYP/E
d5CtoXelRY9n+VJ8o2JkBJ8k1FjDNO4cETpQxGOExy8GetoNUCYppk3FDaaIOGCm
5b6BHsgXXYCjwvzXW8K2Vg/BqrXdg6yK5A/ZVGWiJEEOpUZLbrQXAD4VN2tqp9Zv
w5EdeOjAvPUlnvbQzWRxZST6O2WY5PcTyjkaw259JEJ1XSAoUdqYq2SsbIiUo9ku
2Fp+IdyOzXON/PUkGaYRPu6p6OicFM/Q8bI9cY64luKPZPTJtYRZVW04pLuL8XI7
pGwrkcGsM8jmBpHOOF7YIlK5Io++ThsypkgPjo8Me+scB3hPzBwM6a89mxmYeoIG
8J/6qCcWK7g0j1sVucWdWaXsZu2Qaa+SzsD/gTMiqUGEXcDCg0cR/V1ixAOR+lah
bkuiX09lSmMLFn4nMswCli2R7m83TnvwgTdeuQyXBGWCZPQ0mcJooMVI86BSxKwg
kvJSXuXmOORXmAjfJQNRfn4cDdyoCKaVX14WKBVbf76gGzNmTBvuuvIY03ZhN2ie
h2jM8jI46SdQGhKCMzSDyVvRhdNt3kwvfJe0x5/XYMY3uicYOlcUEYL18RctTf7q
aVVgAqqSRAUyHBop364xvtjae6CG2J/AQlr+rlpC8aHZOH16OpbBTwgyzEMc/XTm
j5HKwCzZj0G2eTWij5sI1dQHqWWYl1Ndk2Ng9ebZyhtWz40v7xtAygwtz0q1L9st
84yGpn5CtXARtj0ZMHt4b/iob4jahh/Ig3w16U1es4+2zPRw3NEQraloeXq6ITLr
44BQqKOg2cpN6740LjJSc2IqNFw0XQ868sKOSV06UI14G/j7fbYnGgomQnS73a6c
L0DTac5NLwnxn6vz7S9JFnFSmdb8z4VZm/dy6ON4dw2Dlx2wAKhXyK8z0MJsXtvU
OsimxIJ/sON/yjk1Bpn1ZPbNygX/rnVltSyYoBSBpr5JafumwNHpoLlzgpXs/6O6
/LNf3Tx9aNsrGzGT3QIpbHRMfJT7cCFndKKvzXoOV2NSxuEJ5gOQmnomnr2zXxXd
0ic+WjsYdAiEDl00wDkMKCQdq7pjkAqktNfFVAXxu20dyrKQ6Cnv5UYMTenUSPpN
2nQANFHExJGFd7xPd/zPw5YS4lxoBZAsroNiUar53WgIXIK0xhUlTl9xM11Cl5Lg
V3J3Q04vNzxmrrJ6RuaAPmM8KgMBuh991SYrKnIAYyyoP4Ykz3YpUm8Qqw/x33at
Nmvw//SnXmg1hW0zUzGew+9UIHLBvQypy15ENmvjflE2g+0ChKnx3Ib28O6PdLnL
qHTq94xCGLkYOJY0XLRXnp3u0hsBhhUB2i5NCFIVM/0XsU9NZ/UubhDAF+S+0vEB
5rzpVS4zSpJf8z6K3JLdd1D41HBkEdLPQMnxx/pyUBdTZIQRDlt8TeMXB5EaVogx
f08GmZupGK32uBKn3szIt5JJNIGfKocOCrpct/3kZLwZJwzr25LmPjB7nSPJQzMY
f2FKkoi6+U+QAaQ96objjuloRMxzpb5AJExBLCMrQzuIARX4/IAcf+loBLTbsLTz
Oo2YFIsyYwVWDV1i8RWuWw719YGFX29efheLitgU095IGb9pjjyjZ40aRCKVSpR6
R/Qsy7gLaaU1a2BEoIM6iNL9ZfTTfqqVAsNSfQ4w6WWSrCUtjhgRB5hLMV2AGS/a
doyH+crapiGvgiwJTkJPu982GV0sVE36dNvxlXefXmTKGXM9YpzHTjybA8+3KljZ
PO7rgPbV6xpOfoailEV3H8Vft1RMI787+MICC+qbRFQDd+dcrdHRsTY1EvtC3Fi8
yoFd+3plhopd7hpQ8dRu+qON2oqlWBMsJApL3LsIygCV6/1lPYroyVGQyDXh4LsR
715CkapXlxR93FFE6D5uTojCvAZ3ItzQ54FR/mKE3KXsPVVX5oQO+qy4a1qLjw4a
Dur0MvUnd68Gde7XdcQwinUK2ClG+GieQc30WbrV8MEsWMyMzLXRWXoINgvscYZO
g/fLnqcHMFoO5bW5ewl3sdfHTeR5XbutViEgVUiVxz3gmgfFZ8o/y8feFWnr1d1r
mNTWg4NL7RTyfYEjam1QgU0rFgpLoMsq6LfP1PEmcO8cMI3l3geJ4Ih5ZuNi9VDi
0Mg/6y9mRjsET+Tx290kCXcnI0wFvEdSpW71bikwJg3s3LhH7O/Uqf62+97G1pur
Wi26s+oHLQpktGnZVRvMkvM4Epqo1ItK/7WK0auFMSQVnBQueF0LnNCp/pNAjckW
HychZ0tILy7CGKALatzkdK1JYpFBZnvCjRcEGL14cJ2H/oAD7/2hZtDwAQp4QxrD
ec0NzgdCsZ14EMEhu0ugLTAG3N+H7yL6lQIHHZqG7kvrBLbFwZgrxCFYFVQpaIeC
1ZQIdqFipEL6iWeetdeBgecS4jiks/wMzc+vKgaLF6Jh7iiM9OPE6ONqAxXnVC5e
aXFcGGkSzINZ5piMhBf5M9VDMTrttZ7GGkawink7/8TXu0mk7iNjxtXEgtTZ+7Zt
TxevcJxsJNRSxIJbJfhZWbNkCTwont4ftsnTZUzUtxIPp55qumfZ62t/s9HN20wB
VU42yb1feO5qyfi7CttYZfWkryCZxiAturleoXKzcLDKWbB/o9jQpfyzaO9f0uCW
6KBYdNLJwzjyBJM3vE3tC4l/XKoQa1VvbmoTtfgGvEE3t2KXo46PQc0raTSs/3Cu
LJRRmJD8c5BsHLSJ84GlTWVn5X3F5kB8SDyMkI/FYJP5XtIXw0SfEPZsFRhh0ja4
pAVbEB002wnLL4wnCTMlWkr19bjV+jZXSFwye9XE7eiEuwIXsyRbOblFW/RZ0jhO
IEt08UYJBI8KY62wYBVHtyEnVygU+eTTv+MGHNoVUEWQYL6OudPQrfDj6+6lVvm3
DsW0epq4q5NlHzXaObm9xPqpwln6IHizufg9g1OvUFtMBjuFR8WhkXfslBiIQCRD
Lo8QA7fqNLA/hsbuNbfQ29UDx00k8BXM+IccQRS/b3yuOe5hQgpTG3mf8hLvJ/eV
WI9JZjaKsfcOMsYkEbXddPITuFw4SDhIB0lCPecuuQH+ySkgha1p30MORltxoLth
WGpTcerMgZtD7KU6JMaboJho43D77u8OixC1iBd1LffC49DHqif1o3NWKr9UvdhW
HWQZlBLN8pao+tUETjW51ae0MZ+fhoH8UkJMoHwPgIPmaYCITCfTByIRKgi+TvyZ
mC0SiebAXmZ6fZ732cS/LvIzEXOZnckGm2u1DshYAVQm71HcEABoE4RuXDtjf6Ct
NkHFar0CN8dCutcjDVOo9obZ4UDp6OXAto0WNM84QUhhnAYDec+rSZqKYU4ku/ZR
o+Poaui+CpNUtqFy6K8FQ7q2w0zzPj75S5lnBmOIc6CygE4ErB1/ZdTsnxF7oVc8
VLc3ffpMqkqP8reHCo5JOvR0Rmn/AcvZmDi/cou8J56tbs9X4Dl32v3YUnyLzPx6
1D29byPVQ+jtglRTHt2Zi4klszOc2VytbYWjT2uKVJcvvwZwohEJ+8wgd/0f3Ubg
Y2LQPqITXEOik3qAb9QhqblWg56AhpNtDvejlvj+8DaTrVS9cWzRllWSnpbZqa/B
Y2UplFFTwV8i5HJmvmrSfJzsgEQ8g/CPHe8wi4SmaSzzfIKo3SceGHECzBPQeYCS
KFq+uq6GErNSFFy1LAx+xImrAxZ70F7MyuyoXz+e9NprFkMbfkZ+5gfwCBVkvJmb
vav0UyVlEU8nqqUUemzKrLDCjiy2Ws33NhpPjgyk9Ung9IR638J4ULh5cDiRlv1X
97IkiI0eA04YPq5U87s3RDrbO5C8Z418WKcQMabUIsET20cFnDkfOOCIljRuYspq
AaIT54n2xya6ILjrm49WuyqZIFVpYMjt8uOzNDPEiNBPNuxjuI33LbIjmW8CxNyv
I/hGUIqCbtGrybZSZpRo1DcZ/LIZ2ki5Vo9ejReAMubGyN1/V5p+I8hPCfvnGBs7
wFk6627qFijMsOGi/S5fAvn09llayEzMet14fyHopM0VQ00a+RTC26u36WZGlUoR
uQ1HqwCGiKysQ7+1gOcPAZRWhQiACJpTA4U1PUpuyG4akydGI1G9GA74TJS8EH/K
HG3wv/E24jT4MZPiZNVWO04rTItOFle0cU9zMy4k6xSvKeEZktk1DlZyJu97O+Up
MuwRpBZG/zVBvGW00xIS+C9Ubt5f8cSpzRaQLvMiLDsFwZJCW0Oj0ORLUs1LkyB2
vYljTjdo7RywrJXRP0PJ1sPLoJDz97IyfixT3NEqDJQM9sNSBm49v49wM3ySRy/4
80igRzQSmk6tFarT6K76yVQzH9CFheWNkS19cW1p9MwJFbXlNtyrSuhL0+33KmTh
5HTwIlbhXE7eZ55wdkKESRnph6vkvaBKEKtfSLvJrnXMoAUPMD9aB6/sOApYT+I1
QqsljXaitN8oM3n6/FMQpjb+vi4EK6CGEuSToju5XDDxUFoenVbSX4TJQkYIXm9+
sVQIweUin8KPyGvwhTRzOi4AN25TRKqQRWdseSKkG05iXkKEEQwuAe+Q+wzOtOMT
0rki8oIM+ls189UMSuXwFQ3NeDtFlqw4l1hrz2FlLiFQGKZm+CbKEeItYD2vC9oQ
ZVjUjN1nISygCDGvhdxvedrRA7KhC/EQZmlRfrlvt8NkpN9rgN2/arvFnsMcodkS
fnKZQXaA2AN95NJHTJb6HHXJ2WqwcrlCyW7J6CSrDHKz2g72JBQOVqEN6H32D/gx
YLkDHqkPTmKI08Ug0hNLs5n+EFbfBDN7j7b1DYTD7wvt0AJS6EYTpXvVqAQ3s+0+
JZP/nSt59L4n3vEKn0fTwxF7kNORUyeB6GyChsOV7j4+6adj2YmSfoPuaq+zupps
MZLGOa/3GqH6+CO9ca7myS2kXMQA2q+Tvl0lu3Rb4VEP7kKMeoejAoH56PIbUbt5
HE7NK88SXFI6B2DpIorC6ckrNmEbZaV9iiXt9u8o+q9XCw8yMpRa4AbtbwtOD3LH
USkxY92rMEDe8BcZHGSfQtxJMaNOqGhaLKQRzfDg0AbArHhJ4RGDWpB1rMTOZkj+
dYHeGIWge+q1wrckmZ6q4bhVng9v0P3mLNvmDla1K4jg30of46XL+vaGoCc+9BZ0
UNksKbmEd2CWQpGJ0KrRB4BSnLuTkrBiH+WK3IScvXJhy3VeHCrYpoYFuvinF8VD
D7MLwc/dwvhl60tacsDRGAhVCkTHUax5GMo+OaPlCCaKXbRv4Cos+B08WI884w6u
IeF0fgCwNiQfuzubaiU1c8QFp9ShcTJpU33k9k2WNpmUplyGU63hLVYlQdSk8HbN
Qs4J8Xb37rfLTA6uNoE03sQjUCKvioC636TXqOCTCxptwkYKLMJwbO2zOyO1vcy8
fw3vu6yZq1c5/9w6WqDaxdvcSeHWubTv+CPt4m6QjhT85xP6kKKH6+MaHHY3yWth
edkbcGq2r7RFJcUEUyhMygQ44L3F+tfnd5VjthUna4fxmL0ck9TPPVXrHYrtgVKI
IePNCBjHJZIJDcsEYQ5mtbBJ+ABqQ4iRWpPl2UW2a0GtmtBcxRfHw2a+25kVajhi
yHre/hNirsFB7iDw7daI7nS67i+Ikxgj5Sx93z7yOxz+WIPoZk9QQ4pUcoYD8Ubr
rF+WOLgWym36bnwUZMaf/2lDaoeSi3+wQ3M2w3xJr1iArJs1sFWvWATFxz/hG7br
wtHbQ83wLjZnVi1t9f+VRkQk0rHmVA9QKrllY4YZwDWklh4xZLeqBat3EcDvElYb
sQrUYuLhIvpHj6P51hkgwnuF1BDUXvIl4++VpiULDOYfxzbOEnKnzpEZWlylyH7I
5KES6P+Op3aJuWZtRpxJG4MZYOV5oqmQXArfKJaJPqn8s+4XW5NSNHZzwYt93C6E
mLyS6hqeGxHKi9dH7cxVYadG1qOxrlpcH5JQCp+WBCLiN2BYZUw9Dw7//R78KgKn
uSBKjH+sb+sQ+9TgyZ9YSdQcyXvlsvzoZt9sigKOhjVm+vzS2UzKjdiSoQKlZdKC
XkyLSAt2vbailgHlhW9sXq33imtYvn0EH2KlRjpmHhaCUndJfTVig4heNSTq5l0A
beKiPdGRJMZ+4l19QxOg4BFE6LxdwgbwmZO7VK+d/TSDnyIDcI5JYMdzh1/jL2mW
BuiCCbYvj5LvIuhdyrqb9vOp2YFPLfD4OlH8MYTeLWsSVMHAwJ7g89x+CYceCxRY
WDfPsD0nUvizsKb5IO7MvdF7F78wTXfYy4v0fghsEcTedkIEKUFrBxPDvpdydv2n
SwPlXUJkEqeGL9DOOpvuj86dr3BRFV8M6af7GlOCGX9DXPzgy3lU0ZVGhOCZKyyE
Pjrr/xowuqSNEhu3gHE1jJAyigGRyewaxwUsk/Kr5munrDTWfUY30Hdejs7smkqT
/gUXEGiC9E+v1xwQ0OulZtMSXA1IPt1qoYQN3tI+IS1peRUt/VPc3XpLs6ZnvwHV
9KXQhvAv4rQf20o72R6fr1IhVumYCQlFawakXazwabzrgDgeURSvc42tC5bqleKG
y1GQWkwOmbRgXDqSA+e1aR1Aa90yExiJnN902OcMV3vsDZqbc2KYUNZ+WPP2kz7Z
cZLSxjG2jSamdh31K3XKFTWQipYozSqGz/H1MewATvP1t3ZFRlV0l3j0cyVvMzD6
VC2+lCurzwOcRL4aEYqlXZCI5Kt63FAGuiR0kx2IwjMksmD5Jzm8dTb+MLde1Oz3
ss2Gk3xfXFZaNcBT1Fmkn7qyTj+KFEKVVcAPNeZM/nmAigHJ19WzaAFvQZ12PbDA
KIAy/xhDcO7dz2OAVb6X5WNdtY4I4Ge8bT0CiqvMk9qE2G5JkGFjUM/2F+mpJ1FB
YCDO4HGkrJ5WywRnTmDOAo2Tpzgam2m4M/AGcyBmNmbjQcDgdhvsE5hB64ItNJ8G
gGf6CfwF90OU88x4tW89tu7I+j/PGOme6v8IBhRTfYtEYZKHk8XfiAxJ9ocZQ4XQ
4EjNl5534KCxjuWPfmjRdvOJbmgclnlmYrFItqUPadPZb3F1Ras4ha3jUoAHliiw
QiYD713GuOyf021uBusKNjDne+Z592KbyahW2qdkJxAvxBya9ESIBlA6sL0UP4AR
8y+gM0m0B27x+gzTKJojJ2Y3ipieh9eSMH6ix8CnZEoKdo5CDFdnsBNYFx7DwffK
sptVd7w+3eEup9mrx7l9pAw88WCWU/VFrHi8OWD9bOOQiTO2S1Bo5dEo+0/ojFyW
NpzXO3CT/zYYF++MsAvIHQgmKxKbvyWRCNbaFpxpJvBXbYHKD0SVX0tVcpumf/J8
QrYOYHf9XXgwTnFx7fVov7yf4dwWs9coxCLTDuwlYmKM0HggqPxRujji5lv4A/Kp
ozm//ZfW4kIqcYzwp9rgYfSZGvYss5QbRslwbcp7F3dXSG47GY1fC5UXdzOOwf/n
zQUDXjiGCkg3qliSIpCacLmX86nlYBWGGZgLh6glYeBTw+9QdjcJiCHcJLf6Fvdn
YztSIgHzyEcIEUBJFBD2PAvzwLOLm5rP6KnnbipQbbM+OgfvALGIHuzSWZQOI5Lw
x5hkYn5EnxT3IFOIVwH7T/YjJiR4bLGIA1IzPekfCN3ieGhoEfWAaMNUMOq3GNEP
cFpOj6/GTjoIu7x9hAx1DMur0SaPrGOg7hQN+lWhXKNJEiodm8Edex3YRMGFAwXK
llWLOldloyyD7MarowUV7STMwQGbcMR4vBDsXSrWtzo8m/T21QsvWCD4HoDz6vxN
oH2yHEZi6FilP68bcSDBG8PAkbq+yG1f2g+MMgP9pNnHpG4dMFKRRAEFt0gzUI2h
Czf/h2wzcj3jXNHmFOi8gypjT+5bK5yX+bCg58IUa4L8qW2mUnFcxneoqO6Bj6c0
lXGPjyFQGoVydwAXAHQ6k5+iQbwtU9j2HBb4o6XaVrcNTYvN7suTc4ArUwGyrsET
NE49B0/MRHrxq2SjLv0GDDc0nTK1UqxlovQuFQx0okJEMC9m/muQilWaDgMT8sa6
SxXzqFzyCO4CSQ0UbDochb4Ea1f1DzXtR44zGjP6tDZu8fGZQAWpt85Nr1HAkswy
dwDgBIWm+4ze/qSc3VCKbxS0+Dd/culyBdem/6/BwqGdLd60vU8iJAfsDeZ62GF4
8KS14V7yOWH8dyRMp+0VKAH2DSl5xu6x4gMqkTwVzXXLUjJHJWcycPo/l9PUce32
5NRksKN0eA06vr7AwvMipUM8wW2CQ0jBgFvSfAsegUx6d8VBGII3G0sCugXEAQGp
I0zfI6YVRAlwSZZioZAWL18Om50pzzCBm1ro93d/K2ILIwvRf9GhNFpVBl9aypmX
64rQfiWJwm8EIWdZPh4YOzHPYFBKTWaf0ZusSHdJGrCb9UeaA/9ZsTTlYGQgZGoY
OSIUURHEC4F7htYxpKtnJoFlMB1yf+DQ52YOvhb3oRiIn4beOi7emIPbB3vSBbhh
IApNVhS9jddkbaKt8MjCxR2OVcPEcKoO84HkuLiwr59lON4XVqmC2sARlR3C66Tv
l1aS3p/lP79nD43YHX64MuAcRc2akV0RFumpUGW3BP3qyZvr4u04nmN20ouHZcOl
xhM0qcQZr/ettxLVLYNIWbdagJaSwlUDAFYMcp/aa9iZLzTE04nDO6l/2+nwbmoL
4s+qGNRTWkTS33zxg+//WjJU5YcSI30wQtt4qp6eHWzomjb4Ieq/onH9AliOXDhP
Fd5bNYATIuRaQLC34aBXMMdYApa+bR8MIcy23wNdAQ4NEzNGIxQSbKGkGjSsRWb2
gt6VkWGCj49itav+6szEh1FQFYbbdLGjbggMs602jKsJuPw2nk/ijxy5rMODK3YO
cEJMkeGvQmZbuFXc0iOibNxq7M2cOAehdxVeRXN2EmwI8FG/5oYPcMOaY9lygEqZ
ROz6SgwEX1LO1u5KkYCm+vgUBArghXnBGIaOMHw0kgjjEKSG81K3vX0qpn8D3k8D
AraC/hKa8vgYKPulkKGBaNsi3A+dvQQiQBKAfww+S6uyP7ccs0OMmpFlbAfb+lL4
gK3eK6dC0EJqZ1bSj+bWi93qkdYeC7+RSe8eFaY5Jde0jZXy7F7HstPxio7RV1Nl
T5YlpneeYUbfJnCagdAXcHiTH+RqoAWgc+8BtlfIDIoiTuaQN8snMz1X66gLOqtn
uo2tDdsMPSBPkAfAqTwxQtCfM0GOLdUXePp3b9EooxlKn8pcmSmS6cM9di+7/XtG
WODEymGFWaxipRMlAEex14R1ChtbP56HNk4/+m/XwAjEhB6KUjw92vmEABg6Q+hw
+LYVLtwvxlzW27eWFItA2GaoMWeN5i0fr109s2JQn6G8O/dQnwg/5IPRQGqDRedf
Rf4ugNQI6rTDf6WzTzE4+cr2w54gn3W5hVPqeRxHIbTJb1nfUCWVMTiTKjGb8qJZ
XTTQZ8QNOYUMgl7WuSnU/LH+kysLvjhP46LsfwydJj5wTVGwxAm42+7xrYUB8m91
8bFbyNt1hNoimfMlJzaZhP2/dCwxXnSEoPfHCAxHX5dROpJQ4PzNPbEh85U43+nr
r/miNiTOt+RlSZa0l/Xkrdm4mJbmdZ3JBHOxaqocl+0I0Zv1UDpB1ca/uz7OThJZ
sI3UUGpO8PVaUuKVqfz8jo0GBoNXSO6RRFpvHmfOIAMLOPM9a/rRj8jzO0o1Dxcq
pKyu5qa2TI2TKADBnudZNaffdCQLZJfRYEjXd1UdJ/qjI5GYNk9iqBDUpewdo/SD
SvKThpwFQ+nSvbuhlmjSHaQ44wrutaryiRIncsAE5MIKFm5W7SolP7nxCK7ieJzE
LI8s9V7C6HZDWhwgw/Jzk0O4FMIDdQu4zEFhYBDd2SI2ebOW/VMC2ikVmeOOoYK+
VZXf121lEKlN/lppVFbobJwRTAy5eBLz2lXZBzlYJh65pS/Y36/gw+43Kb0f9gyS
plC6+famvoKS9BMikS0XZYOoKXDyANYNtctiLleXyYZ2uqluaAQ1L5mjWJouDs4y
gyQqoVAt6oWzk88MlkOLjO+ylizBZVWRCWThOiy72+zFL09Uw8rVojFDMxjefdQ6
avE24DwGWivimOqajdSHlAF2eIbBm2xUdmSYxzdZyF6f3kmioyPl8lA1tCsrso+5
wsYkB6bpp4fQP+YmN/yfv/WJF9iPMLNkCFZ27zyMrFcg6JST+Au2cW+kAFjghgiY
MToiDPzDaEGyUzZQq959ZyDB7Cd0RVOfAmQ1debMUL/cLrS6rfCwfTlZTFsdcAjH
9yAfSOFreS7XsdndQl1YMTtcsHZQu5qJv8+cllLOYQqJIAFAPKd8ixsJFA3ylotE
hNF0I7fbTw985rqnbrungs4x4GbM3uCEw+E/dTAJhhn6HST6UaRJFADVYmEk+V3X
umGeQdgkN8Z7dIiXtqR4L+CEV7D8xeWDAWztxj3ZUQRoP52QndfgE41RV1S3gaEw
1pR6rB4FuPkvkMu2PI8d99VxZt5OwT4Hi/pg9XgMwuiEpi7uS2qHwZ1ZFtChzzm9
Hqrsr+1u/U3+N8oAoKbONXxW+byQAVRFB8VWBtMIoRrUHlcj+IQ1SPd5yIopXHfa
Zi2Thp1kL+c5rJvwM0a0NrbIk+4ET5mfzSVB4fmvgjpMPWVWvBBMdw6tpJie45ea
/HR2z/lVI+zbQrF0w9KSMbVT9EQIygf4PO91YGTrNvEx280UIZZEe/0n6Kv/iU4h
yTXB/V2SvhzZmz674BR3iQyCUB4D4cURrzlLzEXZ31LxSBEMef6bRW1lmgOS/HnF
xeAqMEEU94RGoD1JbQWht3kPorAnqDl5gq7T44/3rTUl8eBvC/fjaLL28LrofWkp
4cxQZXffIi1yVa3jm5jEdFJ2SEmNs5W+HfUs0WDuMnAW9Pv2IfDq5zse/4hViYpg
yTa3zgtsfpyJ85R/5r/ztI4rrq9D+kE9AMRBW0CfXzzC9ptKrcVN6+EfI74HZgNu
c8mfRt0ckFod/ITxPCLCjZBkGlu0S0M01DenpZM42G0K2H8gezllYtKAsUrAyug0
atDW+U5YYPqyRO4oVE263aJqZ83TIO0evNXDs+f0RCxlwlL1Zl2NKrsNsRJjeMk9
xoUKHNl5C8uujIap9gHZKVp45mlYB424sf3F4mKxxHOocSa8L+lMo547qjG7QjEK
TDyHnhQkK1u3f/S98ZOog7RX80PznlhvK3fr9+nGEkBZwSluYOnGbP+UBq9d+Jli
hSzbH6mugMuV70ZpGN4eyBZYGkRefJGmVpoHXt33dnf258UTkMeJCoLxTZIy1roJ
hfBfvQ+Yj/Gq8eBx/obrqn14RQ7S6ALIVpFw0ZQPzXO5G+7nowJA/M1KXPTW3Xmh
de2ObioIKIeD8EvODFuj5ons2aO4da4oamotS5qWCVqb9O1P75ggBlhp7w2B5R6l
7js4jIXdsPvKvOxOc+NVEEuywA2nLrMPf7pAp73Yw/4PSxO+1UnNkLcoINNlZAYN
8u6xq4e1r9/ackSZvWWE8/KniKblmcDS+i2qdZqI13iKfZOH/rXVMt8lZUpywX7i
7WZM4cdm6eACPu468NMww2oT5vHmvBIB3KPpdjKZcCuOyFW+be7ir5IDybFxdvjW
pI7O5cwhDu5/M+C3zCfs/JVCUZDRISCbko5SNSVceC53bL8iIEGN9b6iH4BcOShJ
GOAyJcS+Ca4e4PpIKq100fjk4TVtlqpjA0hIYVg4vhW2KLK0KwQguR4vFBPloVIH
tb/Cw1K7F9gwYDCOuQchLpl+8f3G9Q1Mj0hmzKMt8Ev/gJLgz/0EAbcyHnkDwa+b
y6cVMIVwXdX2XJvS7HeoMhhRWrr/GQg0PUeTmke8DVdZ92buDyR1sVBCIB2fRtdI
1FlUFIWxiP0eTzms9KedAiKGI0bOiPJNAQrjYaBeOTP7aiyE7lAH/IkRYekyvykj
FNTbYxNuQ3MvSulqphLggAHA4NHuyaEk4irc/zgSleVH70e/SjwWVXDxv0kJYANO
iPFydYs3IWjQzV+j0qCJ9cDEmh+1SKUdSi469PcoFad412HCAYPuJvMoNS1gtMop
coIiXGFmvSHsSEmbQto64CIVndZgTIy85VgFb12VJ2b5MaTCKnMFich1IPq84EvQ
JTTgkTsZVBhHl0LoZXPu2vEIx2LNBWJY34DNG/7gK2VbHKRR7+FYhVDQGfmx3s9U
gSEI+9Wr9hFKyq8YISdiZcG0HGYYu3iYz8WjPPbuF4AIPfA+sT9EUd/ZW9LyK/lq
4oLMSTQXHKR/70hVXdaX9UogBdoM2lEv5KW7ROpyKteWLCuZkO/V84BeER0n4dBk
recvZuTy6bsbHJMtP4BjOing0M7cG4WcULnOGqxQghevZfjyyJHW8ASLCk+WXsz3
RD9o/Fho+aOdCW9T/I3dMxxm6fXZWP/SCVOthmQUql7vsyHAnbJJG9/UvbwI3LOh
wj4lzeMUALuVGCYgrq5dryq02QdAlXpUiELo8jWAO3ZZnAO6c5/z3/1U5B7MGxdm
UMQ6ZT4Uzj4KvyvfVAlv9LffnS03o2xMLWpIUqroup08oaugwpNHEdWVkW0Gyett
wLpXJoqHXHGOpaujlpBObX2GkJLdr/zob/vTnFk8l+lQfU2j+scUeBytsKtlMU8G
SUmZimE6r9hh4rOCbqsBPAnxowwp0sf51joCX8E6YYhgXY6VwGhbPP//0O0QzzRp
wXTKXB9gtuPj1XKaNcqvTm8T8ZP64623cy11OMf9XWV260bh1ulDh71Dt3/YRMPN
hL1c71oTd8sBXTIjbuxNLo4+bgg52AZ1JqXV1VxA6F8yBS6KPtoVRLBnaQaIPYgh
Rezl++Jgb/4fC/3yICFeXChYQiVxPbCAVsiveJHUTvGIDsccoRUH3IGbPvkU4710
XWhEO2BXfHbLJwO3jKkOyG5m5DmOz7m1W33hPxCLuVIGCXQZHPn5VdmvvOUp8Q0Y
YZJC8x0AgbI0QJPLHmX/7RZk/GRCgfgLqVeuSTLruhGvllbAAQeTfc/MObKAvVoj
GeYXCM8N6BsY7Ugk6lvUB2ekLMfV+mE82qwdxDxN8xFcuHvh4x4y/YO1v87OxxVk
yCa/JM022WDRIUzy1s1Qb4mhGGOpiWqHykzA8T/JwtGY33BV1XfOcaZenqz1eHAD
aZEhF+r3ItXO9PN2voKkyY5xhdhB7PkkHpqDz3H6ay3qx3xx8N4BEgLSp6at3v7Z
lVkJjiMVJf456ACc7ymVNMUShkkTo4jQSL+IzbI8P6MalOd8F5DOjTOXbSC/Rjwe
PSY3TRFcsdBXOx4+2faIS2FRiEFGmB4GYzlptNqdJM/Nets4xpe27D/1/2+11VuF
XCFmBEBhy3+6HSpGsHoSj6SKk/rRE9IxMlh+A6sUHqd+HGIa6FIXo548zywEhRfR
8BLPCghvc36iH8M1B7fW18FQbQ0awWBQ8p1fzuOiouLIoxpaqS8sGa5eWLoRUhz7
Z7gYBqV+PIFy+tMiqSJ79oT3OBd/BfeKRgXcYdSUZiJfzSOeKZcsHWnKOQkIic03
lcFCwUen+MhCvDc20g8XMzDhW2s1JZj1su9G6/vJmtfKEX7R6TItLQrHsU24wz61
5HIKfkPr4orA+cZqf+i4jMDfjLzrUKgKPNIZ/Vz5T1YqstKd+TNitwuVXT5gt9Fl
AqcM5df14FTFWOqwdVMaFOVozQDic4IBDYCX0eduAW3EpPkOKtctJ9MRRKBUGLYi
098OEfqrH86vQf1rZTo6HV6csD2BoVW4FV4I8/ylBOFM8TgBNErz+gHACycv57r7
pGC03YdHS2OHOrIG5sg/nu7xcUB09xlwir9UErC2TTzu98vCFXM2zBP/Sg0iGN59
q/6ySMnlATprIGrzYOd3VbUa4v2QbkQwjb6Ar9RoQa7i0HQQo1FGNQoE9v6xSzzO
hckoiRMRahuDd3Qebgqm938fW0x+NmnhKEja0g+OYGacyA738dvddfDuZOgN2fpX
oPWi1/nTh5vRPsghoa3Y9IySitpBUJZtWRGHYl2XK7lN+/gJj2D9yUvdHbsHZ+gD
zsN0oeUHmx6yDqisadyomyS5N3rWoJzvmMO3LMS9Pre+L5IRcfuAilGgGQqGfwPc
QoqgPkvNwKQ1SQhJrcOqe9btv1Y7INknYlsEVFe9s+sA6ZNTPG9DmTCcQa01i/U5
oXk9cYG3olx/97+/A88XrafrsbwJBHlOOMxCNcXEW0t2nKRCqKS7rv7vL+vCDhst
/DhSHQG2GwaE6ELQfnI+X/8JgkWnKnF2h9IbXFSX3mG0STMcqHvwXnwvNAVBJcgS
lR9RMd8NWkcKcpnqCDrf9OWBEIeW55JlvW6kIda9I3Qp+SsTiW6E2die/ieEga7k
kljmeZz/h+M5D6Ai8xV9BAxi5n9ZNhoHsPveoXs1+35AnVUBpU6URd49LN+QdAXP
lTR6I8iD2nTA7hGz2p3Fv9VsHu3WGL5YChTobyVLtc3sqbsdD51xdfLeSrI3sXJE
0Mx5T0at2WPk0usKNo7VYH5PBmmbV6Wpmq/QRcrfGaJUvg6xFueHBfm9HJGKtN02
H7EyHu4XEyfwB6InDFc0Efqc12fl5vNsscThxg1SsUchh6mRM3WTnl+IwCof0HlO
LxbEUZmdGqlODWtAsow1wY6hDWikEvsdDWrD9GKM3jEXPdOAgxgimlpHtcfdoF0u
b1plVKrYU0gTtdSkBXFlS7JHXUrtLor9/fiTl//Bqrpof+tTShqXCR7yYEhHCCCo
RKkkO83IX26bhVnoxzYi4I25ZgZuvjI8mfm5fqbJBngKh6b085JBYtnNtqcAlkJk
fq+DQLb7DpmOfJwjGLeTG5ScqH/gIzDDQy6Tw7A3urW5ySwkQIRZXALQCM/UVzIc
0X9ZnvvtqJgH1KfUR8lPTV+dzGaqQvcn/BfeGvtE6o3J2aBJxO9rqT664+IoGUfm
4DBlMjhJtoHZttovUy8fQczUDi9PNAk5OKTnf720fg/r2pOByO0emZac1vdsuPPB
JIDsh8c3Hxqe0UE0e5nNRXqebQw7x/apGMOCSihdw5jkPXUeRP44+2Q3sSAX1/eb
d27/h19hSmpkCSJ9iQnA3zLKMFA/6oIY378vxGaKl5RQN1MvKYXExL2UKnXrSM6r
k0XwYPGws1FTOXb1A/k1R39u/czRijdXUyqIExvRYyH7h6MCIu+p646MdtmVWyTq
bgTvqOGmDBBbYiKpO6YeO4MgO/+kL/MKDjjzxd6qpLoyYbzMWCWX/11Mvx5oGJLc
ISIwDxxI1yXooa/ME2IWUuUUyCPgzDGBjc6/iumpwG/tv0BPG1goCNeYPNWHL9qe
rR5XbgzQKtj9qhT+oIluxKfI1KbBAdabPKcWigRHcaVM234GQduc9lXijU/lO/14
t6jnigXlLgwbUtlr6ih2P8gsLsedx8lHD8of81xN/428U10AkdePMD+i3a5OVRvl
NE8S3rC8K8OVmg7GgTl7aPUcDhfC3pG3o1KTnw12gNqnqI6SuO+Y2t3RvTQWGaGZ
vL/YU6xCDY5kEX8Ib9clx/ocQ2bfXI/BwIKZ4F2wIIEEn92vlj1hH4HnHa26mZIp
wLNoYegABYVGCtL7QkcJ5+YFdpX2dlNaYz5Jv3PDgNzoCr1Jlgl0WP2auYx6q7cL
RTEqoY58H9Z25RrSuER/1bcmBbd0RX5IWbn97oPvyl6tz7ppk6Rlj8HKLXqgKSBF
LoiV6x1f3QGtB0nzEKNMLfkCj3lylbYzP5RerPgRHh9CQavJi5EsKfXJiQeCclBX
zF3rUwVJdUMUAUxHkEMck4GskvTbiZzCVVXJaZwC60nvjW8tf4CBYGKdiE1nowDh
DT1GQQLs9RAk9/LJP7Rq1MCgrBHe37J5qsZSQnJVYjslP+/2DNbfHRnvh9Su2oL0
YXkB8Jv0tgpH5jjUWipU0gPajfhgh1msD7cdR9tyY5ahjX9sKX7WPyY979nX6jT7
m8DgPRpmeSr4+BlJOxgXgqq2zNBr2QHxdHqYmTVZ1tvcBXf3E8YHt3TJSUEN4Ewr
CnwpDomORDkaioBgghNQHDL6CzLF/jFaUMOIyFWACzeJvCOPvuqckaHGaL2rmYpo
z7VN1OWLPxnFuFkISJ6hmBJ0hXhKg21mED+3RVPgaiinXckYms6cJFi8g9FmWdk8
jff2qJ488E/94u8TXfCgmcA4kWltm2KP5bL1w712EoJNTt0DdoGa1j2ZvexarDMA
r8bV6m4ayIYKy9ZHb5NlplkRGnq5MNL4lIjVH+tYeFW59ZgCVyEYf1tj8NWes5Bf
tHYSSGHVq3kdevEfkk87ofPVcSdvyC3XQRnMaDUe3FyLpx/P1hNkWR9rpkAQms3n
UZqh0fpTvBtwz7l4OJNQi/Ud69wauiW5c7G+VmdbyWOcrcl5r3ouGee9D2KL/EED
9EKKsBFX043ZNtpTMIcQf3vaecmQCByhQTqxRzSpUqzOb6kySsyyQBOhJ9S50bmq
y9xI8xylZzDV+OeL708GultQbCOSb5cZsHE13T6Af6ldUTwqdJJQCeAkahzkGfPV
iMBa4iX86fk1QjdJmxD58ginM11839xRl+Rjf/S0mHCuRWf3meLTXPBrmmrwuotE
OLEFns8//jfcN9CY9ZHsYa2xo1SCLJeorEk7dV8Fkuwi8XzF5+A1ZFH8RB+jUXSu
VrOORquoq21Y1GUb5P8Z+eIwqoq3Cq9w21GPgwEX9yRxmoRJbwsFdG70I9UMu+Lf
2rhWCe/9ic6nAT8dqvoG1ql0cL4GoQsNS2Bm/kxIOYvaUdYIYfooPW3ws2B6pW7i
7pDhqEg1aFwB9D51WH/lB9oH5wBMBapjhFyUdV3GevHXXWNEwISgo7HCvzheqXak
hm76IHg7iHIxWIpH4Bw0KCrATsUQoXSK5g4NzZm1aUjEuEO2b0LpAJ65Umjychmy
KPScNZQpZEJgolN3l+2L7eLQUqjoPZkl021wik/x1NmC0WudownmXfQwXCVl0xlb
ZKtgkRWnN5O8auVEaiHJi9aXH+wudVaCHCHpway/oKXIs+IowQ9ni88wKUI1WvfJ
l5bJusHfLkWx3d0I5SqLTaiolpTv7AAl2D/Z5Ww5AFy97mOhM2v+g56AEKWWIlYp
BNzVQRCWf0Yg1IjmUB+C9wBUMfK+bUhCHzAhsezAWQROtpa5mPLsDr0V2OURLuMZ
OqbqtmU8zoeA0O9ECvONwV1WcOKAP1vE/YbryKpWtjZIgxLmnmT9j68QRm25mxKR
wMSd8JQ4WqB9gJ8IK64qU23pjdQyUlBB1ESYBHhtLoKKS/jmDgMeTzoPkEIcK4Ep
5wO7i+m04wwCi5p0ULSt5/xk7cy+LPyjHBHJh6jBFE4ZbG0WxBpMnyedu2SaCdWW
tc2+tqWjesOHKdTgcqLcvJIZOXap07265f3ieNXlUcxLy672mp9xzqnQmFIJXw0V
857x21CoAPdXoGhzSUKMCIpafzKi+gFQd2ObhrZj+TmDua/5bMf4vSg2+qwyNN3+
IV0OswoJz1RlxnHwCbne3x1AQRepqIhZt1Igi94mEwSNThEZD+p+o3k1y/LobPIs
F8Qx7Y5hBLMgCOEKFFADF4UsOUPrFndCGlhZtFi2RLddAxfPnql3goPlMatKbRON
RtE5muj906uvN/JEd1pjd6RW1/T6K9FFi/g/DlHzg3NPgK61UmBjs4A/Vd4Tqwas
fFUP6lnBIKsmAwMBuL18BIazHmMFDWIJ9em7flk5EdB9okz0McsW+AZILapvMSSp
FDjiaoG9k/398Xc3yzExtTIcWCCITrmsbCoF/ZJ507H9NHSQaVnzVinDq2nfeZnW
fBparqHN4fp7ZEcu0Vmxng169UTDRsMTRbOy7ue24FBkdMwlxLkCTVa/OHLP36c/
aF2tc/PvSy1yM3pCZckf1QEOszjNBGGXra/FjyiZHFvt6F6DYSTPZndDf2PZs/vq
BXyB0YmuPgbtM2rXjLyxrRtTuabqc9tVe38tB7+jKWaw3fqXBiXDhiAARoJT20FR
REYhZlrip5x9CDM260sOxpa5HQdxHfpcruhvUdON/+Th5SI2RGGD11PhdbWs+Rh9
U9m+Pyx6vpUmQhcWv68uOKiETtoRf/iZnQrbBtsC77gaCY87dRRzWi4hgeShcLLj
QjqGAkzj6RgoZfrO7pGvK60t1rlD1KHmoLkWmP1t7sh75MKQ/HmCddKHWF5rsq9I
4hAOKtrRBTqJSsgAbezDx5oEQtSGwtvANtvZFSZ/BTSdlQXYMHDPFgcuO3sRTDb+
vVQ7PTBMfmsSpRpxjBAIkUHuLbBTyMRWIsaVgqsYGYZ4fC+ZrE4R7StxU5yp4sF+
quiX0tLMasnNFQE9fnLpKvpQhuJ+qoZYtdjiTYesJvlI97nywRkEB212wNT5NOZ2
ozwV672099RQM5SzigkwXJIU4ekxK00odJC8DEDTVc/7RvSSNkbuog4O00x392FY
HbxuR4xS6cVNHUJ13YU2f0t/ySc0hbe6q3Q64gptdqJv95zNQdpXEzOHpsfNiZPM
KHGQqWzgjb3U8JF+Id1S4l73KMumnqiI7gLvEm5vOffgpuXb6FSxyjr+pKo6jaBh
cOuWmqcLv8oOMculvqSLUSON7zFM0OGSReLKGJyY0himKrO+RIh6KnbiIBrrJK3K
UAeYH7k1EL9DszV+isg7lI89ENiSk5BnxBe2bqLXbJ/uqEjFy20r5e0DAB/zhMgk
waTpfQoUON3QjRfiEwOuNBEbl33VlVTg2N83zrfzn04CEWKBCs8pkFIjWFVLC7Qq
LfzVky7rG74+Fsja6RGSxbTgLra4xJ2twMjqb/h/KVpN63kAbtdKuUZvm+ybsEIK
VNVk75TEVrIYTvy7UZEOE9Cw4jH8cH4YpO7PZj1YcP7RAo4ZPyqLAGv/ucrtIWMK
JO/B756Kz54ZkH1y6HiRPu7El9GmJMnsm37c461jhfqvdaAK8g/irK14HOKBYKsM
ce70mgXQcJK93dVMBu163xPt1cyB5d+iHvpY0HZAtWLacD1ru6pLMAaxxBLej00c
J7iFH42soQzhEdCWcWE17G3kRCOn4wIjhqj+XKkwE8Wp3jzg0v/pSqIUKF7PmZPR
9ijbAAsPUwpD3uLGKKdb16Fb0vJERzmmgaSz5jhgtqEMJbXgGoKWHp6wCwAscpFH
Qw5RecZQEWh9eFawXJSetg1Y4u7dEp7VExbbVbdd7nom+zLU2xEo4bsHvrhcLKsT
TcQ6LJimNNaUqXWa1Jgs2dfyGp/Ba4vD/p/I1NVhzsOWEHHhAICewa7RzLYq83bl
CoqgN7XQxMkFuAUEAGsGQauVTHsKnqSUq//Ccipi61HBNmxKR9dLLBzb+Il1Jb+N
7Z87K4+YWHSOviUfPvcf7isSviK0TrXvnFDr/AlUG7G9A6KfWo3sKPHLY3poveyu
Xa46o7wr9NUfZfY1BjIyw4UU7lRyKrbOYy81ogVfoPpAkIQpJmC6GRoYi1d2Jzs0
ghoWjXgEVWEaXTEBu2W98aPPclrCGnQUOLT/WwUnFGia2AVO98xYU9LkSHhdxioS
zcNz5kRPShldYBcF3D4+M8NfRf7X33uZpCyIMtKNC21W8OsZ+AbeFuumO0E8QSEb
5ErztUhmmLsnmXvTws5FvieGmAbS0U44qa0u68SQYmC2nN90gx8uZXprqFAewB8H
mZZeF2RpfXRP28vvv0jSBvyjEb25v2L7ohwy/V7lHZoimJYsnfN2socrQum6QN0I
f2oXmP5P/wDMoEzib7NpwfWnVeElKDf46uoeTF2P2XmQKOHK/6B/kE47ytpIyQWj
S1SDJA/0ryH+KEFw1AOICevMm0XkOGQIGykCEJegwIXyo5sAm+6OvapV6UqV+Nlr
uJqlELXhnC3iVk0spAJx++c9fc+OP0N66VIvlEIakS+m7xFv9d0Vks2yFvbj4lbb
s8+6vWSEQBtgaBhu9kIwMdo27k72s/LDlmjVuGwYcPaB9BXj02rL0D3PpWfpNfWW
02Dq0f+4QuEx2GcfIklwx20r+zqpwvb0JEa4HfGAA/7sxaRufkTHdo0FT5uKSdad
o6sFXgW+J9nY8n08nYax+hA7ZqnwUNEhNAGAAg//ez6kctMu/anMNaq272X3djyO
NHYdff5oMw2RkfPnyaGUt8q20eSqWd6Apcw0duFP9dJAn2uskvG778qhRRZwRwIH
1i5ACdpLvBCaImwGysEzHvvVhMyo5s+7d5GdcXC7C3w0ZuTx+q6K0JkXu9bbR9/3
syYnJ+989om6Mbvx7pVZVyY642cNY43TYcUNacBCy5JxdhgT5n9w8EpUD7oXqdbF
9Vs8kqN8nshEysUgkXbTE1393OcNmmJjNuclU4qSmx75ZP4q8dYhdBrlvb0LjgIa
2H8dtx6mJENSXRYWyUGsztgpyMChoTV6FnZ4oIqJdRS/SO0Uq7jLdNz+rvchj53O
PcV+shoW2t5pKaSMDJFK//bJd57LOgCp/8Dbv/bXWVswBnf2E3I8wBrbvPCTkDXD
jxu84HvLa41MIHRc2WJg4i96fnUnvzEsjdDrJ2vjtPPg0kP3nomaZ43PtQk87NLp
Mc56m0NuT8vUGwIqopkW7mBtQ1n2HoRuSCfWDWTA2o+4n1w21sghMsIK61nF5aLP
kEdzKz21onwQqdG05MsPUsalD80xDZ8bMjjF9v3/bfZX/SmIW+I56FuTIUndxPut
oqycGtaniT/cEsg1HPC9pNjLxvyVU8pVQjW2Xq1wE+Miu6yBGIcTNpWz2j4BSLNp
/QhZ8NDD/AxuIoK1+pgllNgHO8FYqaLe7nQvT/FsdK65NXmVPU/tWtuh4+/ZKSwb
GN+Bi7zF4+PVGMxVtCw2wd3wB1jf/teoYm8h/e0B232JhIajrhzAUjVfzbybnumh
+HAnARsXxXjDxUE1gKzAZRux6IcBelHqbI/SxAue78uKSjfjSn7efytZfgxptQVi
qAoL7q2tG8AmqRWxPSiWI3uFsLzl8qg6fkN8RsRLq2eGxmgg+yR/nDR/VTEOIEpZ
wmfBDOYiM8Yt5n+ldtz3hDVgbAuGAXA3kDH0Mz+k6JWP8N46JJ2p42WHc7NbUvgH
cVM/gqf3mXOTjlofzCdVGXvWKsS2VN4y5f6c0lyrt43KxXSJH8SDGah1Fp0x7wT5
0zDQjGDX9Hjph1mcYGIJkRwwygz3j+oLVfPSHoDo5mfpV5xvt9/MeT9C5hXJxFF+
XKNaLpoCd+DJwbcXP5AHKvNFk6eiVlPiNk3zUCvrZD4XqMYL9pEk0meme/pac3A6
CHbH+fLaWa+Hvfz/CO7gKRA93LodwqFnWbN7JJX7Lpe3i9OzdIxXT5fKPFYHnv3p
9H+iDQd83C7GOpmhHlkNoZeUBwvHyURph3D20A5PuPV1BvRS2fET49avsrHwij1Y
F7aykDf+Z6sRRfN0DC8iajvAPf/2eOgOLR4VqNcUylg9/uVXX8OaYwqeg0qctdNP
NYMP+aAE7fIfesnanJbAM3McMu5W31e0+OYWe7B+YexOUdGlhrbzav+25c9sSt0t
Hvgj5WaLLoJjYxrn5um+4HYttAS2dSQXNHHv1h97xau17kq8aCqYL8duzAdClcrg
5nXYqQs8QVUYnM7FCvzUHUbmHOE5zSxbYWHAQ8O1cxrHz6gTILvABo9JuKL0nZkr
UWeuNdSfQus5m1LKWNVTcH2GAe9XHAgJ3lPdSurq8fm9gmUgf1xorJiqp63MnlNp
oOFcNJ99HcMScI8E0sFOszV4QILcz99OEsgsKI5G3g21Ob/pseimBQ9Xh9EKW3pu
hSGUuPMsYswZhYow3fhVO3UmM/HYCZ7UY87wwbowacha67O6kJPoFvX75HfwkvIW
+Eoh7zJVCX9fZEE/8T7bA1r4EueQ0SJehCY3KUpF2AAjF0QeoK+yyHMflwdNyuno
BnIOwWblOiF8t0OVpJzQcSGLN6p2Oi7z5BsaqiweJfPK65VOMwJUX7S67rZpUHsc
cmTL8re/pl1OngErlKKtlis3zQ+yIwdo4QAykAThlv0ku39HnUV36jWUpkkeDrv+
K5+/Rk9PeAI3ml5IY7Ll6NCFDR5/pOKD/qgD2K7X3g9I6ChfOMoh1zCRcHDQJASC
AdXv5kvuamc48pzoHyADvE0u6O/w1h/vJq8rftJsFR6HgyTUHuQi1m+/E5HXVGMK
V6bouCEBFo6DlZdsrFlrfXuSw1GRaJPDEhzBg4XCFt0WXbmOrpFUCt/uyABM7euD
bOS4dFcFk1cHGjo9jCE46M7+p9Rfqezt+WA7Eu81ova+NfdiotOpr90cpHsTrrQO
4skct2MNUFIQduSOHP+Uq/m9R65ow708WjdLamK159ofT1t5+QhXX5xVGxfcntoJ
iB/9AKwfL4zx7/fy2eqlVPw4q4a1Sf8r8KWOsJLuixdmNNlPhIrJfQw1TK12LMAa
L4hDMyblWaVKE9f4xnH7XAvrMklpEJ2aQrCBo4ApTzAFSaO696rjJSFAmPvVM2wu
8rDqQlcNNiOQX8qbKa6C05OYKQKBcZDReeUNdF31KATSMbP6r073kV0reGl5Yel5
y2lFZXnkqP0RyvKNfeZYh6HjH3fhgBaYa2iALcWvpX9G/62NcR+LkhMX+m9HN2MZ
GLwSjJ1Caogoy+b0auknq6kB/U5MpIBBBGKtFhyAQfR1YSQjGFvGq1/ef6ME+azR
akZKuQd6qnFlRoYSao5IWqjPHi6Q2BWAXWIP0OGj9TjDtWYrdnQCHo8DUERFu0jC
cMFbgjuGg1CFOnZc5x21S5MKOiVExN3Sw5dGMz/IWMSgx4S6TQW5gs6GBLVVPwUQ
XY82eixKtr8l3V/UGHwjHWU0aWPD2KB+WRWnmpBJhVPaSaoZRMSs2Zf24WBxUpXs
9rJG/J5zD/GzPuTu7qL17Bzgte/Ns0gjMRhjwvZLDKLxgZSau1WuoJMzD3wBstD5
WVXvhhuPDawNW5DNO5mZd2JfzzrN3Q12COtoib5zOXuUnGTCen+0WmCoPmbomS6i
29PJjlGwXhQW2BscIZqZmlxuhrCjFoMSKKSJ5toCLLEwFfmwMmiS3X7JikpQI5B9
qMJsB3lshHFr3YoZoJrv8dHpO1Kv1E37lZT+Z0nwC/2sjXPP/WHa6xfMDN7Zw8Xh
X75oE6yJe1XRl8+prae1A1oq2jaXSJWn0nny8FDnuYFIbHUPEZPbu40cd5abZNaF
E4IfarQYAAqfpAsR+64j1539w/6HWKArC2I1BPzzm4qknw3BgFoiQJlInq40u+lz
22pLIgRW++Us+o1QMX8PCorQJmX5d0GLUsJL1P+zkP7WCPoB8okS0EAdHzvPCdjG
XSeOQd+DAOXF8rGFLX++gEwhuReJl/9YT2dwB/qg3H/alkG/0tcoHJu3sucyVri4
aKU/7vVMHr4UnyvoZZ0+NKZjN0YP/yAKmRY2IzuIK7lEfBxCozrvMXK47Ul21nHQ
MUJ7EGNkDluvM+feQkMpCR6lXNXy9s6HBy3J8A7vx6LkGUFUprkGB95Mymaj5HR3
0mNynMLLxdV+fiwoN4ZaznvzQC6x3WDEcREFUlyJY4kOn9MKLKdN0qzmjA9Bz5+K
JLtBF/HvOTt9hwJ3x+R1lu8BLLY2zUYxYCJN4RDQvYZd4TenxrLX18K69uKigixK
i+aVst7YUjA16Unel7G5ZWg7eBU7wDBKzmpAkoeQumLgoj45eVNIIHkD0c2aVud0
Y63berTFN+REsqcuagxFF+GbALtGhYKopxckkpRtbV8Vi7W7+FKVLtAeIGTLZbh1
QwShBNSV8osh6OIJLSCwZ++zztqnJ+WD4iiv3dBHlSGTlmwTUs/7c1GcZ8Ge+3xZ
BNE1QwB7BKnMuO4ufQUZJyYd6hohjxNsW/8wi/3u1tJEDGPoKIN8++f0lSK7Zezd
HgO5wi7sqz65mf6GLIelUUAvsxFZs9NtnTleEDiTJHtwbcz6lOubaiG/2bF64GBL
Z+eLYv2UevMU22FKoGTsqumFz11RBtIzKOrAGdQfLuS2ffAGyZs0x9kSXMrTWP4P
LLiEVQEnsmhKbm1q3T9HHw/iwOLfMf1KhBBNi5a8wwjT4NF9h2VHxASu3jqqbsdF
PUU/uH5nHQ0to2YScJdD1m3wujd+OXywONJH1ELXm12t6LQMfFf8Nce/NZQM7To3
dS0cAwkp2DTKLGv8XwlgBRhGoU7iFRn2RPPvn8KUAJ9qPJp8dhs6w2ECiP82/rvP
gKk8FL9SwCIM18HC4WoiyXiz4tNDr3Zsctj7W/t6QikBYpG7T7uyknWaJ0UXV2fY
M1Wq3YdHWCqT3gfuriC0qInCpiaABOSsJT2eimLF/lyQBhXTUrPXIBx6HMRlw64r
u0nMV04i68Xg+YxK5z1Rad9OeBw/IxOBP8t1Rq4I94bqSNpbuproeERO6dY0sFn2
cYKiPWDJ5f4aXiVav8m9W3kNs4C5WtVghwYemDI+lHK3n/g3otSTZEPvWb0xy4ke
PG2VkvVnJC6xi1FERnhn7AqgyyhIjrNlZKK5LWUWT4AHqpcxHJKze8QMcP+ZrsrP
PsJBNcOfEgkgWw3R6Do7l2Wk2FbC4K7rnOBHFKztP270OMKrdIl9f5qwRL12dQyp
3BVOdd7QQ3GDeilhPxYxw8xme9ULWx50nHD4Y8BhmHqPP+M046aTlRhni0R9h2v6
2nRmMPuycDnuVnSZiyKntYGDFrGNC1Z8E+Ow6csMg0u8+kCQmtGLeSgFZHSRGQv2
sQ33Nrr78B4y+wCEHPw/vVWRB1TjRJmM2sl0OXl+YpbEYmKnPc30Ud8ufIcFuxEi
IaPEePpMXPgMh/jaGnUEQtJwUjn6Xtp2jIBgslbDj3I6cxHj+kJO4NSDqibjuBfn
llO2YF3lp3FWkrx0ykW409eHKcz9OTdFC1Lsb/amTArQQfgd6q5Yo1NlqdqxhV8u
yADdsAlWLE8/3VrwSyD/B4Kg+ObsfMnJ0LEMylRHiwbDBm+h2+nSzcagZh1FXrK9
oH0IzBz1jZ2oxc65Jq6eD/jTEVm3bOR2Kc+YGFd8OpG3MKbXs4keOkvN653ZxKLJ
ViZmL+4wzmJDL96AQDrUjRZ/H9UGxlcundG4WI56fCg1Mb1JLQdIqzaoYdS5HmPi
AtxZKIm9OoVoaJL4XFgVxWC3R8F3afzGVTrQWf5SjcRNWZbvNq/N5auoQj0RsBMg
2L7tlDiCUqe5a50Av9vSff4TRlnnRJepbjVbFhjv9yaXP+JPD9KBDvdn3pwFC++4
YiFwmWuVPNoCR09ymu50ITO5pczAZ8lURwkY4Hbk32euIXdf6ag8tcjBEFbwYdSv
YSm99i65WK5afWvyhAQLLGLt9BgCB4s3xn+3F+LNUrtAFgKk8B9p1VrJtRLK6yaO
z0kh2tsvEEzz5s1fiqGMhVbMyf+3F7aV2pZSBv1ZB6FptL6wPEF584vLQR1ZjZHF
/qUaklvVRU1sdo+YF9k7ElTHtSa1C5kAUZQKLGPlhmszJTzFSIQwkvkSMKQk8eAC
XoW9LWl922sMP4muW3LyLcRda3vjhig/cZpEc5Xc7TKr+PUEpBlbHGdYc2Vi6lwO
1KT7w+laOePlYVjCOvaqI66LrcyP2uMQxLoq6DER2ewPYQ4IUbPXOU4Kmrd5FYww
KWXPGrMMwODVNq9Y7b1k52G+Q+WsKBa4JEZbiLXflkYBD+MbCUzsEvvj+Fm1zu93
8S2C0l00NCx/kRvUs8KWvLIEl1nGLeX/9fgrFXyiqgwCc0+A60snhhpDJzVP0VUI
w0JTMDE4ktYrUR/SsKdPYVTf5phEzNqAx04iy+NBRhExTEdrs2/1gzaL+4BEhIcE
+vXIj14JYMNZBtFwwFY5T8ZHSjRU0d1jfJyDUjiYOvbtw2A2HJvEjPZvodd1d9o4
B7h4uVKbZ8n6leyoq5vYaYkV8arPqbqIw+7fwAWKzk+rGZGg+FZRbnVBJBnUhjKT
I9brTGn7KwnPgV1l6a3r4G3HZYBo2xwpHTTsH9whKxXBzmeOShCvEPW+mwaIOOCf
qsFfp47KaZxstAqU0yWnqR7350n0S1OY2FOPJi+k4E/Lq9lJQKyoQbd1DZOBrUOv
lbXAAxoD81FHGHyyxYMnnN8uN/hyg39vzVfyqZdfY0f+0cZ88JlyzueYD3HwIwm6
URKAg/4pEMzHFFDfeOPC+pOjdRVTfRvINtQ6LsRQw+OxQKrBh8Jf/SnMRcu8eLpC
0tD+jrPVnh6zxrmUauxIikUUc+Z6ehfc1uWAWUFbin4NcqBSJFJ4zNvi+rZ2o4KB
kVt3nWSzXlLDcryGwYcNxmL92PShkOlAIq8isaP0n8+/eP98+an3qhP+1gc5od0T
UsUUDBceTna3wIydg9Z6EuyMXOjg0Tal2wzBVMqQ6F/0t4Qs1PqgtDp5BS/C/cai
Ha4yW2NSoDgw/ht40ssoWQAcuZSJ91t3tkCky0895sPiuWF7FQLSdUfcDV8lsyep
6QLYQWw00MF5S7OGBl25vqAyZiCYnK5k+lkEkuSQsZjZ0e6iHPq9p5SQWUGZGKin
/fsZF5rRsi1JxBkubiPPoSSJu48vWV0QPLYXfvWeFLNGuPYWtD+OphWVufRKULtz
i0KTxYEd3kop0YAs5T3kU8Ta7hRVExAzXwGqxUJrwCuSh/Lu8qKsEIrGx23cw/U+
EpHRQE4/x44GTFuvUDTtzU4bGyHZZ64q0Jc/wBK8GMsMJeF5O/L8E8xXw2dQwtSn
1bQYn49PoKUYHQHZq+4C/xo2/iI/R84vgmjL3eKO9nZz/RSy5+DzoJ491c3JUQrG
lrLSacrfvcIxnyXFp7dMYIXLx8pox26j80ysvKI5aPm4jJyS0AL3+TIcQ0IKh40/
MmyC89xsPa7HYhivcfXYvCqhQNUKGV2Evm6cacXmBcW2qo6LwogKURBOdEbMQrwe
Ba/6m3PXkvJk7+nqR3zWSgZJeirxRF8LxzmA2WT0eOdZssmfPOQn4i2GqekqT9Hl
Vxm70GmvUKQT3CU8/6m7rqMlzz8dhFypyiCjZ1FwJw//McceP/yBmq+9KJzcwXAV
c6JKJXxQEriffx9V3IPNfg==
`protect END_PROTECTED
