`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0poKzG5kq6QKG/nUt6JY78LabSVvRlBCMtyW5rY2va+6ogCrwE5R79Wvcxq2O76n
+24dgI7PIR8H3sWQzCU0NJ+oXDdHiKnaAoxfJUSPdYeOv4XfV+GznorSxn7MiAOM
FenjlFbtjq8zbzCgLAjm/DNK70FdqstnKIiSAv9XRTQCuMfoSaWrWc86o6KYmr+B
RtQUjcl/8CCNnB1liZamUROzddnr7yRrOu9YBpLkUqC4WMwXxl9OSkVUTv8uDXl/
SQfKlLKjt2XjHUg6lgNOLffKo87w6YM/9b97xEyUFNfjpeWToiKkmuF7i0Fjza09
8FeYrwzFK7DGBjWoDoo/hKBzBR2UBhDUoO3zqwzJV2tlrKTueXJwuMcGeWQy1qbz
ySd8XMuhjyxEGcIrAM0OBa+lH6lNQO4cf0uphyIC89IaVC6Y7yx7ojNwBeFdAS5Z
ET7QNUf7UQFAsdcH0TAllUmHfcfiW/ZNLCcmtmqQBgONHHIT9TSaijtIfK448khk
XI9iSCL6zI+s8KOcwBUxU8BowFfhv6w7LDtHiVh6MZvDiyPURJ59kWXvgCi7GYak
rBHbB0twEp+tGmCgMHjsDneCqlQ47y3bcvTQi5pqB918yzuFo26IZXHPyiBKWx/h
/tINGXPUAq4toCm+Cot3vi9cN1YwnGXh9i3mGu/+HTc/sGB/uBv6Ome/pEHNXOmE
PpA0r6l6x8WpgqIqtsjFsMymerz505RsLdsoGXVIjxBmvuUnT9M1TLACj0jO/Ftz
dlG6xewxvlkCQdYbo+hdNkskKMJeHScdMt3aXVREJp8wqOgGUMu0r7h6eVXMnAGQ
jsqN2s7hMRVUPuh6R+eykuQmKqzeHuhKAsWqrK7eD/H7JeYVewXAQUBJjodfDcY2
srziPZ0oW9ehYGxzsGmLLmXYFNV44vMyaHJ5Dtpba42zhHZrdvivICcW9HW7Gy4C
jdr3twz5A8BbfkH0+nxpgXcENDj+jyb6z/aX2TKIxu4+jmN5MpKJk98NjImhjqai
GXo8EEWNuH0pDwPxi/05tffL/CvugctF5kh3uN/c2EnHeB3fhUVwQ8gmL9GsHF6k
kHoJy+2l5abHrFY0BwPvn+fps42260nShppmjW0MtcHi4bKk1+p6O5xPAEhwOFoj
/IuYCfWc0igaPwRMwoYy9VzMssimvTtmvZXzqMtzL5yXS4gFzVMkq3DK9E/SK0gQ
cLutz/VwBR7vsfIUw6bVHMCQOP+8urr/22DfShTwlWeKhcBt35j9ZJmTPY4GXi2q
qkM2jGwHSUS428IUl51PVaBUC/3Uyq5J70zyQ44gC4xMAXbS0yshM+JaMF1XfigA
jsS9SqrhspNvThEHg/Y3uBM3P9B1ntl9nhURD1Uo5aIiZ5AQtVvm0PQAOi2L2vA5
b/nv5Y/N/hslcwE/inKaDHHBgiUCowxsifdLxK+J97cz/TDt+Bh5a6auR7doL2Zg
kSY8z27vpGvymWFH7y5QWq9OYMiUdr8jj3sVBmRSC24Q2PARA6IMEk7LSaw6Q5TM
81wdoyEOVNxo07OukOOGvp+Mm7AYWmTY0Ive0wNZapBHwXcfOHJUCGVIG6eK4PnB
xNNkEPv14hGkmJWYy+i9H9md10f9Sd+Msf4M1KIzw6gkfiLGlFncipY/ngF5biRJ
b7e68p2h5A1orMh/jYyXqxIakpbqzBCFHaVqglaiUsN/fVjITyRiMiBynzTaBEsi
YZ9M8aZc+mrzlPyu3AKw0uI0dDyqWrjCT6ycrBdYNNC0Ok+q9ALhs3/ab2VGKUDf
T4itVSRjTM4o6etzowEuajvbRlNSa9jfZvy7tTWX03rYKsS1iEN6gOuSWiLTSBu3
wYwqz2rcNnSh6ZV9eYHAye1bygOfNdsJRC24qlnAVB389ylXRR6mirIGjvvObW42
f7Rd3CsoLAspfEsORLfaaHhx6bcay/bHXOYR3dg/DPlMFRUnVToVIjmIHeVkbVi+
ac9+t3H12jt3++Q1zTJAQ8cBlG39Mw7Cz6zRVMur8J9lvwlvDFKcH+V2ib+q2lo1
BATyxq/bGVqpmEPVcu2Mma6o7N9U4d17pQt1Dkgx3RqTMlh73YuZQQr/QmzNdHF8
vuUOg+O2BVrD75AJV5qgixsXBmngXE5QcdchcSa02ThBfMAKsY70Q1crReMpNSzo
XvDq+a2fry4NKAgvCvXKkJ0duMQKyOjCwAi1kuLmHY+jnPhFq0PrwfOBjy7y3f1q
zCIB4g8bwXBhsW65LhHCO4FNOibMN18M1OEg/avUlXPX+QMKwpJIe8Lo80rkYieg
o3jTEdw/JBpZxkkPBLIblvj9Xl/k42JxKoA+M25spHcq29+mUPWalsrqDBFhbswf
nWtcQQLdBmtzLWgPW7PbZJ14c9+nZxy4tHcfxPE/e9SOffOMSl1sxjuYl+yiOH6E
0AvKeGF0VOWV3jbYk1Bic0WnO8La0uhGSknjPoDNvk/A+MGz/YzPMCob4A4Bv/wJ
Iqhhp4teXLO/gZyk9kAI5I27xrsqre3y3buqHfHzxkSx5mtc4/tPC6o+Z/7h1M+C
UtZJnIdrGmg3lZU/dZ9KiB9tWw1Ka0I0YTaOeojJkCR+6fDeSoCSX8sHhW9PRXnW
hmf6qOXFScY/W9R9VLmYvc25jCXmgDjIZppABITsgUiqx4eH+9VZoI+z5Z1ta3qU
r6U3WSkaprQz5xLUUNEckBUubgzX2gUx9Gzylis0gC0M30rjANPxH/x42DLuf0eK
DbLlgilRRGrakJM9IEpzzwkLpklWKVPlXX6VTxWNrX7zSA/Zr/7SbBCEP4G/BbX0
JIspLVjvEOiIz0DOQzmgMjvzvEUxZjo2u1atJVQ6bXtB80jAV4Mce+1zEdeWxLsB
hPv/lWcyO6mxKsOkQfsKRl+u0sRoOB/len+AQUYWPN+ltwCfd4KPAGvUexHWqSk9
Cd+zmkN3F9r9ttr4fkExZ7iAGt+l6sA+Wnm4k/qGCWckgpVXFMUyoqcm5XxlEqlL
sPzXto8hAz+ndjvs2mkreGwK6nHG/HTxoHNrue8+qR+qx6iEr8qFDdfjD3u72eTm
bowai+XkGRmvl1dxXAJRoRH25c2mwmxcKeHvGOgP3j10ZiK7/FsVkXiaqhDfgotj
oR5Q1tOE4a+9LERLVBmgDmTvudVZpNqCEf01VvWppYlin7t8NqHNyvXFDwun7aXf
PxecZFU9AKMXI9ODVU1PpeI/yZDojlbvooXfMpa0aurpYRHGMwj58oOA6TC+BgDJ
rXfOMdwkMoV12TT+q14OO0X+InePMU+5fJ/jBtv8aVOgFiTVA3GEKBXSTVBiGIC8
1xZvYn6bVbFaIuh9MDRx7ceYcJvpiscUelcrFo0sLYJLHolQybEpg2wAy0QJ/HiI
sPS1ct7TkEuOBz8033Y3/Jh4VotinfcnR0FcWnARdG0n8KVd9gvVxvlIaJL9rmA8
aU6bObp50l5Jn1QZ6Gh24pVwT1xbUZ79T/ogoK6mQhmjHxxKbq3lFQE31zEEClSn
+zAdG14LfUq6STCXwYOLVRmzKOUPRd7erYlTgSHEFB/MdF6FB1KUklZT1bS9XNP2
i7TprjjTWZPUEov3W8ueVqmGUZ8ap+qCbJ/Xg3t0uUkvZeJU48DpIStG2PMDtprn
ptHG9cGnep2RuqaoCyLcShnsDaUj8yeLn/Sxgu6V+ANwnSvSb28MmWRP/5xy/vPO
l/BZGpIMJRGInwA1b5DnWHlvGoMOCdEmoWEAhaL6pGxkA2K6qfxhyi88ez5mjYSB
v2m2m2w9pOml2VRMDFWEXvCOciRb35VvavD8Hpfi3XKyTptguhdtiVwmGYT8klcB
ITpAzSJGwWWm0m6Uk76FPGFA9N+s0t4aMDLn5HY9VUjwLzB6PDd6k3RXEAphI3IC
yeXsdAl3OYAXDrfeI5QhPIkncqfAA7kS8XYAU91lXpcvssfVlY4jZJ3hAQGmAPX3
gjvxCj2AkdUyfB9GGokYmqnVf+TuAfgGytv7lrCy1ojG/1KzMy/M+FtAoOXeGTrE
+O9X5k5XntBIC8Gbf6cnCmVk6jIQXbdnM9gjoR4B8jbRGahweYR44jSBwoL7M+cj
Ljy1CEY+g0LIhLiWBpkighp1tDTHwSB6KIfAIy0B+qIbkJ6n5sLbU94vHOEq4tZF
xwaFQLvJc7Wqdo93FlwjFjODKBSRu4yBWF8ZjA2o/0A1eNGOniNX2dfMQBEsKNTO
zWyzCllBj9VZYPi9b10fB+AqwNkPfwdkpBQE7oufZGuA7HhVoFhrH2vWSEP6fcDe
jTCUTs18Hhbxe56briiCJ66hKqdblltb285uIGG3amwoTS70pOnbX+dRLYVx5Vgd
2q2cBPmlxr0HgEW+MiNRsk8BtRLS65/1H9M0rxSC43DS+1YxHVH4A3yzVk5vsLkd
hOY+h2S/qPJzr0Iew1RXz0ghfhMP8SHbVHij6I4F+xFG5qvOITWae9BEiitRRrfF
6mJKxC6env40lGSNCtlGX44LY6jOxAKzxnqwYdkgfAOmPYrflfX/Olg+EY8xFEuC
f9z725tV6iGoeCQ9sPn4lGOEJOPJa9smB4RY2/oOJfoAEVV5vxnfKaMxEVj+aqkk
yoX65b0imlx+W1RPsvFE9X5gAm+Fm6s/p9fm7obSGdgkfbYHKdEH/FH/PmjjBhL8
mh4Vl/Dagx99AG1xPZQOk068T8Ueo/cUqDnJ4ubJ8jwvavcVn9C9FqwyQgKxRPAi
mwrduCkuwyC8azGKeNtiHELADdvdas/z8Eu9nr7vIESA8yUYFTehgXvJsboVhjxF
F0dShjuWcMYujy7TdzpWzLZajFxTQuZ8XJpsAoSjpColgz9kNyHl19doaago1+mF
Cpdqtk7+NISsxa+xinFThXkyoFQaWOUgrkrZ3WHpl6FTctTNQ2QjmDfmcE63Gtt4
kXSGa4eaJ85HWnKxiRVPCvIchVQc+VUqUZc05dE4ZT0XUd29lKfQWTSO/pGoQO7z
mlLaPpY6P3ZyEQQdnanDgur+3csUPUsNi8d1qTS8cyQaAsJi5sE759/yVvnxfevn
6aDnl9TBZC4K/ybJjNTPla4DS2EFORXS43gbMyVpbSMD8hByH2Mv9gLy+o7E/DrN
zlV4wdxzn29y8nKOX5Ds9pvGQxmAYvYUTv+NTYlyfvMO6cNuazjnhMAw08VHyh6j
o2tBbyHqP1CksoY02vTENYk3groVPHI/2vzO4pVYJJCfmbI/C0i+CNS/teXQwGYo
4qVkLjinxC8JjpR9bBT2e3DB4Gl7/WNCsI1sBVFTCDuZGApeoWRuUbJMbBYhy51b
TujFQQ33YvMtbuk+v7NJcTM3Vuukwd/OzKrV5USWWfh9+Wq4hbvkDyI0I6uwhrQV
2Nm9orkPADb4k2q29gHZpEDMB5xFbGcxU3nJE30ZDRVWMVzJTY7HJsQTLLJ1LfPf
mRn+156yqmb4Nun4j+Ht9V1L+Cl1RenIvNt9eoMSKz8iIWV6JDUZxaKJfDtFvf4b
26LLGU3snBbCnp9qC38HGIQLl4pU9HgrLsBGbbzRGRlZL1VA2bHi4yqPANU4WgKw
TRqjEx2mC+HUz6PMDeufoRFMmsHjv9MLFugoiCvQFDxukDcV/AZOvj7UnTTg1VBC
3xExVLxN6dfLTmQzyDfy/+f+g/+FuDV8gaA5gmfOB6oRWp/6Es2M4eOOCTnB6Of7
sY+dTl7kLs6EH+8GOyc/V+TwW2ywL0DErfsoOImZ5DB/C1evmXv6x6OAZBbG4W9r
w+fR3eVpZOufV7BkNyBWtIqjk/dQoJ8gWbwC02Wdz7AmSaUJhQjDwgd375Syr7Ep
HFbAZ8c2kdTAqF/dTpmwMxFxZyr+dzh9S5wuTzicnEfYfdycDmBdsUX4YTsf9orm
FoLZKnDTUv7UGtTSLtEFhTkTQePHCPMV5AgujyNQKgdy4MwHXjgIfVWbGNEEV3s1
KiKWvu01ZS/DXXHOeV0sJ8/YxnDOFaDhilkIrDe3noCDCb14nR1JJoAmagwXYIVz
c7ofKP9FFIyBwznwjNFJ/jeaJj+EuYJ6I/YZ3DQnqj7Ie/XtuWEOrzrgPkTkdatz
HubQnuNMkBslGyDx1JzAh7OguUOTagexvql5PJ/Of0MIEg3Qk+Pb1qk+V4OZlijG
/7P/4RyLc1hxtMeL3XRW+WX9EKY/P4a5frIAooZII2Wr/imGlHqgeuxuxSCQqr+z
lbloyvuU2iABTmJGz+6tArLUwDcD9C4ITFzajx7iXpJyHvKO6BPMmULRiVCaPZDq
0SyIWP2aEsw9uL3u6LnCtsMX9YDIW2yYRD2q5Qvx/D7LYQyrKxs4qAmiV+THnpBp
8dqetDxIFG4vDzWMKF9vkbdp9oQ395t+1UlfwQsbQ3dIhoXQ4oEdA8Icro1lTvS4
E+vTAO8IZkuD2kT84Ds3eHDLBtuV1oTPodNRWJlt7DUWD4up7pmvubgclYxlY6Dt
SQ0dmIARbD7D7rqzx275IpXKWYIkbPFYugdzvoux6BBO6A9pBbzuCp7jxxbSji0G
MAwf+51MW+uv3gq6oC38Wmlr6Bt6HhfT/wed1eioFK/S9cTeXzenXKFj8H8lSThG
UV/HE7OT4hPgEz6AAsLrlTTY7fR3F2FsX6A2+i4CJBvQPpxljJQihrNzwBgbBSw+
7f8BFyC3meF3u3fNHwYjkh3EdqvMLR4+ge8EHfGIqkV/FQp/AoQ7lEnw6FzxeQqt
xEJgKG5LEkST+uH19euy55r3jgxVtIl6pDOwTiSoYK/uIqshI/yjW+iiJemZpWVi
KITmILmehXRM3k3Q7rPdVbVjD5kRPhaCoeg5SzKeFYlMCWw1svd420Smu4KLsTGR
+kdSehpUM8GSxrmQA2KqomzgwJrcTerghLcxX/AGWSK0FVy7oXvtBBCcwaNsLHOm
t/fUr0Is/HpcMcSKj1uy39sQSS3s3VnTFET+q8/tcGC4Gzp9vHb2L+2wQQQAUMkF
C0s7l1vmugTtwJ3g8rA7JLblrt0TR0CowwE5TB5a+YVfBG1wAPQFjLM7ioD7fPB4
k8X2jGXWa6rniFNoy5ocU/zdaByLGG7S/l6SnmkmKabwuQPi2K5xGDnaCzQCYts4
3asygI4zA+/PaiBb6sa1hQyWZt+qBdOtuUUu+QAc4g6DgSFjkg6cKZBuKexMJ9o4
3L4uEQ0N3O3McOxebtC2+iPYwh6N7LxXFAhFnDNp2O6ZU7NtuGy0KU3suskzvruR
VByXHgV/f7MTeek4EBBUG2zyhoQff6ObYXR75O1nq08NIfu+HvX6Gri9ZsnYSsrU
R0oaTbXAXOyWlZ6p6RH2g9MU0rrf2mQy1f9mA3Wn3f6E04sVrhJdIHqm5pwHFirS
xbZ5r9ox5/sZa0DV6aHgOvZ6AkxQvj4NkRjvaEzUDu9KiCoUiiiIqJ2AGeHwNcUe
wTfmZ2sE7LWN0NCn6djVObD3tpOEGgcz59LmTVRod1Wro/u+hKae0AYxa8bSAdCi
aa1U5RDt8pGkYioZfKQ3FZeyDI3C80bL7tBN1Pj/xuJ7o6QvYaR/S3TpyBC0HV4A
/PSjL4ResEq+bbjHrfC2jPMq/nGPL8fnkDSpJERn3hrt7oPCW07pD+eVObhXrj5O
daiO5TD9K0Qx+H50UiYNR3CIL4i9olZp3tAnvlrLCSuI354BAKAygFLfFRZRp9Lq
5KHVPcBLeJ+c3S8Fx0/D4SAPQ3QfxOpQF27DBWi2JuaayX9JGRqhtgMO/oKtNnnS
kABvTJJdvlP6VqgweHCq5gSQA3n+ANQJdTXqN5WBffjGcnPA8E1d0b7H2QP/SKkD
4UHW9Ko70FjDM07HFmBV1L541cqg8CH2vJ2Veu4nuZsOG5MMz18g7jnjuQOlsJky
QC7DhN49AjdiSscYN0KVToF4NXsVI73CqzzG/jZOGXZJ3Of7ifi1aoegP22zSMQ3
7R5GkrCQYHh864JZ+jkINCZUoJy5NL/fzfFSwEAIoo2HEfYUa7MLMkEFd0pS/ASR
8ZzqqJX4jmg2R9OJbX9CFWLbqpgJKEqQRbxh+OgmyER/MCFJIwny3uEmK57fMFZM
x8lgSNSa1NP3Jy2wZ+E5qMz+F0IkReH813vpZ6AqRC9wit0oPk8O5NvX8QNhD476
hfzWwni12lsds62aMF6arfe7HKxXPuI9CnKxilhkBIp/jctpR5uzUK46OXJE0mG9
4/e6Lz+V9h9HcvIkROhQGWI4Egqh0y0iaCr3+sN65OFQ6t3QUAZLe0fjBvKuv7oh
ayJ/nwn96H9EyriVZsQ13Sq2VzIJ+j7NYGXoirqjCdDo0cnY1X5SFZka72kChoHE
cMUFnBbpwMUtIdUZCW85pGzO8QbiYY/8NMA6N6ZiFood12EYMjMhk99ifhyzGR3X
s4Mx5ZZHCmy1kWYIAxgy0O7tWP3mM8jCJ9MULiCdPcGb1P5YURl+yr+sL7SrefIu
kM53MDtgRE8wgpT/TCg78rM+C2FHwpwhojcuJ5l5FJQtDaM3dtyxarDAxYb+3nNU
GIVHkFIRPKI5QJd6QwiBgrRXKpBpihTx/eYJYT9oTASi+yiVTKHPGZVa7xc3pQBq
RrXFw3Ixf79fIw1zUfNvkkDUo/aalMmy8UOmjLPKl8lN4E0ViLW21aJx20LkM0bl
Ec1t1UhZntkkFgVittmBdIM4feHoGw2Q8qRq586PQZMUDnW12gr58DuUtNn5d5eP
UQrhuxBKw4DR/Pqs+hIEqYunx9uKJG4Wsh6XnPJ3YkU5oEsuLBIPk6cxHaRzwKLt
XQvd26dtfkiRSeh2cdOsvVt0MHX575FcOfe5rk7V708AVpyTlK+jYdNdO+1K1pYD
Q19317ikaE+giIDuVe4HyDWSU+LebncyVtsIvHrZAbouSC3KG3sko2N7AvyPliqZ
Ftp5So1Sx/PqwHppXiGJc4lXnkwJZxDRX/HMpOc8nmN8P07TKK8shtO4j6Cpg9hK
ip+8p+5hdsWMjPhUj+HzoBUKPv4Et47gtHAP751irspQEMH4l1FQwT2XI81Hsz0m
5h2fYgRiLieMjhsGSk67KWJIdD3etcJnEXiGjM5+m4a7Nhyni2TUglm1yJGZoAU2
6A7aorgwS0bzTQaAyln3vOY4NF/fsrsTGquaaxjROupWkTw04T0AeyRS1afGGLVh
qtMyIjFZAH1lxezqN6bvZ6o5AE75zaml4WUpK2NA0r4y5G4bZxfisWWQojD15jGP
PlI9UfMYnwA1Tx1dDCEOJLy0Ej05SmJr8TdM7YCmsNAJ340VuyPdfsvJTy7XDvVt
qPt/n4Mol9/yUqL4uos0C1Y+aRQk1tBJPLCcOEyB/3PDsYSADgJOkgni6V2oxyss
Cr8GWWXJEd6tq+Dc0ObBZI7f8DSaPleK8Ddrwb69fpskPEIlnInwIq5b7eLlcKrm
LUIqxHD6nGnj2IA3yX5LPtmlgzAde5y44hDdzbHlLj8vJvQKCK9GfxJqgaDh5hxX
H81L79CGqf1IEo4MQxR3a6R1k7pkLAOjGtnE0hKlxNM2SSucsQUGaC57Y6hnMpaa
vpH5kIOd8Wh0A9OgbuFId99fcLIN/jIHIwrtBw7h6yez1XswXk6pzNWdWx1NRraM
qQtStxyyCnVeiJYQ3+fGEM8Fm0S2GucL9fF6HMR8AmF9Rdtthdrg4MMVxvIIrWt8
eV5PKuIEDPp6MvL5VNUlCZOGixWM9JjAJ7mQmYm/aylQBgaoBzb0oiXKanDDam1F
Y7J2ikm1b1PhNVdijzzqOrmEi/wfNcrupnjIu2GCpBVCxhCUHRg/li4oOjrTM4fe
9iVHhcAEuy1NmTSmMTJsmiYRPHg7fSFPL5S03VE8+BOFcogK6knIQ08kjn+VBUEP
PVYF9wfRByhcEUe/kmnbMrviIxpx7amZ4M1PD2SY+3AJLCiHnVcl1WBOTsQ3pQe1
KnfJh/9USwZ8SrxJWZK1vuwHuhKyYo40B5hAL0mIB6EaXY7y7c3TAu5+45jurCB4
edJywL5GoKAX2JimFalg78LJ3d4BDRGIWJKzYnc089lyWpXUT9VdIHg+blc2JBdL
0YVJSyozHlmxLyYB7LYxufkjqIy88tIH+RrP+miE/5bVyqJ2LJ0GS0aE/EREZLJ0
bpagEo5iqyeWbxD9B1as/6M0YKKIe1OQ5GfcOItejseD+AlbiPH576yv99414gQN
ZGxpUm7urm7JEbTwS6Kt4f9bXvOg0WqMHl87f61FwvChrUUNqVP1kpZg8efBVrFJ
SuKxs5hr6M0Clrk+umpQ154qOyKCsVcOTQ2CHKPI8FJwyonj+RmNq/9y3QrjwOmf
lBsGyJ+9R3oXXSAOJNN20N8jm0acP5OHAgwEkKAn6CE51bOaLnFC6XWArgrk4fSU
BXrpKfc1Bhz62GIHBiq5vy7eY/LB8F8CWZ82kao0pL6dfEpT/1zji+YXe5sHuP2m
qdpxxo38FVnWZImMW9rJdlariQ4Pcdacf0OOAU3iP+QKVm4fjxpVrys3DvoJzx4z
q5Y/0pvRPtpVqfBej94YEAvOu0lKSYCUO2iUiwXzXLGbgaSK/rFICXp4/+jVwFpY
yPOIiq66z/no62n/k28qodAFCIQrCWQbhlHyZdcx/1xlGinrviiNL1zEqrP22byP
sxte5FcJNPX6xCaCZ+HohnfjKsFupETrLvIFh/5FBnrRDwc7Xplv1jDLVgSQ7hYt
q1U8Ah7R11sL0RR+adGzOSIACZKJTyIAOYhyVb7+4CLM0llos+UG0EtnV+jB5JiU
wZPtpsGXFKdnSyK22ZU9PQr4fnZDWiSzDnJHp8JkP9fa2k2vP74WPue7aGA3TQfa
mtsEL7MwNn37ZwJXWsDbeevuQXVVKA/qmeN1LvRlec7QfUUS+Ecb2g6rg0/4uLgX
DX636GdZ50eXCxLGntfFaiunLBG38sQnLcM6wIhnxTe4076d4XT0tTxsgzHdu0n/
h3QFOoCEu7NJ1CmnSgryL5hcOVTtnDXSjI3/rHYgq4wh3v0GjzktxbyMf17y3U0H
K0Q1FyXuC4LWZFXYH7jR5BPL7No9wf1MfetslPwbXJkPqGtsYvgsXC1pb+DNJhO3
ctjM4AZAyR7A0yfeb5CItFvjr/qT50dzbbyGXm1Jo4U6uJ8xuFO64nmpki5bF2n/
Q3NY3+3QiuS+0CDMwjbrD+ZYEYpAE+EjIXLPNxcElbBRK37dkHygFtZWdyxq3Z9O
uVeH0QDbcPj9CbwWgoJZUiOBe+r/5mWosXXrIUXuBEbgc/WJGLjdpnng8sQUtqOy
bTsGi3BIsSovpSzML6xWh7WsyH4NxF8fACMfXlb1Hauh/plezC/Ba4a1aVRwXPIV
V95VYDqNjypz9nH1oVm/M0IYKmIgGfc5mOb0LRrRDexGiyQAQCs//FFTvxt6BCiy
EiEOISJzchdwrluc2T2El2QrdL1mzFM0XCDpXYpLOg0TBjljPi/LMJCLzbHFHtz/
2UUIjoErhxpd7QLcVhaPbkXkOOO7a9KVgC96APv/QYD2Me3uD7PD3cf1txDAEkNP
AMt1hhHl2tR11nPXH8EvFvk+CwxYE/6ry1dhoHIBjMhoCsJWi7/IlPnsxpL8H0Wb
mj5wIP+Kr4rPqOL9n0rQKA3BDaoF3GK9zCAMYqVq/KkTJy8cLlv/IBKjyvnDDDga
P0oYnaSJdwtJF67+Ks7unghgL0p8x+NL2iLDQj6XM7KIzyYUG+aU8QsFt0LmedIG
LeqO75TfMOlSbbmVHbbF1GPmKHyypinIuVsK0w18HnKk75+jRiXuL2TJlQTxGzg0
vDyGSqt/0RinuAIbiAvF9u6xbYt3Iz0SB1RJIdkoiGQDz21D5kf+JxkLgxr/HVG0
fYBuB3swykO6QlXlco+uoLxsb5NULLVuqzI4QuA86yOF3+OwtpHNstKoLZ7zhjMd
bAihissjgeQxpF1cJt8MWWWw0u1LUyhKkMd6Gu9vZDPi1CBB0gxjCmHlN4lgD7o3
u9Sr0FwDBpsz/quAhAQcc+qIBPOM/Y5UERd6UfAl0Rw3V9X+84dbTpr6UBSizlAv
brpRQdfcuXwaiWTahvj2R5m5WkjR72WQ4oyu2eT/i9nLukUTb12A4GTOx5iFRWn1
4SVL5jahNi4hJOt8Bu19Jjap4jfxBvJYZXuGsFvmcfL081QXVzOYOqmHPNNqd+JA
3eXK7msyZG+eZnehcS4cD6SCIy9e6mJUWfRCqzpx9bF1+igv0Tpq+ZlKSSIpQjic
z/3acD8aGQmdy0O4SA7yMwkVDYenCXaVvKte0LxyGMVUnp2Qfw9gPGKtz4/U/TM2
plxhG2IHjRipwDtguvxTUOXe2nuKzyFmMEICxwqyggXvUY+jvhzUlQuCisGnNPnR
MZsZb5j49ao9R9u5ZG3bjOVZEzEbQmUywcuYXGEfBKlg5qm3tT+wAFOZC+6psqCX
i9D5tf1IqQqBfm4LvMluDzHvqdIkELPhqyJX5REfIwgXNitjNsJxr6+dyKSSr6Sb
VdEoiNUlXiPGa8KTk5+5hE9I2UKwsX0qFDiY+Skg0i04++dxMoPM8uSk4RBMKyRi
Z387RcCpJKcnnwg2Lc6bum09XL2gS9F7hIuXMV0wkHHIaHjn7b4qBkt8hxpmvuoS
EXBVkdkiH+ObzOpUQMa9CS6f9qRzDnspoT1PYjZziw0kWjheuVcTm6QRllQ1RVRu
HHBn+v/t10F7eiaf/xbBZ2muXb4VVw+x2STDdeD88riFvrfcjYiyrI08dL+i68eZ
rBCyw4GKpmQ/h6tmJTg236tLAHAHzb2xx/vuLf2nd7CPo3JYhJsEa4wB8LJzHiQc
Dopfs1f/uJWYd2uJmeaAcnVfv6Shzu+KtzhvNcSjX2yA8ZCk3rM6E9I1hmWSeVd0
Nt+XncvI6ccX5RZMctukNJmcsf6a1ye1N/wU7odttrgnlS8t2Ca6DZO2xHm9VDtr
2CK5VwiYRKa4gNwVgCbysdNSiC+48bHPDJIU1cYRe9Bp+OMvRC5ogDF4TqGr9nBW
eRZk8JmHJHP9f9T5EtH8JfbpkuQxpFcP4QcAjpRqiUjatyfVCCE7w6E7Oe0j9IPw
66wtBMxWp4X0NYg5YydzwJbnyOD++n5bYImkS3G//OYgVKtI5zxzsjqUUs5BGlUd
p/NtIvTDiGOhCf0eWvfUM95gFv+XlEEH+PrgVYbrBQzv7vjYGvn9BbhsrdLOmShw
a/8fAmy+VZLNwRjEEnzcX78GVikSBF1HeNLRkj/Du20/XkTpPS5sb0ZeKCOUpP1q
fGk6lORtKUPtVZo2Ep4IniruIBp7t+OQWI6N9bGgIB/DdZJQgqZnabJPCFDM0OWj
KpF5IgmPXuapRqiuINwHBVxL6nYMBQvwUu/AZ5JvRnCfaSLTBTx+ZCN79fWrXyxm
mFixPPwcrOAgnkLKug0P0CUaxv6hFnTarAjwCv8+AzHTgVlyxmh7DVH8EQBOXRtz
N8sD26LoZsgRsEewXOKo/HiWE+JtHEi1kA/40n2xXSQ7b1RHNHeEDnCApyinbPiS
8IfiChSqMWDKRvpAzYWp0NBZHK0AHDB6dUZru7JcgpNxEguEd1b/moqIJ82q1LTY
9CEvBPB+pOCAkK2xQwq7ClRu+yLYqFg9obSaSszmTY3sqqOWcWGsilHHGEUD2b1o
zjSZ/6XuViwl/xx3nz4AzWvhcC52QghoEzEaQs7lCHF2+kiZgraRL/RL2Udp9x/6
HIwhon66kRlrYg0FUEMEwF1lfJ4Px1kdJBpaXYTIsqDgAI//6uVyYkrYExKpURO/
Y5R/eecoRGyEBU74DfkpUOYtYrGLSEFiTnJWXOdq24UjithJOYlvEH9ITWX7GJSB
8GN4gLjrQmNI4eFQSXhoXZ5RVPiBgG6HURpyt100lPFJf/+WafN4PG2yDK+k2Grn
iHFMzx8KI6sQC6hVDNE8aWTV51khir/AiJbpj10MdE7jf//ZmGXWrfJ8s2OHbRxw
b4ypCvwg80MauTUBlBrkarKKV7uG61EgI5lKO0x6oCS0vFYerS3zEHdyC5e5nj7f
oyrMoGqh7FjSPhUJZxEdi9KSFxRJhNBUzEXVxbygyFzrAEEHUGJ97CLvtolZ8lMu
+QVJhRuoOaiNBqXpXHgJV73AB1wzhfSH9Gm4v6b0GDLsf6DIaALtzRDhRrSeSTaB
m3lI1nNRdLflF4A/nnYajyU5pgfHAxVgSav+cg9KTVKG8+kOE2FPt26VRtwiF71N
b3xa+BRzGVwrXZj80CjLpIOBJt5fnvE9kLxriIugNOTK3VNpIAf5Vn/k3fuzeb2z
V3vRiwjgrEZdMtZ9pRSHI6fLnr1GjmaTXGKcJx5XQfyn9eYiOIVDjnQ1K3BLolts
iTrHu4zzHiCP4xC4dgjH4CL9VcWmAMDB/bFXyV6fRqx2us3aHOnvmPCqkuUehHh2
FnQ0hlFWsML3qasaIHRIaXyJCfmXKpAeULxQRiQFom2lOhCgbniidgiMKxZ/SsbE
3ovrbQXdg8nPTF+FM4pO6QkD5eVtNGJFIvlv+PO8SlNw+4orYraHllxIW73fEtbs
U2E2axPIN5Si6KrNV8geJ17/YxQiW8I1sgz/gKakWGfcnZvyt73BTkEZ/5uquo5M
X9pSIVotdbcI2622RL4NqRXanEmn+R7vVbxdz2MSzsbtp7leqe35YtWvOnaKO/rs
jiJBoDxffXzKxg4G2rnbPDw0oLyhx2nEMa250n3UYPsFiixHkSxOC+3P6KQob4a2
TXzT1WdbhDTiPIkyjEFjzBdXguL63Yudn8uNBjlxGc/5574T1LW5WEN1DONFyCZC
uJ6Yxn3hwKKLtuPoTbF8Ofp8JX4yaH0IS2pJ+W4UO/mR9+bm9loIBARIubnmMjhK
6QZbjsLkiF39o9Tc8IDHQnE0OGfbYAu3T+GXsEURHzSZB+ohz6Sf+wI6cD5xnIFw
9Lq/KmpR3w/6b+b9hBLnKxlxLh1dN8GJpVv4Y1YhWdTYcq4rVDtgOyBI5iawElW2
NQkOvN6F4d9sM2y+GgnR9wGkPQGgfAFBQJYu/GjmUCA9euEgDlUoIIVm1uY7k4w8
u7s8syUq8b+KQLyOCJ/i2piwD3NVzVi5afM0TLOj0e9x05K2HLS2PWxjJAOHPwoa
VIRzeHe+EWdHeBVtnFGquoZ8A+xoXJsMuVKYOeFKfJhMloSCIJuHyNJxvbz34iMc
pj0FxPcLyjHsJchWAoNDqTkzTI7v+PAbIzTWbO6xJoSHKymHNHy7gzixMBRNV4N9
gYrrsaav7zCnWamnB3hCB7LmOffeHi+cZJkh0mgQLjtmUc5zXS7clr1Qgixh0MxR
Yjw3GIsO3ppuELIeiNqMK1MmXRygAtmnspn9dUqA8EoNgdXww/i4wqC6mvjxEfoZ
zJJ0x5lD0bFYjT2AYGO2g9fxzyPIRjto/SWhIQKIMJyA6zcNseUatzfcgexleFuc
KkumWPmdK2zInIw1okvktCUgHMFflrDoSbjywVMFxZ/Pyv1jn8NZKUsihlCZ0Ai1
//A0qtE2/eqVMuYgWw8RfvdDPrPixdYkc/Cd6BxXhBaOMMSgpZ7UkcUnxo+01GTY
5h/T30Dm5Sjg6alf60V+zqBAO/rgr7X9knrVLUQDTLpEOVCbrFcX6k0khxaw40Bj
KgWcCr73OgGKKtoMaw/lkPAtpS/0aVKzfxib1ESUFocVUx3a9oc5kbHPYmXpdc6h
oB9BuShrTFKByYJLXZwfrEu2K78RoUCJgGB/6AO+tScwilil7uaEipvPV7KsrKSw
IieYZyFRg0UoHmZacTz3z8UoAvciAuEEnfgJ9gLqJXb9JX7++k3HWVfbvWYlvTe6
5CFfBeqwZzlqaoFakxdU7Kkuxz7EFOBTRtl1G75B4scxyNt6r/zbr+5fB7q1HI9o
lXuuUCIBCDkKKj1LgKdTWS+rRxnB7p7baTtU0jWrmsdaeQn0XJ1v/Andx+kvRdNL
0J+3+2vhch5sPrE4I+PElZ73ICG39vTXtEeA6Hwe9pzNuCOoJbX7w8UrN8tM1QYx
ZznryVYhE3sg71HSi25I4kBhX97PiB0qnHJUKxb6vU1UFddOjNjgDzN2EDAQ+/dr
THFRfJjtcDJ36E3/r6tIEpanK54Dtdog7bOpZ5kz3ZJB8IcGXDAt60iVMBC6KmMr
+IPlLP/7GfLFfCQXzVbLoAqVY25DrO77/RN+CgvMhB1uIDRC93A6YazpHVnUvRJN
cwHzYH/LNFW55qZptAc4ZI+G7XZCMxIUA6owgMmB/czIWNYFoSJSlyCxFYBBsbih
AoJENtExcIUquk+htb84S+N/AJEoEsgPShUtvkkG/WUkQWvZhZPCWyE1w+5JYRaD
P5IIkUfeTU9FBdEmjM8YrSUEh3NFdXWPk1PmC70sUhAm9ILHRqfhLLKd7AM64joi
IbDF8Wu2VKVtSadzk0KuODrSh5jVxSOtDVf10bnnrvVkTJeEUpRWVeBrKGkihTlQ
w66qBrv47PmnhSWvB/y6Ta3O0hvBboUqI6IErrN8gGOm3UGj1QyFmSPDE9W7Cbi9
NabYZlQydeoi6yPmvRqdi2288ODiG1vrJC7pH4fd9CLdBZhBnW8Ae4M5BEss8Md4
O+h3gAQd9Qsvrjqrx/ceGtvkaHvVM1WnF5WUbO3bH3+vzaHR/ga7VjMsLR8d+X5b
yUNaDtUiUmw28rf21B/F4FAH5cd26MF9d3PFSA1KcwUbH5mL6qT9ggKsR3t4dI7y
FGjmxR5jK9X0wn2R6b53f5jUOz5aG5y3/bEF/XEuMF80lH04RMoXHiDWQI5YB0cV
ND+UJJ4F3VkFdyGWIBrd9KAU0Ilm9TCtPJ9yddFRlzezsA8kQ4nI5MbNyJSvB7wn
KO539CL/cep12MdpY6FLmd4j+SujCpz54sbJ/CDwYcbhQqrKK9TuBacxESly2WUF
R3GmHkndclIyPJaEZEiE+G82owKTvx/AZhaPCHkLSw9lXzqSO2+WiRqDFi3ga6Gm
R4DiFePXs2oVddaxyi9ve0u1kl9viTkh9n9jAbjexxq9weyo/qZ0p4bJGOMxgX/C
IVJne07epqy4K4MVBPh0kttd0U6yYD5364Y3R6ObyVsF6X/6mRrk7E6rjtb6ICiM
tGaMht46pdJ+lbvY+Rab+dL8DLdx4qTm2yxP6Qh5wck+Z+sPZvro0yviLb44J+sR
Xfs9ZA24xNGIhm0qGHBfhoHhk9o4L4/w8eXEw8wiLIPj3YFE0Odl0nv6VUDH3dPg
pBVIvYY72Yf2KA1TTSduI9GXh/OQJN7BI59rSNlxiOj3/oRlHE/avPsmoUOF26sV
rNwiai995dsPNxNAqecMiDUivTYClPC6LInANhYp9+vxvYVHwwKENUyDNudJ7kwv
4zre6wjKO3AGzdLMBOq30+U+HdwTLVd6tRsUr5oTfu7tm9o5euGTap8Ay0vTKlyt
uDpG2vX4slOKG7zkTENdlBO+XAR7m27PJ3u68glqbxTdxaU+VGKmfMu/ghS/38Vi
qdTgP9oMRQRyywvHg1QHcZIUpdaygchJ6JudbIcvxYMWcXtc/yZm9gKDVoqY9/6E
pqgmDEarMt6mqJ9FXh9E7ebXbkNwAUw26f9uuCTTfzEONbFPC8S+mIu+VpZ7MEyA
5XucJGk/aeh+cVXLFpKw5djLWFf/7SJRCJuO7ce1gPQGhVO1LBgxDiwuOUEM7Xrz
5TGGs1enTTLJtwkeIKxkU68DylYVqBd1RGGMYSCYNwNsIDrrLhUkyd3n40W9wtnu
BW/QTKx3LfMAE8koxP+duSOtSCNXUhTT9Ub4Wylc1UXms9F8kRnqsdYzD4LgBnHK
E0VkXcWnygqzdV5m1eemvEkLY4tjFMiHrjgIARnGDO7QmWb4aVMi9BalaHg2aUja
NqqaX4FOMlUBxBXXX1zXRDuayW8CE2T1ikVELCcrMdZ32VcHyyYxpNfaNUcVX6+i
hu058x0XO/ewPriGBt0v5+YqdlzAIiC/6eccIvwzNNiV6EQN36H/H+vD4gTZqUwp
3LbqC9NFX1oWnovOTo1FgOb7FlD+n9jvVhFJcwqs/wXXVgz6o5NxlrBmz2eA0+Zq
g6FR8Kt+Gqut5PAgD3AYCt0/NbGZgdS6imZzSe3of9AsTkq7qHCXQwjvn7S+U4Sn
LPbkYPqZydQaY8zwIop2S8mui7wdQlvT5YSnta67rkyFgdo6hG65RUwM79MjgvuY
yZEQ6Fr2xVzxak2zqoqggc2vbJy5zH4F2bow1d2Q3hCMq36WSu4NaMV/eOblSHQ1
SVoucTYs/55xty2bvubggdE0bwgd20GPViHjsEU8cNg74ZBu5BvvBioi7n/JmBi6
86/CKwSrXstzFwDXpkGCDNc6XsqWuLYr2eatBFri7d2M7X7eqmXPDu5RgLe5uZdc
3LEBpraoni7oSKL3lxd3an2V+8QAbJXwwPvhvR+fJcWVkh+Al0a/47o5dwZyUit5
rx9Sq5fwFJsZpJU0Jxhhr0kGq+djJxEvRxKf4l7lkP2hDjXTxpB7WmKN9UPwVOvJ
UyFxtoqyESnpkrTDg3WiMcTFQNbv/qJRzrj56zVy9RnzRUIYjUb1eUTD2ToPsS6n
H+tXxk1yVs/7Gks8F6LY5s3Fh1G84tWS0Pke07Oms6jhhqe8WeFN3YVT4+gkfMSE
xB+K1su1lVGs2ThvDrxAf4bvCFpv8dijC8nHRrh/W6ppCqTxGhA7G6OLc6leQKO0
kCOhIJXOtg6dmLMf0j6/mz0JrjScrLShPOZ7yAmF5S6t/Wq6vz3YDWmiVwfi47m5
ogIwtzS1Y92IlggdOS1DnclNWF6vVpxrx+TVHmYCu+VWJYCQq6RCosCi59pJb0sX
LENI+pPzMVoXtAhER4bbfY4uittyASts1GlgLLvqQcDRGbdFo5G7u0IY3kLBpzej
EJ4aHlF3FC9Kb12RLN4OfX0dE+4FmUNUik6dwHyCf3GZdKjE2bSTNPqxiW0Jg4ph
buKmrw84EM2Zhjhh+SZuhHQYGf28jEnmCoUaa3hb6UTd9otAYq+qzJcENiRtRqjE
zt9QyRaKn7YMjuRZINxKUZpmkkJk1GYc/8noj4zTzBP8f/B6M2Jg7pkK8tGl6HxK
FUBQ1E/BA9qm9kCQ4oxCKc8ecwwCFZsBTYFysMYmVCvazr1x6e8kr+Hrzjdz7xuf
ri1/6JmxXqhjOf/p2pB8loeD8HdZBYWyq5yGOtMMStmgf0100GZThqGC1eS8Bcu/
3HHOqDEw+v77k1Auyqdmo+59fRouLLZ48NaBkC286O41UrClD7NKwB9FeRYQSAfL
fUCJ9y7NkJKAWO1VxY4czTKWI0AlEIuh+bcVY1Oa0GxDR4bXTNMHIb/rmauj6IO8
OJV7muhlar+v0kDjmTQW8jXfgJoif8DnXTwRc1qmOafUCjtcgNKZqNwTIAFuPIhA
ltYNxUsMuAUtW40RYmXRZGirc77XgUtpqHhfbd2SdNQOP19P8a+FMWknA+f8pT+b
7lslE3ILBF2cTcwxUydkb7lBh22rG42ggFIBGL/nEOu/IY1aRPzwMpWQ7DpHoiLz
cxoC/inITfFxGIlFQ7fSzfA25GQo3OIEe1+BYLweANGZhEBwwdYnJgtPlruX+Rnv
HIqk/33st/h/T4CGov9UC8Au6uTkqBlnzH/vVFGNmQCAHAfEitc/eVulHLxPZgD1
xfdRok5v8Hu7YSGOHxDUiUP+BvhNPWQPtbSV0uB3kmP7agFaPb+Vce+grfqJ+ej9
Vb//rfMdC2/cQdgzDUlwkjjwPKjUON9KcEk4FLDCm91tfCmXZRaNlKDwIGx7MCUD
vH1QoB5Zy1naXoHgG76sMYTokmGm8QRp9/3dtK3vrTns+djyqMvPBXA6t1wVjunM
4y/SZ1pbcBwBzDbJ8wfN0Q==
`protect END_PROTECTED
