`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IYsc3PCXxfzGYqgDqz3j8CwpRHDlhBobl/JpbqxiLGoQiTVDB1kmi1fdu96rzd2x
HXMHW9M+0Zpng7jFDJ0HomQQ2/CM59y6rFiVKO/8h2+nmFMgq95vvUf7/yPOt7OG
iNdQhk2ajxDVvoWX5QPwOAZ5tTLg29Ba5Q5ENVvzy/hNiDpyzoP7M3UuMNMDKOfC
mdqfXdrWLs9ZhNFqKaSQ/2pX48kwdgtdoKBApkRIVRoqmkd3X7mecN4qt5Oio/CW
y06ZDA3YquTpjCDqauPL3U+Q9KF1z7xLeBZnHv/FtNW2QebW6iNKXTYjKIoaDMj8
RcBfu2/uVp2FXcDnuLZC4ELr1//4x2h/prCXearVozQM6UzKWnOFvuECPbGm8RPZ
oz5Lxp0Rygj9kqMqK3sbe9JHfWEaMn36tmTWtOXAEZML2CyNJbSm1Uh+RupMO3AF
FmjZ5pFes+VnR5etaoavoIyJjbVTyNbu5UEnb5iYVGhn6l+q9TVI7amvyPpIiOns
zh2KEctDOH5xMts+Uwl5MWqgcpVsEvcbsJUMG0GPdIX0O2FP2cXGwpN9Tq7EbCaP
v5PIPgSKnqOWrouq0kRxNLaYbjdwcNlvgTISocVHht65BhiuDBvm5dUHTWWGK1qn
aMyOqlEQrQR1rQZqBR39zLH6nFLHC1moeIbwO5IqggniXtUeD3KJrExvH1EgAJA/
xB/xjm9m+ph88Wx1PKFprPPZc71Y7SbnBwZ02doFOFBUkbYag4d1b71KEfUhJ8AX
NAeqLchB5ySUAR6S2+Tg/McHJzE/llXAnXZF4IRD9lqHaupIy2e/BuvaxLbzPQAA
Ho1eMFbEYOv6InIQLxCun7AtRxHRTZbK00fH9mgi2J2DXildlzKUDbR6mpFkFWqC
tAlxnt1Ul4spxrz7dTuLH33xFEIIjXjyjdmhg4SOOr+P7+CnHcF4rnfbg6oIMpcp
`protect END_PROTECTED
