`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
naeHxLNf3d+KOga5nV1daU1vgR/nt6nLqFF7KcCJ5EpjalY6ahshUVBWuqpa5kVi
3T+d+nSx7YH8aGW3NSb5AAw1WkKQ5hAsssjjHdWKYgl4xp7kdRaeq8tSuOegxC2N
gFDryvbxKZgnW7ntr+5LZUp8hMw961aRpiwPMdlh6NIh0uMusRmQU8co98qv+rvV
4flY8r1OOsKPfgVwsNsDWb//ZbGBm/Cjk+rRrgy8iIgeGxzQHyy12dGVnHI4BILd
pm0pCv5zkjiHfApF7Qdcuamjj1OKQMeTVOrmQkARiscuQd8bijkptNQL908WRjea
umdC/iyJU72v1SVNDZ2BTWwp4QwnNBi8gjNqTY0qtjxljTv4vbLX+Y0MHmhN2D7R
ul/KKIha/46NcdFGZ0sNyURXePpj3O+OusyQhLiXzNRxVX0uuBILDy2YjidK5mP1
VSPL/p3EQQ7suIwqkbqCnUdEjSWtUWnjrJURUg4G9Bov6ltPBGFpcUmgY/U8mj5M
z6XodWSdsbAXGrCRUvdqYYbVEQ7OTJ927ZJJ57nbmBWLYWGetQK+jqOokmy9aqdX
I74pMmg0Jsmz803KX4BfzPHDTlgZ780L9pPvCnNetowrYt1hofBdEfM/o/zN4Hpm
0Vuaz54saIX8Blihg5Nn0jtHnbWYc4Qi7/tgnhTQoF1a8jYitdNo84448Ws0YHFq
96vtFUDHE0zK9Wqy51DK/1Yp463eiBsmaBVibFT671vgqZKgyVE+pF4xtWmruPoN
IN3XQU/+PkWbu+38FrncEynGdAETzB1bekucNxoVcwI8Lp/v2z6vfA3AOMRjrIrn
WUq9PanszmIAeoCFvj9XSPf7Rq+Y9q1X6zNWxg4gA40WdpCud6eyiuqXBNf79ZnN
VKUUxsLNwsNHupcHe6xn5yu9ksvdmSZ6yiWaEwAczK3SzdacSfpJTlLjjMWM2p/4
CIjk/3EbEGFq8UW1aB9nHJwARcM4SG4FT52OeYaGMeUsMupKx0sBQe4/1b87CZYX
qMtZ3Su/D7ROV9diMg5UZJoJODQYbi4vd+IufAwa7nX2RoTGe/HFnmszJZDRVFH/
rm5E0VMWaWfMr1wyCYB8mpyOL/jF3deLEiXFDXAkbnTpOLedQNwhzcu6twNtDTB0
wHMi8VuZLvqDHiowPVS0L0G3kC5vLdXf3Jr/zTIHq7AlOLRMjpTgC+DMdAiTo6N8
hsgoBS1ZF+zD84hwI1cRh1eOykHlEb+eyzFEDzM649fyz7qeIBCcgILugfJ9A0YR
t9/ubintrrOxzqzwocb96PBCmBM0N69vd18hvlKHVpdyDL9KhooOCwbJ776lfd+Q
ZJYFXlEi1Rrnbmccm++Hl2WNbwDxRJ7R10Rp/IVaVZAUX4Kuq8W1wk51ToAujuob
lUcFTGcqWCkiEcuJXWxTcXh7Inka0EmNTfHJJBlhHWgioDZZuttmh1P5+4Y88AuP
mWbDupTSxwDzgmq8w+Jb64bNU+GiDJUUrjXYVaDRcFKC8HS97v3xN9x0WgwSneGN
/tIiQLCqH4QsKldYo4Wsk0uY80YQOKKUd/G42cfmpE22zEnzA/bOwUTg+OIXbI/4
PbTYmscfRJUYHtaMb1IwqSXV76Li5EV9ZK/TWCaQz3crHvJkRx5ey/HY9cV8nmT/
t5pGd446O0gkHOABHFcib9EjdH4v/Ug1r7OMjuv7eAsYQVKQXkT/KMxiQ22fceA8
tf+vVEL2387VfJ7dkOFLOuw/EVwaILzGWj7p8y9rh6cVACMDoFnyF/FGAhsYfV3w
tzA9x8xHov67b0ECe0WIllhpyzK/2ZgXFBYYXFdafJpIDhW/U8C5j0zpegyEPmuS
`protect END_PROTECTED
