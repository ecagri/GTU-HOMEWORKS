`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cj83j/Q1IPnDZ3nC8xio3iBADT79IrLN4VCZiKOxqhMIV7JwGE8SgbRCj7jPGeOo
5bD4XljxSC0bHtCMHauxA2y5/C/PO4oHOfG1F8NO4SRQXrdPH2tL1whO70G0Jr0l
nc+A8iwht6G2uKDVe1Om1su2FTVN2N4x5Jzs+LDWJbwTb7e27htTOFR1rTgiOT2x
3qKh4scXJesA0dG6MOx+oNH47fkd3hhrqZUy0LRO34abtBKLLp9nktXmZb47HyiP
p8Fs9dTdHHJvSdOU5LRpVpU/bjUkvyuvMb81rgZCGz1HE2SJllWtay2qhIEol82x
0Mp/SmB8dhSbjnv2Tqwuyzx7S86qFxj4NRak8y1Jltwc2A3pWO3noAtIbrDIhIHI
AKRn4xDCrKddh+SvB2mkie6bXtB370blDZPAbKC3XE9qy+wgBua0X3Ql6FE7YTYP
Sndh7e37u6s0fI46xfMvNd4nz4Xm7CodMthE85Jgn0NB6+NKXd/tK/OuHTmO/zSo
GcTBNCTP+rlJCU/w6FiejtBy4edA1B9KVOEfpZNflvC/Ckg2WbdXgy10a9GCsteu
1boynV8WNKX0e7CUEU0IbE0KJs3NHU+FppIpnN6anB6mr+1cqvGjqKAW+pbKCWSG
LO6PkD2f2u8/Vozq1AEaSd2fYsBxW68qT0gHyo8H66UYNZOvjkXd8VuNvn34pMuY
yuxoF/jM2oIZe2qMpFncdEeIyfYmUoYtm6AYtCpb3s+6U9uOnSvHQHbf1EupfIkX
Qy6kTHjBzhIEXU44OjbXQK4KJu6o4HcjUFTCpSbGLCP8SacsneNb6Kh2jOkytAa3
nwYoXtLlkr62wJIlRcyRDW8+PqgsDZQxo6d9Ziq/f7Au/D/hm8jID4ESPAhZ4CqG
7zJnc2IKrTVC+4UBb9lQfQWyMhJw1vjpCDo8RSUYjpMx8+4CD2GfVMz2+0Q0//WG
+ylpElfB4tI24+Wr9zgkuTrl+CWmobi1M4wUHSk75+Tzut7yzjid1L1888oqV/uf
9H6ZLysjByqvdNQ3xoVXMh4l4eRhyxtCR1fFYAEnlZUWqvLg4ru+DSTMDDhk7tfx
xN9zSd/KkbbAQdrl5lCNXo7FzNyQE+dwc4kzUJwF4qNF/7t1mu6g7qGYzuTvQPuV
pW0d8IBncP28VxmMnXayyv/+MF8G0KXxnNpRaOacuP3F+RB+oY3V5afHzMmJhg/M
ltJNdm0EKjqsaFBgD9Odk+re27c1thfmDylKH93SXEFR31CLUiDbFMaEQj4q3vD5
V1WPdn4vkMtLdpckugFd7HteXLUnTPAv9ji9d0e7wH47V409xHnazOeN7MMRarC3
UJX82OIRMQX45PjOurqrwvVqx2AuturUs0x6lIaHrnGueAAsYx0g7BuNohKjHm84
sJaC392e9m61d4XxAf8OLSclTkMdTyxZwBdIZaOztrGIKrlaMdYRvKbvZOLCVcwo
qr8AnyAHGxSEGOjR/7BK9SyutHxbhBAEeseUUKRLnrjv/f7eLbm29SchBRSkj6aM
Crbdv3y5knMOAq0ahe8pLZTt59+prMUT455zAY7MVkr5biSvWV2/zHLTVLqPfiqa
H1PS0oif/Y38k0CwqdjUhpkBMN6mGd+0cSbNQuPfMQKS13UweenbOYfmFEIx62La
1IfBf/Hw1rZJ3aztpk/8Uh4ZZRDXKIfb0sITqRNouk78oB33sD8aZtEWACSiyeh/
ieJLiNu7m5LhLJP8sTvuDJNXWf95G3xSAIfk5MLJdIkQMFyCIjpKMkM+pxJ83Lmw
fSLEQuKGlD18eHK2jfzv6/PYo7kRlxlCLFQ8wmP/P8RZoMJbL2lZkVRGFzLzRitU
yWpepuCrwbBQlaNYEAJVhie06XQF/WLkRdJFJgflL50OnLTdSEacPcPrMzMqUOZe
6YhRQBTcusGi6LkdvE058N5ZzrRKbm1vYMt3VQsnByYeqLzsC1v0vh8RrA2I0pDj
c4b5urAdzZsROaav96XaG6Yor7JOvEI8TXChh3sW/2MS7YaRGT7ucn5DcOu6fhJg
1hmbDrsI/63HUEIngtICm+DdmCwUcMJz7ZIb9aP9QEITkfdw8cbZis8Ry4u2NOGY
FT9ZIGtGTkYWZdmYoZnLy3DhMcn3cVou2yOmUz/Dd8rxxImIJ4DIAacnRAUoE6Bt
s1ur5NqoTswU4E9/daM+RUH3srxhkqjW20CNVv3arFNpt+K7RFtWCj/TW2tcu3OT
u4D3mwY4DpuClVHbvM/xTek+L3H/tJN/OaHUohISW7dyI7OE/H1n1eErt9ZVoqbK
qlJZywgbV3cUBXFF+gYQl5luizDwB47Gjd4/4XqqE/Bp/Cqaa9G3cJBARSul1fJ2
pyxdN+J5zc61A+gYWusw5TOX6YcdTu14iDTAEn7kJ4NVTNHEwNmCyHxa3wWjFCiS
K0PTV7HH5hSyHYCsxXk/T819xWmWkUMUQEXN+X/uYT27iasKVTUGpMsUQIM9n43N
BaDvxg1K2ZqsaTU9jjGu91SakW1UN1Sy6fMtOhPaaOQgtm43fs5U6Vsglz7mWuGQ
GP4g5Kx4MJh0bPwZgocvA7EdXCEGzfwNAJqcePwbnQWIDoIRMCOCy7LoxV788Swf
lss3hwDTJtTzHJjxM3cYPFygkINfoXgYLyG0kngGcs5T3b5cufOmZr1MLOISo26G
yM2iSEMEA2Xqp/E5uJ7wx9jBdM87juM80hEC77P4+L45s/oRV19haQYnxHVTvO3c
hJe9rW8iwjBMkytcfxgxrDIMUxY4RLLEiZ54qVQTQFEyssZDEys8iFIJ7053HKxt
r70WNxZ7pc2CkuIuM2cvDThG0KKo4zy5Kcec0JRKhruUjxi5z5H+t90kfl/I759o
1591wV24gR1EXHFSChPDDnpRYYjdvbIQDzT6NxPIGxIfX2Wp2mYbfxviC/C3RAN2
3DPHsVrbfqVDWPOqW4EFNNQVpFmZCbH2mQkHxp6PyPRLvoRuiOSNHIyQoL3fHBYh
IilPYSrGG42ne0L8VY67iWhml5+9W1E+id5z2AHQ/BDgifEZ/7LqCr4g1uSXhQwy
wkYwcjHvPkWuNK1BVFbl8MOkJ3zcgMJoDAqiX/ClVRUB7MdmhrIJ5PH4h2Aq4ob7
4OaKxfgHAvikp0L1NxHV+e/GzARk3T2VN8K6pWpdp0IUw/2Lb4w29l5dQm+yLzPC
sBMwqf7v0EjQNx/IyZvl4eL/r9elFSGEbTQG3Q6tUbu54bcYfWS8xA5sdlFWNSmS
LNg9gAA39ejs1bcQ3oZi31Eclv8ZxwWnyuuSRNFJUP3YI+b2dwCYpUgJfb9bmzSs
hp1J+dhWkGXJzOTmqwaZMkoRpORV9mco8ayQCHWHDkgg7UWXmd/Tcc+tiMZYfNF9
R4fsudQSP6Q39SNy1t7V2qt+lT2Xir7RlMwVZ15lqjH0wCeHgnRfykhP5VWPk4T0
R6y0UaDr+Rjig6hUw2NZpzRSnuFcJHlFgAUZootYMLDGc1Ez2RutpiC1QToJM8DU
Irxw/rDfJwV5jxRIeAq2N5iLWpg7EzIMLDw2B6XCAgkNPBPktG4F97gNiklBwO7e
hk2nTRBXYtvBoVuyRYMKto9wVV72sAZoOcWRVJHqNhmlgmsXfHceAp/RYCL8niSw
QPUNAs1kVsW+TaOICAw4D5U//ph8z/6ot4wIv37iCMfQxeHA7MbNlm0HdgToa1b9
8JDjk9WVSk3Tp519mMllAxl7AXZOH/snB+0BicHHpENPayCSQV/6Bbaa9Km1tsQL
1TcBuyO+UgWIHVrbuGq6hDhtubvu0dg1VhUDWu/ycjQ99X24Cl19mxZtF57NHYKK
u0QlfGG8lkqMNHiX5rpCm1GgWBPLZMVsd637l5cOw6790UIM7SbqxihthWPLZPXu
VJ4Lzx4nZEHGNOsWB6WohHcXeql+gY/Ra6UAAyoxpkivyBlxcKwQMuy8avF1uj2P
jx9h0X+kSBb1u5fHltlpPFVK2JfBt+Bxu98+CR+VHmvbR/tzgwk3Z1KIoB2+Qz9q
PWcpixpuFxcZTGk/ySTDNQeb6uemZ39zLAskDnTCeuUvC5sSSsjgXsz9BR48ig+T
ZP0b5V2aVMx87XohSE7VaGT26OUqDTbM2XNkUaKOJ4fwXNqGS4E6wr9KCyJfB61O
qrTfUcOdVmzLmpKgcY/pagR5d6R0CmiLM7hrju1slKjvC3WyivX/PlphPVF344Zs
wSSbGsswZE/q1sAyDALL8AZwmazgjZ4RdJlNfzlXQ1QggAs6el8goVB03xuquD6a
v3I60u+B5Y01DoTkXZySpRXi1yYQpQVKjTAFE6btNgnjSsvkw/WOmLfc4bomPCd0
/JP58GZ13W6jhFzYN3rhXlU4XlgSScHzGvLmM3oxRjAgabBNqP0ZyDS8yg6gsGRu
ouYNJ3PKnH57qomO/K5UeKyIhQUn+ju5FsuKfSxiw2PXjV68YogX9+bnZQW9eEuN
zGOEuHIvObQl3tk0MbCzVGa0ngzmHDWTGgNPZy5b4SLCbMwph9r/SY+tqFtsKC6I
m9Q9tFi+fYjuOe5RHxHaaIHlP3vcqniO/nX+O33SKL6+lgLIYmaMWRo5pwxohaap
cUfnOg6mrljcNS/aAbMj7y6iwvmFmcDdHUjAHi/2uGMgPWiK5ukzp/RxC8uYKapH
lE+5xjF0O+GqhKAk+RFTHC1aGt3wIybUtc+ueiO2GY8WQz8TqJPibVRR1fRxAcym
4isep3IYpqX22y0vIoVgeLBaEecCxNVpybWJyzOeK+Yq6wwmBry/jhgBkyxX5QVC
qtFkwKtUo1COVZ5kNyHb8lWdxxbQ9Bnrvz1c3lfrl7KJBnub0JJTld5MFKgd1FxS
pJt+jX44NnVEf8MpgUKcABq26bcOKjy7zfXv0XJ/yb/FYr4GOtuwAI6uwo+G0jIC
MN7hnVsrHRT1Rg8Q9TDxCGoiafCP8FjlZ0VxzV4BHKTav3pxPNL6OJrvkDW+JKhS
7mqivrc0wj/6Uc9ceaqKB0E8yhb0Ra7InllNHbpzGZQ+7M7rK5Tbe+P+TzfRa16f
qZDE9pxbHwoUtAASOKHjVBYspJ6KO2XedhuO2fUqHv5fum1fdxe4iJu+O9dFHaBn
9neLwzi0RjKmUh4mY/qnBbkRpm4kHPAQ/ARvxeBe+FTNWmDAyvcftcD9FQo/l0Jc
ByzJ0VLMoEB8OPK0ueWUK2x6QAFOilAojbA/dCN0e1EK2oFGSQhbh49nYCTXG2MK
eR7WMhHor7fv/pLwpM6fePfTn/s4WlKc7KNfnJ6sGDma39AqP/wIJmAq/+u/KFZN
i/bmNcWH+d1rXGQ1VW0/pnCUOxklX34RaMuJyg3Pji3WaanpQdSnDCeTsoP9MaZB
Io6m12ovqqkhSi8Cxh+rcy5nqyCghTMJFpdT8U8limVEQo+FtcDHbTxgpMOvkTZ1
u762KOM15eQhX+3sR5nidM7cEBhOYahP87wbl2V1kHoUqpUvXKN0wTC7i1t2kRE3
G5KCtzD02MWgQvDce3uZHFPUxRNlqkN+RXfUxPj+mPrUIdQX9MKF8n2Ky1xQAlPI
wRtvJo85L+kjaF2x089LIW1ZNSHzbi6ZOs6lkbTJOk4WAp3CZSnxZ2Tc140sPfBq
i4aEcRpz11H4QfLOQ8nhlJZmkqaXBxxy6z+u04WW3Q3Qmv27qUjsOyQAWsbM7JD5
ffyORI3RVc+9EPw/1EwDrFE8DdC7Uil2x/MUGcUpKClRHQeQkEIKmPBtdqBZWPFk
o5fCGiVEb18S4RjqvWN2P/F2bEJkphdksn7707ElW32mk7yCboV/GCEJK9bkIM3A
TlSPAYeJNoY+0bUuwINwDqlQu/ks6EnWYZTAqLycT4oJBXDariQdKlltN5Ddwt1Z
UFxnSxEs7VU5uBtukDTRSnI6pwWnrxFoYy6NgLehPl/QiatNHgwwvHRZSiKNp2YL
ARsI9DqkPXm9GNdDP5r6G5t+PlKF98bDKbK1AXfUys/Lax/Z7K3ro9izjRdzzpjY
CIHN2AiI3ksZ6LTFV/crn8P5GWAhUfTDUNLPe7ASDuLFvMvpTCCat5R5EOEl219a
Dm2qIT04a+RuJj073NcBOTNu5913QdHrAi7Okb/zodGhiwK0k2WDVfjgxxihsFuy
WFLRKeDvUMCW1b2zplzs/Xb3/MT5yT2dIscCd5+i3idpSJ7/6Nytx7bXVt+vCAZH
yKzEYRyxicSJM1Q1BChnwVj0E2MRd+KF3f2vMsLlopWeSKgkD+KD2xZXanj9P5MD
penAOKbds/J+GV1XBnvfgiFISYsGeQVmK+ZqDjijus0lb7VJ76EGm1rEMgxbQSw1
c8Tx/QoEBErDDPYY9YznXfr09A+yibt/gY/TMKpxLj8mMtnUR4W611bk9JLDZaRL
inkRiZ0LKxYEuqtE9qLdnWBi8nVR70wnJUE+y+gNLa6IE8DkO8iolMopbAlqvVwd
iJQ0a89HrBeVIzORrjs/MbdWso+QLVY5E8FQ6Ky0FWILI8IazrVk/Gz1RUhK3ymB
zwo0RVqULjVMeuyAiwcGabFg+rMjzttyW3juxWQQtM9rTBgCeMOXSrUWEhKU2gEm
Kl7Cnsubb//AmqciLB+WALpWFJ/nJW3mOATnBDLvOiZ5kl4CIcrmKHDaTJcELRR0
ZUi99y9IpiVfRiV6UlD7ioasRKTM0PWH7DFpyh7wImkyBL50DBK2ZCBkBxomkzO0
oJsXD+XggRd+EJsXIYfVs1N51c4F7QrGnbfIImkFVOsew89/Jg5/NEDDTtx/us2q
T8408Uw00joWajybC6HhhjOabi0tW9gZo6aj/kpyfF6xWbjormyVewq2VyeKD9y2
cngr9snLbzMyB/5I1ioYwgewsxvwJWAjXRlLc7BqMv+2asJGOPpa2UIIfzBgUEPK
ZUr23383XJDy4vILbsrbyKlgRpZj0N/t20F8yjY7cH6Hb5aWNm0bO1TMA6OLO3UH
+UsZ2trLaXvTbiLQd5OominbibK9X4HC1eQDKi0tSPYbd3qhbUiEnJuXBfZg3MVM
oLW969S94a9h3CUcgyY2iY9BPknbTTAGA77AvwtAc2XtOmIjbZ5Ir7xr2m8TUji/
FTH5Lr77eucoWqAPcoPE66FkHzBGaLcyuCASSNCgiBt+bSExT6DM/pPbuo0E0O01
63lFxr1wblW+n2W9+tKfsEgFMz+xJKlYQRnGuWIndovf4/JuRTqQz6qhuNumwQEF
0CN14PZNnVpP7MybdaHg77k4IriWNG3G6LLY/Pwrvyawnki9+WlKAEw61q3VRTTl
mjwjTUHDFmSSgS7wmIMRVlpEso+HtYiwS6+6SVZmSBOf9zjek+mzjz8lW5h0vCZd
Uv/ugpZtyjUyMEYeYueFchaWGgfa4VdqKin/x2JgP31Px2HuNQhfbfftEYiMW3gT
YUDARxnsX8wV+7PZlZgf3fTWhUzAIg0/zU8OAck7Y4/7syxOt4PKhN7+5cCXcIv2
QWB4xgfmw3gizsaYhurjeBe/h9V7NBm0jm/CZ6OUTIRXLpjfQkQR7YEr+oUKaKCv
5y0DdJNVf+nXDswJs8VekT8lfu+5HGkAvbNlBrc2tJi4RXuKrOnQtdNWclLOhYBY
ZUur3cXBruAqB6hlCowgU6mWCSB/Y6k55rCReqJYz0I2ZY9RUT9az3MPDnoxV3YF
6D/brIZN/EWb5ayKqupf+U8p7Q5aCZIAnDH480UJb9LuuY9ZJ76L9R0gI26iF0XG
/UUiYsiWnnZu1BRoQmlYXvi04dH+ZehgHoA43EqDFBvRCFJfpVkrJXEgYds0nsEp
k7Ey46ZRTaBm8eTnvvV2WWskmi3Mysxzjq78ryretObYf3wG2AjHZdOQ/fx+hwXP
WwNR5PeC9zhLvEyYJJmxTWRRjrNRMa5SEhs2nbdrh6yX9cbyB6BZSk4NmgQaWcg4
0GnW9YPS7/Ntb6ZcaRysrBQm2gGr4it8y7yabD6r3c5YebJgkIN375gpIib39O8a
TtFo90Cf37zaLTug4AtEsI8P6zCBsfcbzHAELbUH8tW6UsufDbB+HgtpxjeBahrf
D6mmnvpxQ13ts8bA5XS9uRbC1scZSh66gzfjXSN4eEml5H5juv1naEh114G0jPjv
WLiEe1N469/DZaJK//bNioP8n93oUijhxBUzyqOujl2VcC4FuLXh/lh5ytUx8s9/
AJ1vVjQ/YcFFX7EaG43Lmpt+wtZZeVHXOO+t0PWmCivEj7KCcMl4QsiLUuBwMxyr
MKMCjz7PIG4UPw99i+0z1VwYx2Id0B2pWCiyqKMcj06WbGsesojzwyI5Zr6lpfek
vqk3II+0kP3X96xZmGoqxBT8xS7+yghtyneWNAYc55ToVTtuH9woakxwKtV8HENC
a+vnNBQXEZODotgMCfMEjjbecRg1mXqvjvDvCMp3fM48g4eUpsw4JMH8t8S0UbBt
pn0IcoNicRDbDTLUk+HEwJ3tJur9VeK7IO25VpsUDVhwZtNDq1JRLdpEnk/oq3DL
hfdVlFTc4sb19Dn9qgg2PPC62iibmk+2S4SLGPvEdc3Iz1IqR+96BlUXhfXF1URr
xWIOqPyFjnbE466GKekadool/v4O8gACM7AWw4Wm9blxNv5mp6oDS8zdUf8sZpfX
tCgDRky26A94QvYLWAV8FV+AnBrrWPmAP5Olds+uMtEFhvv+CIh7QnX/DQo9iVHB
/d8c55mO+pddJcnoRv5Y9h+Hs4y9M7VQcTsNLQlzMDRFgtmOyq20JT+rJziF8pLP
ENacNo9cCrYrezmzugUpotlpQkaiH01P3PirapriCJsg5j9limFCVv/JTOA8a2+F
CGiv7cqwNR5DT/eBNPPkcmIc0FgD43qrH/Hzr0tpru6JSWsHWl5bTiOeybm920J8
/mfX/xsxNLRgw+r8XCESmoVRfGDQacH5oWoLeghS+3HYQKn6RwHO3gLBv8iESBdo
nmXCBqTDvCUN9c6NupP8ZU1UTENNkxj+00qwKjHZf+Eg5tXRdcj+3tOORBNXkQ1B
pEzw0bMqyoKxolyST0BTUB6xgWvn3H4rwEFKCVQPwmDqebfGeqVDDBAXc5n1dQbP
xPZZoss1vQkS+fgScp5Hf6QaGHoMMpsG6FyStw7bOJYA4Z9wz9lvUU8wXaW5DhZ3
DK8XEYUhwHH/vFgwSPCnOkUpSQmYNK8gwEu1HnMwjt5ROOccNuU/HXiQwsHM3QCU
IsvOlCGz8P7gqAEtxm98ID1GXF0IBzpIeWZh4eloyNpZn3kMsUOWKBpGjuaE9UHN
EQctJrg9DlLX1WrBVlu9yqeb/y/FAwT27j0t2AOp5QqGnhoZDf0rWCiKYItEnrYC
rJsoAs5gBHE/qi8liANeRJfN6TzObcY+yJtfYObxJkrGOkHkDxPvGMyZZLPv31z5
plTEeGQikYW5QHfbayMcg5+2s6mv1YDob+aS57u0B/NStljNHEglE9tFVvXyXVV9
yQegExh/YxQ2HrzW9oEymNB0o6I/LFvQYSzhBh109iijQTk0uulHLWk9cBElngh3
sOmWTLgbf6sgtPige7XAOUAv/Ox0s6hzi4BV+w1Np1r70DRJAr+nQguJejCzP7kV
Gj9ZqLY2oWrI0Wu2KfO/SvJzGIHHycPmKbhrLu6O+HE7rJpC1CL3d5do2tKiTUll
eT9oEvWunC40nMneV9PcbrZQpKtgSWtlwPFK2dmXJJmlmaUO667z6bg9LlRPxDI5
8YtgXtG4miIFJBj1RHhvHbLgtTWXQuByuFds3a3LdWeiWJcLdmJWxwBJmbxTcMXa
D2QsfS1H0ldiVe/KfZSKwQM3uQireP+mcSbvJG+9KJ5vcUs38UNT9pmFFFrps2ms
iqn7MN3NYZ2epXCwN93Gi5d1a3N9EjpIkrOssgv0JlC4SOHY0W9qYwAY+0Tfm2Df
D7FpHVflgp8pZcF6kmr4tu9dB8ljkcOggKy7O6OlVP7xddU6JJTrnvqtZ8JAW/tG
ybjZp5H0y3nx8L1YUfhQ5cfTHYdWz56PbS5eAIFWUZ+EtFoz2YlSJbVm9hY6fKGM
82Ack1+RA1qp/xlrJxejZW5mQf5QuiQ1S0UL+M68VkNOBrGAnlRPQICaQRHHVEFX
jThBFFG50Wpir49PLLlNwd7m1i9rW+D2+xIyav0TgnxxsaW+6ge4fHl6VvpGZfLU
vr5VboFLzge14+TqqkMJ/Lb30L1yvVGu0c8UkyY2QXhSadDB5ryu6kftYqAC/47X
wBKIonF9BM4yeeG8B2U6dmSgC5+NhrTN1LgDEToh5FVE9za/B1ratjabJ18RXr19
1EHK3EKK6Ag2Wj4KcGT/cr61HgT9KFXTRvdSRzb/dUZxijb5WpjhQdP33ivRJ20L
kCxiqO1Qz0iN4uM7+GuGqpFfbGgtQYLXtIXxtT7ApwLe8zAoSo6rYbytoGHg3NQr
JNecPPxgtxIkii9IGT0Tec2KU1SFmgkeqJjccBK2lYkCUr1nxXZmYfheXYsXEA4t
zPpKNgV5yGx7d/vwB1wQmqIy1dXalxYQaDVfI0znrfbaYPzSzPbBGOhvboeE72QF
UjyoljhyoWKWkTZjMGcNedCzEapoVWKhtHxC5o1/mCiJKTtc2nU+zXVy3a2LeZNR
7Zn37MAOErMHRZROEDbkpqXW1RnW/W7Ay/8dM5NNlwdNJVNK4g5IDovIGvrVS7Py
/TDvmYKt9rNtAJCUrRWnx5Sxz4qKaHKqy0X9dbi7+RS7FEz/zDA+0SAlKAR5FFZa
tgNDGzfup3Je5qsCQvFtF6IjNLL83GROnN3osXDA5x54ksquMe0+DxbA+PGMqmZM
v43XtWtAGSSGRVHaWitboBzCrpFGE2cvK/GoDoCd6A3pwrbOZrG3c0SlkoLamg7Z
3WeYZwd/xzfMwgpumOxshPyKp38cYqKsaTdvxOfx9Dva7zTI941ypIOwAueQj/nq
MQxJqh/znLkcsxYpS1c2cgwhYxuuUfcSHUOQl47dbUjsjAVEKTvWU55dD1zBFw4C
d8iDy7K+ymMuIq6uTaEcDACu5vHvRjgYc6dOGZLNLIfCUAkSbBuUOKYFG3Jb5Ocy
VAHgliLUXVe/qJg8lMbS1yTU+3+w2jQy1CvSggE5f7lrolB4EhowwdVedHYj0puy
0e6CQmBSlZPxBbgFIYuHiHnpv1CVHWYkmCzAvWfc21GaSpxgxJmz6rBwdq2hOMZ5
bDHwdq3oAeobt7KY7EOQO4OeH15sAypkr8XZRGZ/QJxFWCLUARgOmRiuaxT10HFx
BubSw3WE4+xLVKgcHBuagA==
`protect END_PROTECTED
