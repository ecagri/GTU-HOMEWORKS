`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9/AnaHYLDfNHP3l52I9MhTtYd6aoBIPx004hMY4mvGAtZ2g1ocH9Rz2P8fTEg0B2
Xlx7EsFop92+vuz0v0CWqvn2pkIqkmEd1I3IoSaqN5ekzbaCvps0Jq26zmA3rS0K
37us3qV1lpO6a1I3t+WeRXRszQxFImSrfSdbaRcTpk4WfSH/wvj3+V79g68U4wZ6
J4jcynfNRyB3XoBIA/IC2tiQiNu/xez9PsLTbuc7MoSOQNWKtrqLXj1NIJd2pwnf
qwy/ITL5jHolz9gwKWV2gpZrn614A7Extry/aPsDCIiq18zOoRq6YU7M3iAMPn1i
pB39PbrMUMqwOrHujPaCVP6/Es8+3P7vFzHvzBsZFbNYnMKUKFGvbdg9qyzZtkK+
yCtBjrTIv5gzkUjBzfO4Fn1b9mV8PSvHPrGJblq8a9mdFNIqPLxpxvpBmHlGLnT6
9iUURoEkM81Z5RpjRq5dC/hYhWlaIZZXLbJQd69lBXkXAADtkCkl2iAXVMVS+L1f
313IAKx0EW8Waiuejbg3oy/eEI/lX175x1riIw6nzDrVEGnk1spyUTF+nOFMwHlE
lYQDPADEXYIjAy+6TRXLfEDnalUtO10SVpAm74cf5b3bU1a7IcS66DYJtAuGZWMV
JG5nlMRPg3Wyy2Glj41GjSLmz+8FZDqjVB62neiU5lpH5gwQzLmu6344ZUMVw8N8
nVDqnVF4Rs6gk+Die9LbjLIloEnTd6HzVNCWKUHC0+sYimhsToqyF5iqQ7tqO9bT
cQgWmz5dWnJYnJ5fzfgDTuTlZUBQJylkWUpLjCu4zPBpNqbNlihnw8cBPSfBSuXO
t2QdeAyfZrCM7hx4A7f2IT2FEg2FP46h+F9UdcQTju69OvBRwjuRRpupzUIGb7bA
SS7iWTcuj8b4OCZBt1ZiRMWjLw08FPblXA8isPvKJpAOt5sA1cplFPhC/rNb5e9J
f2mkXsuvVrqoA+uaVYdHnq8oK3DD9i1lCQ+B75bOzD6szknMlvE85q+G9eDSIh3l
dltUyqQ8D/mdHuflIAUM0iEaN2FCHRNfd/1qpEFmArs9kAS5ob7kItGQufS7CdAf
aFW+0hIlavyFv3jM7R0nZNFpODARYqt450IE5+2slEpyvdGMdX4tMZE/d//ZWD61
gV0/TMO8/lbLP6ILKaZuJ0Ym/XOoEmJxrNW1uZRUCwFpRA/O+0avoB4WEcPZhOO0
px/i6oT8rROGO66AbLCN2aIt7n8bkFMOyR2fcPQzqoMPs3Zn2Wd/PwBz4i6IagYi
mlB0nMAzJaG/ZRa5Kzos5NHB2dHkL1kkQzloENasCmFDne9Nxmo+6R3E5Rchp3mt
ZOipIHEouj4vclp7iSgB92+jRnlY/D9GJQpA3Lql7b00d9M6jIbXJnrrapJTz0Fx
HKpNbbKdoh5WTHcg2r8YBpD1oM2Us4Yrw1XxscqbzsZJeWQQCWglwrOYRlXCBixq
psnZEK8zSOy4LbUV1y5nlsMdEavlKdryPOGvCV4mCG7v5zGM9lcBxZMVlSc18VaG
XdWy+9sYmbTK1xb+M+F1VguBKR0ucfhzZGacFkLULPy/Xav6XqXsS8c7VfVv3pk7
oVY8Hi9Jp/L0QTclSyHNOzNH2m0+cZhP0WO523PzTko/aysd//D/0ebySo7tIYXo
j7dtiq9WrEhtKa0pInGqxmqvMBCNgij8wkRZiLbgolipVT/ncaDHVfiPvF52GIWy
6kLGDmi2ZdPNosON4frXGBTsDi+1+na3kyixGmZOvFxeytgPfvyXnk8Gj+XPJKVO
yVsbneLWdijyDZWQCWDnuJxRmzJ9HE7WDsvHYRcvZtFdKxVN40vEs1ws7Am3BqIY
xiGeaO+W7O5jz9c9+NdEHKhkW8piqWAt7z59ECQ5BZ+2JI0mVUXEz3geM118zEtf
bsUxVwf0LokggiWs1wVUYzkuBWEOpF97aG8V+wVhMbjwwfKwnMpLo8wfwBnRYuvD
mflrFwWLcEzjMptI1Rxb6A+HZjNFcqsIergNfKq2XHbiIQDGDzqAIDcLcYlXdLg2
TB1nNlcLHk8oA35GCb0v4ptyUu1Jiq6Qr8Q7kfnCn4lvHYrrraqGRCQ4RTtMVaLD
nZFZY56xee88j5HqfnlczfygNivUP9qPcIn2OuwEyEhYklAZv4OCYU0tZgVvxSLk
SNHxCAfs9DBSpvCW+XQ/rC8nTw8ZSpZclu9EPfZBWC8Zh8YMlt11PQwM5w4O/AQ8
m/8BsRHcoqsNOsO7WIISMk/G/CtbqlaqUpN1YZ3/4jVZLglhNRmgPI0AUYbmUl77
DyGAQrNHSqsmE8A1oCJ6trkZ6ofTWSsqzdg0jNX/g6o5RTCcTUmZQAKTZFCbUhLP
+tM5bF1PWi2DZGLv9qLODdksMykPndL1V8dExdUEYCHYV7iU7+jStCiwDxsImcwg
qnlrYw8kMNTO4bN+YG2KQqK5p0bLzgFQOVvmVZaHEi/WTzHjSF6vwldULNrOGsZK
+joMqPiaSKOeODRYUb7roPkt+yn1MjaD69bF4KwN1rm/3ykNSyUYpYYIHD28rpmS
yhlypV2D9v8TV+DUnWyi3/QRFrBNDSSdkq0O3mZY5ZvVypSKuIprFCEaZVLMbxLh
mkW3kT3c0p9CFzHdtsarmdFWOlGeRaBpzwR4Bg8KPgPrWd1ZT01tePESMX3fzL2t
gXUBruqoKEULybpmhP1o9g85Uh0Ds9PIMYcbYlwSqeeJ5/fkWDbC1UM5SkWqHy5S
PyvQ4GX/jIcTEwfZUz8dmi6o9pvpxhGBA2r8WSZC/dh0KybvpfUFNxkNRkWEPweO
0XoxicG2VsZqcP8oFfmSL9SkkyfI9dYU0quFCN5OmiFe4UwrZmAnmTwzPJ0Iugw5
prFs34jWyGfbTdvHjTR8rQ/XtSFbUqf/j979IrAXF9ZbPa9xXCP3TxwGsTGsB90q
5kgKcbTyTj2LyOBUqddaEAJU3zycYZCwrP5EwxiICfRIhqEqqsCHS/aGJPMlKyzK
zYSihI7VuJRBdteZasRe/APTsdbSLezUD/Ow266e/OxDF+OGyQB3WInBro/jjrYa
4XuYnLbBHC7aMFQiIusc6qLvNWY5xpQAA8eKq2S2EK6XKgm1KxgWgeaG7KJY2wU9
BmqpLEB15qkJRtMwVPqTL0v/5kikQlMmZTth+/RhcUOU2pTXK4X9KdPj215dQJYh
B6Uqg4+pRVSAw0/UdUSQphlcf17LdzIFkvKpllHnwaakXz9pii6bpEdIlRKEiMhC
qChB2Ol64VZz0kxXkESPuK8Ilwh8SCQPbGHFWcKDaORsAJhcC6gULy0qAYWQxWxY
13NVEk5NJLCkgJ67qgA45L3Va4oFE9Vn78rEqBwPz5AdrI/grVgbvxCE53NQKnGh
IqwuY8DTkeUEbzLAFLb0MtaedyYq7Epi7kVZO+zKfT4eKzeh7ao92u525C5te/PJ
8WRfDqRwOT4360iUv5emd+GFw5xSP/cikdlNwllhTQD7D7aqVExpaJNWWMaEvhCd
LxJtD1i7cqfSEKZU5v6bRvCR3+qwzRIIuqjUruYSO+OKBcm0n2dRSoEfB7JuoPax
fHPDFLooMlgVqknckxiZl98GFOK4jlEfhnhKoFjdT+eMQAuKWetAZ2PXRmvcUrcU
AHt6/kLX1BK7Hn/3sStb04p6qZGrnlUpp4ERz7tAzXR404CsZty/tR77qIVw065e
wpm3cMfaUEkaTHXVso3g4nllmINY6QdIwiWrRZUjgA6le0C41OXCuDzoQxT+TBx7
UDJyucbYx0wcdZ1coXdo1MRktTOs2Nh+bClqlPkdePz37tCgJl8yl0wLPIaURLU4
0Mv+ja0L+dmTadowI5s8W/i3ivt47lOruzSVM5NHvC/y3JdbH01H7CQUWUrzhZxy
yR+ahP/OQbQP5CdssMELMsJgEx4K7J+x2FVBwqCnsONM7gL5SqsqTvxStOvMMrYw
Q/+vA8IIttB4/MwcY9FiM60L9ld65UECjMsHMzVrvnB7aQGTuerD5oIzo4iclWx8
M+DVGoSizih744704w/qGgPYNuJCsLxAb4pO48aOlTqVLc9lAju2KG9nwSsNkQvI
KwthuZiELfSeMMu/A8UFk8os6ffiOX+gBOsb+Ipqea9755puG5zVE2Zyf9Cyuto+
J+whtGuSz/GzbC2MGjmJ3ePMEiUIbEJ0yGjOGWt2daWavGFC9Rp4E1mCswluDW+R
YLR/HUTw4wWdsDUw5t311uPh/rO1xJtJYd8f8yDy/ghzzYU6t3tew0hU21RtbdGp
IgVgLO3VR/UbaXwStISA/vru9CCtDvPCTBK6ex4zEFWSdUzpGC36ALoJxxX5Gxu9
6BES6QkpYdVQKi6JyMTRteTOTDEEwJevxB+1idn5iR5JlRCT9mriVj+AR674i3pK
T7D8tGAk+tplNc6D6vREuFha/US+1Ip+5iEQx7cW03M9CEHYdqpTKnh/W4SxaaHk
0OKISWnhTLVCkswszEg1aZOWca8MmFlmU2HJlOVWNITCVP8zFLblp0NBjKbRhzt0
zPscviyvRdfTkGeZlN2cvSl5NLItAo+wlNfr6JPkjNSp1y+eelaAWCUFc1/26s9L
sMghQtH65DjB/SgK1bhgnzawmpSfZZYz5HzOjiasscC9b2LMSpZq5uB87CXqRDgF
heNQFRdowwE/bQ0neKb6AvZQNSsi1A6KvIw6loKCWA3kV5qFJph00kzL4sypw+q5
w9QzAKxjRT279+xUBGARaMeVdZceQflrm6sowRQGUXyoLtexDeOgALfqnzqcFDYP
GUqOXDFKrdzz7W5qIkR1cRc1Fbsji7Fo/SpOneoMfqRsnyGoNrw8hlOlijgBU7TX
cK9XYGR6q0h4O7zug0ORNfCRou5Jwj/Bm7QxggSUkq8gLSUvEVRpSJ/V8sqfjcqj
QOC9QXkKLw5ySRfyBLnUHcKZF9KohbrrI7r5Cv52INmqV+tqlZF/2MaLd7F8Pvj1
vthsSSCGTIaQ0bQpJg1P8EZnqDdIKsG5F7JyxMd+kuO4Fb5E2ZEVbqqQ3SQJzHO+
Zl4CpSd07iLJYcT3VhIrzuGETWSPJ3TqkTU92KWxJyFa7vb2y9X41aFdD8VldvFk
X4yVKvqjlHimvLNONlTndpi4G3PCl4tGhPScCOy6qnUhQqk6T+TUdruiSfA+c1L9
iLVHGrvT8tVWr+j7IuKUIyI6lOVR7s2tYT+ukD3+GcDnbiXBixz0q4+KX6M3CpRX
3t42Zpq5icMuXnX3LLQQA3h2Qw/Ca5hiPBjI5XdpLXUbuSDXitW9/jiLs1EgD6rd
qEUWY4iOYOH2gZ5e045b0fYaZflDltx/9iQskMj9O5CIsSWyArWAB9i3RvAeVmtW
NqdMIjXnGMKPF5kkRADSzD+LobMDy9mpkza1RdnDn4Ym552vsRY8Q5OE9MET8jKv
m4leMbYg1rxv1Gx2chIrZzT2T+9JBpZSoMGVgXQ+sOZSQF6jvl3+m5sV2eMZ/yiJ
k4/nrBY1iKx5TCfX1sScpnPWnEOpUPb1fUGy8ZtbIRMz4G1nsYOJERVmD84SQaU1
utr+oaOQ8XLy9t2dZUOLxw0uUePuEGZl50kfnwKO+153fnruFygrL6c0YvevFe4q
c50UdasHhqlbnUGfs8GfCA7AnXZcrvmKFKkTB//waBZJl/5BLp9pkaghouDLUUjl
exgNpsnzlM0fARXOXAixufwCgv6v6BhFeWgKh42lR6MfCVbArTu0FjH9GWhyFyxp
RyjiKi6Q6f7uGbVjiHVPf8psTSdFJb+dhNvbzpLUsJSZ12Upo2GZVH2Z84kywyw0
t7HceXAL6xl+r7RUyfM1e4CsFEq3D9kXhtpU2zzsKzW3dxTJ0U7zCyP+DSuUxq85
7GPNftqase61/ID0mJ2ry1SU/XIQck/Mv31r56ugMrbV64l8f/bj93Z5s+qoVofK
yTKkoMw0owl3GDsGSQu0c4UqnuZoLe0potLqDaI4JBNR/N2YYg/M297OTopAAv24
o4EiUszNqf7ZVtOtuaPPOGL7dCxKsZJtsFYKjNbDa3rBrgIwCHJ0qY8AvHV6Qxlr
0rsP15iSclDguYvggpQZFSJoQrDcVJic/wfMQ6fCriGb28lWtckS47zdkRTqG8tp
pkxw+r3wo8kcDzISN02JSovD29Q0D62sz7GR04dDyZT7kKtLuOc4Y8Z9WMzp1gi6
kHl4C3ceeC1cCcdykWZRdnRyyfSGUdmFc0BN3UCVssyZYez7goPYYtI3eRGJVRQ4
mFN9UG+MZTnlFPfaonaLnq4E7fgyS0ZRjM55clC+H9o1iWrUZe1aswxqC60mxl4q
VWeWuQN+tpFQmT+ICUsJLuYljKe5ULLDa9yweCzU2bCd8JrPW66aa47owlwoeHVH
Etqi1ESNfEMe9L8XEIQIHEpaBREqOk7PVofIe1lCa3Xl0OUrMnAxJf4/VAa0yvvv
IYNbOg3FdPp4K0U/H7mMVWlB2YXPFA6Z/f6paroSpoYvjaCCueam/EYtKLqVRV/m
SWS1yPvPOk8XwT9AsKe3Xzpw57UD+W5Vv91L2dcUaYJruOdcRZ5B8POWCIpwdX0K
222WXocop12FspbhgofxNy+OaamYcEFg1qir2XbExI0jqhkN3SBeHHv6+059sQHn
99VCS8K1hkTHNytRY6Wc+Aebq2I8S7ioqielgcFQmq+hZ2wqwJkaYCE+f7+N77E4
q5E6HeCEGHy4fdwutThdxWscfPg4az7bN699Fs/uvvcAy4oBMD2PRtK6KTXiAap3
XIOSPtPPj+3mFD5n4nvhAViZHLX+3BZlRGlElkZ/Uy0bH/WGg+MOBqg0XjrSviq+
DOSGelsP6Q9gqLOT1lmHb3LNt0+9Ep+xdAP3/SCIS+FqdeHnZfE1pkpmM7Rvp891
6UrLFz488bGeT9XsDCkdnb0ECzjAZjfgGP1pNuBCSmhlauKm2NNtbPBVO0CfjYvt
8oqM+fV4JCD0CMQpiBEAU24Zi29IOt1E58j/ln8wipX3uCOu2UIsjsLaQglNdK4w
j5QrwNGJpZZBZURMOncxji0jZxTeDMlVNp7RYunJrwLqev1sZTUFM6pq5wfkQsnO
WfKpD/ccAZvP/ixeQS730b49pL+wfNfGBTp6/d5FiAPOUR3GYfT2dh7NRrIUxVBN
pZW6NEObAyUJjCaSOFRl12hwbis8za8PaHGJVjOOd0NOsSyL+eP2c4WSmvSaH2db
Y6u3kOSDFyOT/nZiXkb5h8RizkIgonJZbljWgCVXEp8/YhLDCjQm0yDNYWghmz7Y
jrwECb5TVhI8ZdqVGT+hMsJeKx1HDiGLf34c/D3M0e2NxPyqpYkSxkS28H1G2Cba
z8+eGhFOHK6XMj8XCaoKP+UjR5PMzztc6orFuEGuy1YGDM3K0oD7L8WKRNo6fBRz
hcUAIE5iX21f1Ksw1IgGWJylP6NX8gXGe4UCg2evuZXw2TLJWB3sKAK4iM6Zh+av
JTc6DzL9hwumY5K2l5OPncaIkyV24cvSJsaui8oqvvBawFS0VBYCNrOhxqitQSfi
fOUsSJjFomXKUjFwXymPVLRz4mxiSCgwhMpm9Ag58ZcVETUzQrbWpg03Xzgm+VKP
B1ULhCB9W9nwxHQd1un9JdonmbDFHHgdAubr7CDIHkuQkyfj0qfKedRP7n1WimNt
/rwLQIgZ3Zcu94uUySTV3vHoVQkOVMbOomRi7FRFHnDU2Y2eARpES4pxNhBaEx/o
vtzj4xsRe1cQ+7mjgJUCyrGC9YJQWfXYFzDRDFM8fjuGWBMaAHxDpkv9dnQjm3pu
dtiorx3+5jG8Tc/OETkdhvEFxkuUJ6VwmvQLTwH87gwElW/ICQaHBW7yrW06IKkl
5+tQYKLyhV0mmbABa7brlCDFGW3AQESVNh1sMUCx/bnccNMN+fRD73UyTGiSW24U
hX89YkmpIwAwq7nN9BsC0PQzFpiz6q9hdIlSGNosrhxV2G1iVI1a+/p4qj4F3J7O
0qHUWfwTEwlsUZWrT9dVC2jLZqOUbbMAGUgv/a6g8oGSAqUzSWU9HnTWoOkslojf
VCpvu97MGL78Yd9HFAhcD4XNzDoxM7jsiiTumBs2pi4rOCpgooQI97lMODJw91Co
Jw37LkniI2CbFHhYVIdMfTDKdaApcch1tYHaUrRsZd/KUQgT51e2jD7i7iVakmsY
g2H6DUbeKJuAzquGFg8vLzFWa37Yib7WoE0oq/Y52NsqUl/ZPFab1J2WsrV5kqti
zqVRjKXP0BQ9W6/T1ziWOQJc9aViIGkba3PAVhgtMXeyfAk9cxXAACabtdLG4eyr
XFUM1oF6/iLNUgTSFJRFx4RdClYeIdhOvwA+Z+UPHslS4a+lT/f2nCn8XRDSMjf+
SU3nPPeJfEHSa32DWdBsbtkNAtlvHN6sLnfS1p/GUdq0kOL6pZqBK5+4eBAB16TX
ILICB022LnDCsK1VGOT9jh71uy5jMFJ13BwJoShspcu0jieawiC1Dhk5zYY13bCB
vuxGKGgNRCvfbFYLUOcsq7DQ/VCeavGy9PYgaty7k2egzt/5u/sYhdw9FNfHKoVw
+1axR4U0iPDdEtDDLzeV0xTVX07yb2ViI1T3PIMlV3CAD32bLDzluYcVM+saKGfk
mIOrq5e/S4mqgrgjFVUrufaG5tgwwZ7qHNPYinxawjceJuA+SUjkzfAS4fnoCv3o
lBCmMhy8xX/fNTY4rBoWDecvWxuDosZgLCJbBo/AyXlIgdgQLVgJXT7Se75qYOKr
CqBvaGKVHZcMl9KfpR3xbBeSJ1YPFtPwsoTbdMtXbtYQjTjEl11lwaPcbnME+6AS
gGzH2rsvHilOIbMcX46WP3z0Zsn5yBdyyNW9cQ5QxsN2WdsZlYtmc61dew7OJhrY
6TBna8I0a+/KXN6zhLrBjEd97K8mimL8U2TBaCkdybZBNf9kYOkowmdKFKzH3JgX
Vcm8Q3LsWmoQEy8QDeST3EB5A40wIegshk0f272eE2R2WCRUsmcixwk01hETJ+N5
i9QKLGR5wWb6rbmHyUqmn339+yPiSHNdNf6ru7bUh/DSRVjnF0RB1NOiOBOvsjuB
YJ2tXDbi+6BCy/QJ6PBsL5lvGw2BdCLsxjLEmkP935/k1zGvBrLCqqx1yIHybZqi
7ZRvaF819CHEmFqaekboyyjp2BgaL2NBKJxg60WW1/pJ/CYI3lPZXykJ0qAPGk8r
PN0bkd/7hv1iKS4D6Lbn9P+UZqhug9Aq5TFmv9o/zWT30aZGVrVl/Yxjm/pa4pf3
e3AUjiuTaRWX6GTQ9o8cta3GqWLrQ8bKvf84FX7f8+9wCIQNkw8W8ooke49AAl5L
Di98vXvLqkY24yEavTK0gg+HxvoIdoKkAyDLeixYKWt0i4OZ/DnMlGowUiVsXKjI
jgfZE/ajRyB4HRj+Ffen5pW/2W59lcuITDQ6vTkIwC4viyhAi+vnObH2XA7LaqRq
1SivCjFU1WzT5lARe4wtuim378Dx8AdYiQlzL7a8ygTs7OxqRTVyB6XxikgAfHYG
L38iPICQMUefweOU8hU1CcNDaC8TBzxTnFon9RB8CUMgZLe4+GgdssoggzdSKU+l
fpikFj1LYkV1Ocbzuocle7e6PoEdNPKDTOi2rpNwrZPKEQiixaPw8QR46i2ZXYWE
lPfhkGOS9oEt9gc9ZvwoiGyEqBtojAwcQ455g0K2qvwBeluwZZ+ss9ZwEsr34OH6
1NhtKeQg0b94J9Ed5bqchBVo8f1/VTB3M4ci/A+6V36AP8r02uPLvNK3YIz6JR5N
OBTtjWvwnS++L6yevVa5+JP9Ex42/CHpv2LuI8zy2GnOnsf6bjmIsvLbw0F1bo2S
lTKfUHuELYaRl/BPaXA1mcXs8+LUEqMH8ulGxaqk//Ig3/gCOLWYk6HsLv2h+gg6
CkSi66Cbw0Cwq5Lnt3PVmWXmgyrFPgvXUzdP2ChFox/mTOq5OTUnbS1ww5aU23/J
vwQvT+/ggbVhT1CchSd/fw7R/nHF156TDpDUW+iS31jucRX+mZ8seXhA1CJXSfKy
AR4x5ik+QobNIlfHySqlXCRQAoo7cJTK/r9lnUsidlSzi5HXkHq6Y9YdZFdv/fxX
54OqKqRRC7ugYkUzaIwnjMgXo8pM7h+V+MR/cK2itABQUXVSv6jECJ2OSdrg0VHe
j5pMw9XN7xj74GoVpZySqoUZvE+D19LSj+0KRpVp93uN7DR8+WEPDQ1bQPsPEe8B
IXGQSh1z1WRK/XY2JXo/7N5QiKEVHfW+BF/hRW9pjpU=
`protect END_PROTECTED
