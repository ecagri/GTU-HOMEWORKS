`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T81bn06AxttV3gMcItuRukPL5DHQqg2/MajO6EYt8XeDAiDGkcdwlnhjzQOwVkf+
onJPBkk6TqacODgYRuDTDS4V2MriGBthEme3RKOzjk7US13V2WdzAb0rSq8EKlCE
89RFL1ONsEXZFZ5otEyS6rDhRLDYU5ei20JZGtdcwBhXAJOf6Rj7PZ3bvAyyWsZw
3D9bcNmKWSVexoCq5Nd/zvVGVmAtKG15gwQsV0M34AMAxd8siIh2uSnVRwV2d1W1
i0wk94Y+3iEZibsWC9vhw3NYCH8c4lnvYb906warlwJU3FRc9bj/bfFI8lrsPmRg
vsN4BCa5iJmkrsgRib02Q5N+5jk77+5LXwfjR4GNmi8Pu2anjI7kOUS1Nm40Ys/m
b3g4gSwndFtYMMtnRFrYk6IVhVxHpe0sIwMppsMFnC+0EpfVIrhPm7NB68PASiwY
0dr2jGw3XV7pmcIv1o9l32lTuZCXeGDcbXDHTUKNqVAeF9pXORYMwNIYbjsjXoE0
xPpfA943VYrF8LdWgq7iV5fRLk0SPZxllsbNEF+C67hnIUm5Hn6V6OtVU5fZisK3
AKXYsdf1fVKmAk3+uJ9uPb2+tju7rPK6XqQxywdR5F2e32yuljmPrnmP09FNNXrs
X6Om+tkxPBVXZ7NbApsgVwroBA2SA9dlepl3fwwU2ch4hSHbCpGdg4664hk6LALT
fbK+uavMd2kFidc3pTV2ZlWo/nckhZ/gtmnDuRJJDxqH+WD79dErFgoUD2AKTkd5
S5WXHPSOVC/E7z5j8RV0VKuKUfWfZrdbOdyrldthCKdFmkQlXPqv/0qGoQPQZDlD
Rfqrz2htlSO6NcRrdf1fWfvEYHgCy+v1cJ+pLskLDP2zV/RL4LhnzkelwVCZ8Rh7
YU+t306MSJUUZFPFlYg4lXfXziFaHRN7IK05u+HNpZSKEdRBgzflKfLZIYIBgEs9
oxo4ObeRRUGB1PQeqDGMNd0htbUvLvCrbqfpQmlKFWj23oSOESCyt9B1U3zwPhF0
iSYuXdhXlTyXduDlu9A4qlqA8fuUVjqPn5LBGNaklN7cG+h29ja6y5aHHZ3Q7qOa
vGgC+XmFzKlPi0c4eKxbul0j31XS5yph14xrId0NA6D95Pf4ti57UUDHWW4/VJzv
z/LTM8F8/EjrC6HdJulsl2zAonJqmF+GfUgcay1agErenLXuyUaJgteliEay1rol
rrX6+DsbAOvvVX2YEwQFvOWKgCqmHsQpKaSazNeNxg44ddxNuG855J8QlyqNEYKx
`protect END_PROTECTED
