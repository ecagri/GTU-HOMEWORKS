`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EybGcZd0nVzxTisSLPdPRn18iSR6yYWm6TIHojQlovoM7C3Fa6unqnViESNDgJCy
fSIbGhFl5QmQd2X0V6yy1YN+HUXQR7q5HGW5zs2qdArSvypGDC17Ys8vg/EA/p5N
Cd2U2WXEwSVHELgyu8M5tvSPqhJqDpqgQNfJtfD8It5dVZypO168B6c0hCctkhs+
NhTTxqPdTQH6qEQTYMdjy3Z64eizFhqa5ANMqiQy7AKDwciWC+9hQm8YqLoXLWLP
m77OccWJCUQwCdRyO27MTOiUORqSRwnV5QoXuxzuKMbgtDN34zp343hbEg3fj9BB
AUCUycMZUlyvcbyv7FaLkeOK3kMZdo2sux7of5bAUnDIjXIFWfNHUqzncs4W1D9f
jW16BI+RSQEWLEHA4ulY6mhZiRDOHI5pFo1JbRpWNvCFSjcWYFszhhMgqi6W6QT7
apeaH7VDcvobNhpo7Pn6uG/OYXt7NgCffjc4VwgXfYwt4kwaKJYiiHnd/BoURs1t
HB+AsCkhVtZNTUse8ygowZy5IkC195lTr7ALnluIf223SYYqLD7ZvwEhT3WtQ7Id
8xhPqspcFHn6fmD+LWF3PnciyYCbUwmpKpnpduQ7zTEN4VAQeaCbASIkYopQxrNi
GGnrXXhJu8ffxinIRuTxD3OlGqYundxPqX3hkWJzkWkamSOEq7kA5dOS4eJDj9SW
vfP4m0uUPg35y5QBuJJGtiyXsj06biQGU158IsxiOX7DtcGWZfWkCPMMJ5KRM4yZ
MNBA98KcCjx3GPR5/H7wMuwlU52rYLl/MvmeS8PL0YHnSs5Tk1E3RHnuatO0VTFJ
foNNHPZ+2NM8aQruczYUkI6gyvs6nhAOwn6sOtncyIMup+YfHrHzqDCMfRsHBPnT
fY5qWeYZAKpQI9PYCHc5Nx0rPSIQoKuWQL07nPbo6LIp3VC2XuV8Ugvz4fkbngvG
7U7d4DgCW57bv9Y5wj4+4MAnzrPM3eCjIR9rYJ4KTZJ2p74dgILCYAprUJ9vfA9o
7RPUW8lmHzyQUp8nijpwgvIHI2HmBMqxhsEEdMd2cP4S+ahtTVxdd9nx2JpZhm8U
ZBbIK7lU2cO15O9C3UCEvwksy9T+iWeTKxhKFXO2ShOOljgJPqrtf6Emef+nsEeY
8WTH+FI0uysBQwlyF12oLbDHOC7buGYUZILeqlaedlS8jSgbhqaMhV7n3/ewTPhJ
yU6e3Amn8TJK/wgKIQGFr9sWjAawT2Tk+T48KzS5tWYdx02RpoUBwZ5Obt+U1elr
ViPVtmBXwsNgczYtH1rgx37j6JrnA6Y0B6l+3AhNAy0Cuv01gR5iPOL2GAzntDWd
9ZAHthRB94xoJSO4rSp9QRrjjUL9VDboxD9UjAkRI0B1NsD0u2uMTD57WHKFxW7J
kUhG7sIXzuxesiCaHy2ZQG6FqpQqbQR0Ix30kcUjeYlSKCcqlEODojSejP5psB21
TYuCLeH7ideOjcr5ypXQA/s9oQ6E6vrHOWzhGFsA5Qscm5CK+wVxWCet3GY3QnpP
GeKtaciGKyc7gtwoo/QIW43rs9tliSV8KZW3zQQpq+6MS4Yi87gAxWzMkYAnhj1q
Ttp+sx8o/vNpCBRNpZWrnwDlg1C4/Br1/PWBHsxyvaIKRjDMqmi4F5+d7qKOwlwi
C0m5eN0MZOavNHrM5+AcIZj+HcjGOzi+XzXcagkX318RBNTn0nHs0qsyI5QhPwhC
KKzF9XUeiPUBUrk4FUXiQ6c12hjI+KLNGLe3/iAHp+ptobg4itteSyZOQSvt1FWc
2+kmmZauqwJoXU2ztasK2j6JGPBuy540npnt+ad9ZLYN66/zfgOkvHzrmBACk7fk
Be9yIMv9Z5Rk9fgcillg7KErySwwBPt9wYf04nmRm0cfAVq+YH0P2yT+rE4taLXy
8Oheniq6wip3zcNsB+0R9aMMQWrvEOpRmS9/st0/JATR1pa7wmXGHuWytOKbAx34
6gMLhkGFZLIQmTvRbcDw21ESc7LqSleorIlb6uttVTtVQzf3b/iJns7EPm70o0Z+
RKqRiha6y4nw3MSLbydjgAZUqO4Ei5a5F+aPP5idFL1W/+8MJ1LdaJV8I0oBbX+G
as36vFMttubXW/mCqWcnPy9mgaRrcBtXhzg45r2SsrdvqCqgciuvRQr5PeOBmz0E
4OpqVX4Gv6QFBeIYITFtyC8GaM6xTdkE+BdyUO/kWy6mnqtiOoPx9ejBQvkqtstm
2ZvDv6MZZoHg+exxPWOJyc4Aka1x0ddjWFVar9q0PVxyBGVrN2V/pi5mdpEKPuMS
KhvD3PLcvw5a/PMjYwxrZTvzAIhvb99OamgW/OfjASB1XsyxSrPd8E5+1objiFXF
OLMiZY+4qLYZN7q1jiXkSKkkiFktG28J6hx6btufZSUW9odYT6/wIzY+7IbQhCvC
vj3or9TIBj86DueemQ4tzhmHT79YAyRkT/zl+9EuhainXKiN7MTb6mzVmdfleF5V
ImGnEqbBMvVMJXi7pP21hBvnd52uQxAIoDdiYART44y43deP9X/l8e1fCPdt3gMF
qi0tJufBHgB9FlQCepFpSFlkTeVUqNvg9xKfC21fdcUyz8uxCW8d5E/apihLMd+j
lKKp0QOiHk9F+LjbL3NBTDoY8+k8fKuJEdO4lB6g2WWnfbGckii6QooM1i1Yheie
OlV5+ifX4pDjOKWZnHnE6z1KEav9YvHWYDxqAkmdI3SUW2pzddWYQgNnWl0PVVb+
7+7fVlWvndqAqspGwn+IDQJY/DL/2aZN5EKJXso47rmihxxAKSfAjh7suqebNPbS
127sIVorPIgbhLcWG7vc1mJQ/DIqgNtX+GggZFxvCByilD1GdX/dNikcHfnG/G4d
qtBFY7An3SM+OycdQHBamCQK6x4t3hp5OfNFfEs70Uv0hP3aAhXG941mYD0ppxwn
K0ZrHM6ZFKcw0dpHgk/HPK+4n3/Cpf0EYd1dwRPpA2PyDsbLazp4j2lOQNmCSs8q
7zvWNiMo3JT37fXVzHUcvmj0wxFuyDzb8Rk+43jKi6hbWmOHsSZh0KUVJtSGCJxN
2UrSqcqNuSxOEyfY4jlPS2aQQC9hF6sqskTmy5qyCoOejTEmo8qIvvng1bLKaUsU
bgCBCdzfx2H6e0PYLirnzFz9fZ0gB+DKKPfGgCpnW1XI9SiCOJ9W/K4gBDw1CqSL
Gn7SfWrtX7vQqK30Srx32xcOz5rNz2rA7KOBtlz+0ip8AX8mqJLGly2uDu2KVSal
BdnpTB/iTKABQKiT2wQhJlCZwPod1FnLGT+LJ3/NcHG8oSzD6ujE4pHcGFh4MNOV
cCvJwhZr4ungfzfw6bwTwa2Du1A9I8CupsSMguILq4jwSPL82wT9BG4kFdTOIubu
Vmv0nnGmCcdTTKn2vvywu+S5dYItlkR/6qVbXZOVbiovFo6Af9RsuGOmShBXeL9k
Hkk1qkH2UXTJeQFnqUzO0uVNhDS8sU/8pDU9D4D+xJY4jbrDcB5ciRmtw2k6dBlQ
2YrutfO9HXfQR4739I6yOnAPo1ofy4DA2Opm1F0I+huzG3zvtMwz4qWceyEPhkDN
/BWI2UiFhHDqs2o4xKe4wsw5FAeTwuJ/H/98V1wADw5NeHS6POGzs/k59e+GmH3U
ubLUhjdrUp9t2TIENnAIzPTyDF8gfPPv+KA+PhZhcEt5IiYWQq6Hr94vHkpbLJew
V+NqPPjCsOGX5lZytySjOCNWQwmXUBnDj/yPpGJjADVPajU5N9Yo4/V8NmxEownE
9nHAf65zYK6uoicNeSt8YYVQNx6KrV8OCihnDKUeXJcEzW2AGfkgnPTonw8P4pW+
PqbhGFvmV6d0loIulQ/9jPf/iiqiBsZVYqV5J6LWQ6+hUNyH5l7k6YlFAANXDiDB
E2mcW9x9rviDAu0JBbtuw69px+30/5iJC08d6Hct7c3ansCrNY6U7zM8bQDTTuAt
QEUv+m6+9fv1YyK1XK7CzHt1tGgkECRI08Ap/UUgLbuovz07FMj1t8FoqifFERds
XHqpg4WAiNFt4e6O88USKQiQmGq4zpkvl15zcRlOa/MVAzuvB1aASdJdSrYEnBd5
UMnnQlksvDmcxSBFcOhwBtCAq3X7cq8oPwiKFCS7kEskW1zFW8o7JHfvNscb9Ca9
NMJnjZf3DCMLGYdUPI+YJIK+dZ9wmHkVWS20RLGiTga0CLnSJ1fvLMf2u8ahn5qm
SsHEDZJh7dgLpeHiIT3fHdarbSgFkksuCtjDz0HCVFJVKO5i87XwmNkDsdcteLqg
2uoS2jDWhxmDF6H16FW4x9Bi5weAzwv5bqHCtbRl9UH+tFIXtEjB3jcHqCjNjjH4
yIUjHIN9lZZNqqLWZXkAth/fse5dXpn9LXLJZWSaFu7kgLYGJXWK+OHMBmaz1Eog
ZRf1HUr94aCdpmyN7Z4GPwGVxG/RVPnV4BQYpyxfbHxw/i8otVkMqLypwTcjPGEK
9o1Qt9BsO+3JybeETlN6jKW7LscmHxfCGY9zlNMSnoWeSjefG8ApuDhr0EeQrC0j
EeimBH7czVm60ccxQU6E0aP+sjNMLS81eET7PeVH9ioC00g4URYNJn63mluja3HV
YdgEYnSkRv+BkW2lOxWNKr3EQ3OA31W/HwjGrWbMybBTKPz5guZHDP2mHwrSAk7E
4NLoPktieSnE16Fh3uZe1OyaHZap8PJqeXStfaMfrxeMqslpqT2Hpf/JxIWrLW+N
lkKCvTheddNEat5Jbxx/aVeyxp6lOYPToFr32UM9ykxhOSvIopePW6L29741j0MT
2WkVFW/81Di3eQqlJXANRuGG8vfC1nn8PNQULU9c/iBAJkaM8h4TLF/M1MfCIf8a
mWOF2zzP+IxtLGrTFIJDM4M/PjXeeAOhdFcu8SPZzuR+O7w47aTTcsX5zm2Gi+zY
ifZojmOfWBNx72sUGzoMODU0VykAPUbBn0OEr83LfPvHEYNYolU75jLoov/XZUTo
vbzDnIyYyZsgDFgbe1rgHaTv/udOntcx5HUCdYsITZ+FjD9HWLaumkobFe4JTKuA
X0tSEYZmcecy0bH89pv2hQIrXpLmyJdN1xBPDyZquWxDNkL4UHMjaHrVnzLvl3Re
fZpRib9Ag5Npa8BXbVkPgublcrpRwXXlllqEUCDEy71+JursvHlh1w/mi3B6/FoG
yzwX+doeKTqYWfDqTuveLjyWJQhezUv2DuAQpYvOZcw+CpWIZZdpfYywJ54e6DKX
GerW0C0N8cna0wKW6ff9LHI7T5kwJ2CgR+PUQkLsFsVwrD2J/U3YVIvSSsHfnYI/
cI0THELljpNgYPP5bscrWvbLCgch/5L5C72eIMaOlGtGcDUlKPSc0Mhr0W19J/Pk
PydEUdosUwq6lyLattQ/HJ4Q2TjPuz639InktSXlowa8fDk2LLM0ROfTmvxLT6Ci
t0/LAcBP5R/I8r25cSRoRDvklMhpW2ea2sQuziSWbr4pVaDfFa2m6EvCiCmHrvfb
Xj0hsHhcbkSmg0rR5Lqx1RHkN3eHxk8QaOt7MdlceyGwWID259oLw/4VUjQ8kBe8
viJrYXfkNI4F8PqXgWaXHkzmLAXu/E9YJihOoPmHya0x5YLPULR4FUwuqP3KleZz
2Ysg2ZxjfzBWFnX7H/SIDgSbS4DCrUP2bMXppAq745TmWKK+CJc2lojEOVvtLT6O
sT/d9Z64WbuyfCuDUK5VDFfwjYrVSUnsc1K+vffD9NTXpegraBv5QydNtVd/DJCS
sfnzvcTYxAdn5TNEdZmTiRZEGsRLqijflXE685nGAUcyyWY7c7lD8Ly01i8pfB34
ib6PW5KFXqA6ZnjJ8KrPQnTgJ0udS4dVd+pJ205nWrZI6E3w+SlayWYBxguTWVtC
fHwm+8swo411RVQMyquC1BiFWE6zTmYDTkJtCtbmLMZowDCeMBl5sZ15ge20J3/3
`protect END_PROTECTED
