`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ILEPIkTuNcUBPqQ5JrLRAcrVDDapfkrTVLH5wcSQo2jgE3gry8jcvDIYadIh4dB3
cQ+tULbKUx/I9OQmKlRbuQPXfzPzaZHW6vIbvMibUo/kZtYsGb3MtxIlMPs4Tvsa
dhXGD+yP+CrqdRIUP4dDQqM0RNqdMO1pRSfpoJIfzFwcrJ5ZVJGreDZDklFMRX8e
H8bKE2WHCJiYYwiqxkHcDCt2jYoDtqtELOS6Pt19ZzpfNLXLwoaByGkAYMknizyQ
otNV4TPO6Zi21fJmXDw8VSWLNo8eroZpj/q0pm6vidV5ZtmKHYhLc2UXCCXFghwu
CFdKbC9VtT7eCukBUF7bG4o4JRA4ItS7+Hg/eALIKzgcfDFFVbTWwiEBdwNelBlu
D/gdWBdkNVcDtq6/pDQrxhIaFeUsSRYYpeM7XipQCF6p1H1K2EmeEHEiFw+pfzPn
p+SS5z2V2VJ5nPH00mmORA==
`protect END_PROTECTED
