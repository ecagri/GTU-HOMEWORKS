`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZG+7H51CMcppUhOAsR5YwXJrLKEOZw1H5GrnwrZZkFUsflvuQKh+qpJzkPcinsL0
kjBxesPpq4Re4cn4T+lCWgKQNYbsjytIiA2Q6y/XCsD31vUrrMyQph/wODqoggQf
K9nFov4GLIMFrhSamU76pc+BZrk0pqpegxHF2euCob55ZxuJquHDxiX1EXmo4MGw
cHsNAkpmtRj2U4AcYYViltxDrX/inoxPN4jdlDZznjPI3Cr66zm3rKpdeeMt5XfS
tGSqkoG+p+PEip41RGj6JZavIYWWRNxVVJqnOIaV2Xesl6GXv+4Yck+HXXhCcB/A
V9HgQNnjEQ56dwFdiMShJiDjsEcZAgHPip8ISJ/uCmeYDeRQVvVHESKvKUCh5L3S
HOgw1niM82DrNvQ1TWi8c4hQWpUJxAG2qaFD9U/Kopir+WTlmBHj6qS0MhU81GvS
0UyrXvs77Af4apmTzVsAE6iiRpWp9oTgsTRxWDql/Jc7zxg6QF3eYhavhG2cevG3
qXz3TDDhpEcQ0XqYNyCEGg==
`protect END_PROTECTED
