`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zySZ+7sbiDCEsqLyQlVaUhSah3NEm4RlcpX4rV31oB5rQo950Nhp9JLJJfySezGf
C9hxmBDU1OrLy4/Vzvz15bOggW9CDylN/+ZyJ7qW1v0vSSXYE4nBIcuZm0JtbfQU
q9UX/83oxzvo+72WlbYFC9m10AHv4GN3pDxgWSRbPhwVO/OE4bdRp2J8pxXBt94u
btos+7v/q+jfEEVgRDMz2jc9ss//FKmKHEaphOM6bgeuxH0XYQIL6yPp0STh6FEJ
05829g2ti2XLKT5oI4XLuYUOB8qPQothlndYDu/QpU6MQ0IAqs3geIGGBeWEL9f8
orBuuP58R2qYjaw/HuJqAMujQ+oqDkjTXEeRvRfgYwTbujRQiSlzL4i4tLs1Fw2F
FDxd+NXWraNnZ/uzu2MqAS4jucU2vBk4/z8BIl79thmIPolqd+ZUbYa8z5GjFM/m
VlgIsGhnXFtVXlV0lad6F0MN4PHFmiUhu3ZrC/HU3NPHXsJYIO9GhVE/XwRjbtVl
SqJ+FSeRYKOZBYvL3Y7bjvZgyn3gN91gOwaQK0l0624RBJtslCebaFwkfwuXzn7v
F9jfrVrEeeDtjF8+jxBeNMbXPd9F1Q8KuUTPmAwYGoiGcu64w1DUi0rCRX/bPPcy
kk0RRoxTt3iuObof3bNhVyeuKNDmL5sC/wUcG7Qb88Y39M0K7WilHTlvrOZiUtil
TUv/KocnSuZXg/W94040ilaRejaiikP37pYe0H2IPhUfGOX1HsMs8e4/HvvJKZHo
swrSiPUyvngcS6ZKJwyB60EYsmEfMOj4/AlMyq8xuV+0mpqHdaa4tY1t6Aie4JAc
PZ2ofZZxbT2OMDeMith62DGIRFObpaevUu1qheuHjlDrGGZxGloovWO85pbf8Flm
2MLvufMhSVHBciknuBNeSKoxUDaOy5BmyyIPXwA41VE3B6vvW33HQ5cdI6LgB8lV
0v1V6RXQTTYn3Rm/q2Eg6tgRgpB+TCov2bObYJj78RXGV3JlCXg0pROQcsbTnrCc
D0jZ8Z/FtuQdgXvlECz+cjAiJST34d0x7vbUvQrHeD1Ubtb9gD/4UgeBkSGVeQno
PQ+kXfOlJ0J+vfUPf7tN0Q7JOgv53grL700gQbycvuZ+7m1apkuWOEGyHRSm4ale
ObYP0zhOvIAF9Xv+cmcu04uZIdQob+P3q3RnV/iAv4qK4tDkGIknuuePtvtPbk6S
5LKicoVY1RRtshHAMF8tfDol4eZZQPyGMyBm4Z4XaBqeXPJHvTSUZyhMt1gOwtVx
`protect END_PROTECTED
