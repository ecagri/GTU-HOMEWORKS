`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+VDkY0fl7G1cxHkgJG0wkfvwHY//sJ3UChfuUAqbpbXb5S3SdPy4ESNRQ7Aq4VSd
gpRNSxsPHb28j6cXYMBshZUanYMbRFPQ1CLLGthFU7T6MKwRD8IQMewYdzaDLzOF
rrKnDTy/31OW+PFug8JQnQSapQTtGjxN+Ir8sjs+f1Yy17gmgctcQef3QbzmMBda
YxiakiDkjHNm/tH4NVg8PRwBCMYsWFaV/mnNRVv55X3f/GAq5Q86RiqIMZz8T6Qg
SqR7rtXVSW4ucGuz2tDlau1rrTT8NQRs9xBNY+B91U/v85EShOhDXx091vwFBvPA
D/hmPA0N2EU9LWiiNCn6wh/QixOcHlezNQOg2BfXEc7UtfE1eMJZtoX+Ba6T290U
mQeNyzeuKweYJMjd60qFT0ODM8xSrYGnmLV2YRpnEms21D2YVS+0PERuURoVDEGJ
ywVszuSEpB0xo7mIhcqJm3UuagwbTlkG3KRlZM2n+GLhiwOuUXHZtb+7377oqlbF
1ocIpW+T/R/21aByIqnNfGlPMvRhWG58EbYocXEIC5sgoRooheWUjf26VsESQ7Kt
xamfhOLI1TrR3t7Nk+N7VqRcVWSR7RMx98m3xPvyE/m8FwcHGSJ1KrpLYPJz9XZn
WvYWdvIMq2YgQaNVAqn3bydfzB6YBrWV2tucBKJGdtgeh4XQZVqL07MRNKjUYTaX
S8fE3QuF6jLrVSzWOSZvQGh/qt6dQKLXC6EvRYVPEJElORmarnsU3R9lxnBGdrHF
7NZldLoV2uTqsxcYi/UxI8cafjQE5gIhcXTUwvZ6r1DE4hWekolQDWbR07fGfLoX
C21tX0m46Ih+oSG5i40EjsX1cdv/Vbhe4paXaf9SplGnce1Vt21ty5INmibtL6ZE
YdM/hic5zIgfCLFrYdJ5JJL+2+w2V4DjBiy/hrsQeSORxvfRvSe8T7NbHYCJXcv+
CoQNIxdRztlrPbd4UJBI8aP8QPIYABmgIFECFum/11chyaWSSzGn6Bk5sWgUgpig
1HLq6XRfDvb1DcYTpUMzLZ1QExmVtGXlHzSamwIl5A1DSfY4vbKKvxvRCKlBPCOe
5HnxzVwgoTAQWQhR9dg2EhAjVMXSoHhNc4Qd6mHxJ1M0NfYskdaOkX3kYozRYD0j
nHeTmVy2wNIocJ2VqsX/1De6OxUuEEMW1l+V8VuqAia5zThfY0e7nPO1rGneHT/q
n1Sy8NW4J4i+EEbi3K8AoB3yNFowSIk7xb/CQtnoCsY9CbFkIaQkPcueEfYK3Vq0
UuGbs5QuWiv4mltAWaYPAJDc8k8MCjz7diYK9EpNMd0CI6S/zz1DgjzaQ2iYv9NY
Jr/dfVDNbbwwRJQTP/idYHvSYUSewgeqi5erNIxeEcrsS70dLwJ4oDcPIj5koKir
0YklAL6+Y1stC9HhbNAWBIaD10ug5rwUBEBsxduIOfNL4RWciMgRzpFc68sH3NWZ
arDLBvM5r/Y+QjYD1sxg00f70CbkXQBMZM36zh5bAaHWnu/K4NunWeSUs0vjd7iK
9H0vuYDtzqe1C1Aklo5FYTfWIiCjFnSzBrcYF9CAWpgs+5R78wVFEiUZj2DQ8eZl
9hGOa1f3yknyZEx/tR4jc5GVGdcyd0PS/LlK91W2Af6xqNYWGBbWJrAmAu2rx6/2
WlyBhS3MTVdKP7BuurTasQ==
`protect END_PROTECTED
