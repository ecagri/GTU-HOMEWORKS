`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9U4hr5l52fS/EZCxUF6Jm1JeZv5qFyXNBtzk/VgkD9/vuKTzp+wlI0fjbyoI9JZL
Hv8+i41eH8QavRA7rc3iUK54y2526L5W5TXzhWV2jCOaesTNnMYImQ6X5zwdMpUS
D4DrxTG9+NA+OrlT3MKzkDFLi3498icwYkSM3PIzlpeBsH8Kv4IykQLBd7vQ7pmx
AGChFpPVtjsvERLBnZcUrEB4mvS7Sm+KVUtrreL+nL7AZkcMklRygT1vEZc7QxB1
JFjujVPqLr3i7rdwdPKBKQbs9sxiMF7rI1nkOdA/iRlR0uOoAaAW4+zEYN6HdHfY
8GzSMK4R10d2uiUZyTEOboKJHKD5VMjuaQbcmk8wSzaqMWe56Cmhxum7rdP12Zv9
c3HWuhshRE3Wp60DRWS0Mnfx6/HVaBKmTNJKtmYy90t+0fRk5W6rNOI12e4imxII
2eRaT+8t0xAvBKRyLjWJZ5/yKxaqU+2ZO5ZMKiwCMj7xBSJhfYJs/wPb3UiLZmUn
TodA4Cmug/FZLLRECUnH339zlB3IO9TGRGaVcvWf8PhWmD0l8RMv8B6qT9G1udVh
BxJ7/wknMJJXdz1f6LtZ2YtmDPMR+HbxS6X9YFnAE4vpaxduyXT/pueX2oukSA7u
jJKkHhohOLtMSzRrYwy1yDzv/V9XRqv2to7XXYCcva/kISnZlwHGfZR5UALoiOP/
NjVGPrjvchhL3v4rM0yVcfp2bsVmYqaXs3fmm2J0+Ec0p2g8CFbomlScqtgMjhlY
7ihhSRUBl0R5sehZ3zwYuWLu8CAmp8QcFo71tqjI4bKlDkaHaeO+ZDnVJPmFJB7o
onTCG+uHyi9XYYYYVoqJjwkAwVcPSnj3e9Oflk+1oVVsE98aG9bI/+sUL0QskTWK
Vks6PdcbL33CGNTyDdv2teA8RIPiKPnZnqGQ65Uz9raXB/Yt+PNvy26PKObVfd7k
if3VbgUV6nZ1X5G1EdhOiqo/FoWp41LhQL2X2pGLFQSTFo8/aFkh1w1CbNu6opLe
zOJhBjM91ym/0zLet2rYFDdY3KWlWYhTvyrjt9XxwFx72EY2IvrGzb20FAOl3yLG
+M3xBI8KnplcnWUMXWZSTPet1r1S5jTQ0sQPrLjTMFIrRDnvYe/019LrMb16W8zR
kRUdCK75QD2hEoHsz2d3/hdwud7xyz5u/5/gCCtEoQCLuRpU7jDzm1CoiSWB6BNB
iJjcUqloPSU9esWhjbmSs1+1HjilfxYTEadX8orQJpMmgqQnWwm04IUQm2tN2x30
eGUyqs3MlRaNI7Ugjs+lMLkbfh4/+gFYgZ2qy7iFpq3hAZlaqxle9Ar7DZhOjyA3
58RFScVDR50SUxsQHwKs3gV9tUoicDTCepB7pDTG43fstqaIVJWr22rqpgog4SA6
A7YezZZf61Xizfvxbw927AFt6UXe0a4phn+toq0v6+tjouc26GisQVsUzFld5zw3
c1/p+Zal/EX8pcC8wt4HiSwI+tXklnD4aEZq8ze4SHD3d/lxKXec6h7TEXbvIGIf
Q5atSHK0kmdVZkJCsQB+Ogq8rC/UI0g+P6fvPg2wkJreUJOJDhH/OpGFpmkNPnPl
r4CKDulyitUuh199E6C6QiINs8/1wPfP+BpB3u7jpoBE8Bu33OY77xqqg+6zbkyF
k0oklstafggFHzn1VLkfJmSp8ENCUAnhUgUQVX1XELAOP0FyM7SfJxqVzawLFN9g
8u5HO/EoW5NKsPupCrsTpGjmhseSdu0pWJlkUxLiGD6ZNy/RokqDCA3tSGBisqPU
3gFI0/ykeH4B51qYpGuEtLuYb2BRKkXV2LV2Hb9/eFPH45gyqzVNeTb7FDQeogxT
8pM1xK3rWJUiG8gAA65QN0mJvjoNDJY0EJ5H8O5G835fcjOITgTmm+5cF/oGIf71
yeKOFJzDOU5H40MgIlEpPQ8cbNIX9jAdLfj6suWnDi5u8FveuuPjq0po03yozoml
Ol/LN4vkL5NbvaS7d16J/zb31N0C0aauiRh9RtKOiD07XgAWOTz3iyR6KLC542LS
3eVA7SLlPH0IG+UhwKnX/MuxUtk254DiUnDRwj1HZ0gbJnGSmYST4XDGA5tx+rcH
2hOGz1uGy1IOdPMNtIVPJLcHnaDNgeX/TSa3cDLFKu9cnY5YDY1lCJttg+t7heZQ
siHKkx8hu9tnOJBReVHWThGxyBj6wsdE8AOF4vmxzZJPn+cnYUwfTYaE/aGDfK2F
9o2rvjb7Fs9KuZvrQckDVK6z42k1oId70u+Y+oJEoYAPZ+0U+LKFxVael7b4mDSr
lGM9pkJyTpcdv5y3t/9Qi7JdEi9FfIHqRe9/jJwlGDFjHwZ4za7Qea1kLCrd2aYC
to/fb9KV7SQ5X4c3DqZcsW/y4iHgLDm386mYwy3ickTbgWhnsAuYxTmHbfZ82mSp
vvM0/Y9cxZU/9wpRyySFe0mwYFnLGjwowYFKyEXE4NGn6CGvxyz9Xhjk6XKznTHe
Cnh/NMvk817fJWsT+oxAmCqVZqmLrVMh9Ag4Ldpewg93h9qcPxVOeoXQj6aSgB6/
QMZXtoxKdNE9f4MeUShoJ8pl1obf9jd5lJCwA18Z31jVbC/88J96QFT+B8kMfpNH
bhfPsQECV0ql3n4JrlsYeK1FgZwjcw+Ek1v0cfW91aDJiMT8UH3MP+LljXHVJndO
6LABTGIkMBQE5nSR0iGNm4h616PxOdCFse/pGMHqybliVyZed4obsJieXsJunJCF
z2AT9iH/RdUFw82+JpOg3ZsTc+UH2DgnhdFkiHd6Xnb7wXHaFIkwmQQQ2T6FTvxR
FE2L3U6bXPfLfwhD3+Uq0VVDe4spdMXqfWKcdCI96qH6Q5xbIxzVQ9B5BA0OS2Mo
5AqTcyE4+G+eKO6yPGjb+Gx5zCkjNDEaT9fxuPP4v1y9smZ6hVDrgwQ58r4K7YxY
dGq1z/v0z5bI3s5jBWXVAkOyo3u3Apl30CwMGqPYZeSDiae7gmCbiDbfZAkym8sK
0bIYErH8oT76k3fu2cAKf/MPjRSxPkUIdv9sSd+WbTBXcyCnmNFzcchwQ1hCTE//
uYfd4QQmIW9j6oJnC75D9ahCcQA/5Yxu7F8tZ/lbycCUbQNAkVn0kT8P4IrzsmUw
duGr9cA/d0ZwZUZLTxg45N/LW83DEdeO9fAFWhWy4oXJDt2yM4fHCzUba1/4TUPH
koIdFFEcPNb0FIIzQmSwHUxf2OLBmuqKYAAfvoUfFl9/H/IEtRK/dffbVNNh9FAU
S+dsCJpZlFWJW+5q7Yj5vjz/IpL3UkLQaHyegWEaVZatxChU0PJltkq8ReBlGnJz
p89FC7+ZZpA7agrfBzRSviBPxmeby8wiGlbwSMi7btVd+hT51UkGyYqBtHKd3cIw
FiaAqQkGR55J/yz6AyGy1J6fQcP3LGyExchHjsXX24vqWcX2AF3Hki+/5WddqQ6D
9C5fX4DfvJHqSCG3gIbCAqka0TOghnc5yNMaG4BvxB35YwkclowLkm9u3iEc3LhO
ymc+H8bry7h1lJu0VOMGJ3ihTOCJoTUS07V5Wt/mtwRhu1EDrdO78QtJFpEII4Kd
r9dny3itROSltSxKB3mVU0YY6uWrhdbBXjKMd7hA2QC0KB4gi50pyEpEG9aYd1+r
kOxwuJquktetyhV8XLP5u+Sz3yP4BK9YP+gSgGzgIkZA0Iw0BRmiChOxnk3qNvnY
Qf3Mu+HWSpY+E8P1xYhWmdI+vIHv3C5UPn8khodXhLbtL6D+7tepfrxwlYRKxOLX
s1HHJh7xiuFo71ZdaYvsokqnwyIDa8BT4VhTMKAo3pFktFA5UA6Vb5JcqLAZvjvg
v1OLehSGWPZV+37I7Ou2st0UqtJllxQtT2eKLXP/8XQu1p5eOduH16nUKhyRx00U
LCg9sLQ+Cb18V8LGMhqR8Emqhk9mnEngMQBjB8dpQP2Ez2yJenELidO7+azw9K3o
7+WQjnUMaQr1I/4nLR/vl3xfwwmsJZaMZmzP5Ti4hdmauI8ihGjmvmVnfkoXyGxi
fom2EDhA0Yg7uFaLFZZwS2zCn0N9q13YpIc0Kucwad2Nae6NJhBYq9bUr284DFAs
XrVk9w4lX45yjQdAoIqqXc5UZYttX2r1n7fNdky0nd+a7OE7Ct26V6Vjutf5jcfH
W26Szc4OGB9ljgaKso9qjmrrsyPCrWmTepWm6fGOl7HtUlJL4kRBk/VEgYTQD0TA
dWwAGUE75TMn9CllP2Fopz7fg6/500sfe4BkXcm1HDV8nMazmtyfiOFrSL8od5L9
SWnIKtexUgZCeHzuTe6bXoJjV4JxHQFpwu3g/YPIQnCfESpuw+vTVEuAF+03tXJn
lnmL2XxU1S2C7ZTtSQ4Df4PFfFhMU4VNVSlcT6Tye0P/tlUnhN1Ms2RA4UGs76ud
Vg3mgdTmFjsVQ5N1BDQnyoqs4XqvG1lgHmyQBcm55tb1mE8YJH+FfxW/b2+dOE1K
w7JIv5V1am70prAHrlO5rwB0Olj/QVKiIlAEejKZ/b+9H1LcbV6KhboU8+m0av9C
bG808pWsZb1r6XWiEJdkF7Oc6XXUoEqwjqEM5aTqsQFQBam52pFL9Fwome0rWDSp
j1/9nPp5JK7XIivoAlfwmUgzBq+bg9Kk5P7hbid8uG+DQkLY1R2D396v0QjHM0PE
2mNkw9NToLLdM6znytQOXgXZeDGfjkJoaG7FA/49DQSDEP+sQk0eVu/0Vl0/2wTB
QVF2/ER2upRkxEcepYqEUxRkEbWiZ8VV6N+Lk7OYXNVoLB+ArKQh8tCtF4k3FFfI
TO1NxEyXjK8x7mlOuTF8Fo0Qu7wndAPtebMPkSJCSz8E0ECDnCDfFjHs1ofSb+Wu
WzUikE0RxXpwVpQtRcG5v8zDZsCXAf2lR9AsTI6i190NcVCG7dV5t5Hiat1VOpy5
OHqdHTOyqynJunyxt+0v1YshPg6u7qagGZaAQBelIRp+FP8ieog86S3Kid/W08Zv
qQdhLSFq2nWSLgL4dAp1mnY1zJE/qoGpCGxncNAT1JnMvDNOUedKF8d84O4QOkKu
`protect END_PROTECTED
