`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LJboqeh1Y3VBjX3L2aUzTcqYwIRNRKki+dtdvzbg9LeC9n9pNwIKkt3r0Zr9ciFI
EGF54zswOlrh10Yor5zvfUtnkEdC7YCLH0WQFxg15+INKadKj1DMBMce5cWxrm2U
amWnws0w9ta8hWFzMjdehW13jjXRIeRXnRRddL3cEXU4xhyfWNoDnTFPNONg1Lk0
R4wqLknUgSS/peyWQrABWMW+LC8xbJLemzZQKjsYFyVzFgKanNl43Anye6mfxKzQ
WuuqYDqJ4ieuy97A0lRBreLHvJdxfWak51jsW8+qNN2mK1mGAQ9pTsSkuxl6WaZO
14Yy7bUbrBlQjyIkXgzSNlvd0GP3nDQyh3fpaCAsmrMfkHaUs+7mXUlZLww6GisC
c4wi6+ga+MqAOD+8QGj7rGEKlVEOGJKrxmrr0wV4u6VDiyZCLerKHfnh9lCxKt14
ZTUfQm9Qot6qGT9HRg5tK1Sv4qCHmq8qr+XPNIUThDImyDZs+Btz+tfgEMpIHLMp
HXYxTsh9lEEnzRB1NsacOPZr4UAJnIE/qkBpA6QhO8lPE6AO8OhRAqP6K8rkpBj5
5YtEqAOKBe0JnkeWab2ka7lbowrCp2gkAx1eAg6/WXpmpxcR+PJVqkSNUE22EOG0
rdXkepp7jSqvT0rD5ocfbTKmM7ekLZq+0xTtRJ63yBjlVhVlsesZOp9VEH4IB3z0
iZRW5+OvpONEy35NG7rKNXvzgeQsQ5DgdKeookeNYzRiYmMhZbtC1OdQrEHgSIMS
5xb/l4LLFkMlE8d2ss9fCJwT1mj/NY8lQ0zHvQ5BiQq7eLvK+gWY/DCq4uVpMA66
jWVJ5+ZwW+qPw9J8q5rAKsvbCeKgPIE8wLIuC3l705eurH9NMXVhzY/lOOiYmX7R
2wjZls8MITeyqKQKDqBTqlXowKTrfE3uY5f/B86e9vaNEJIpAi5qAvYaUybj4b7z
Po8ioB4kjkZUoT+JbQh/oVmjV0ZZTq6aXSxPXF27/YB8fqZ+L3daH5TbIsw7yj1O
AS47AibV3GxqfWKzFyqzg5DL8wKzHevCxW1IP4/2EpDvuXWaGT3KA232/VEyF9gu
5AcfB5PsvyKqAcbT3iKZTxUB8Mh3HGWYqo1Lb4uDfbnP75VG1maTUjLDqjVwV5y8
TCLYurpMBCRtebnk85jBwmvQswGffn9qk8k4BoRoJs3dxhEw0RF8A7Wa3Shz2QdJ
uBpFJTmgFdPF+sf6j2TgiWeICWFBZYL2G81qlgf3NbPur+wPMi7MdjpyeD48YJ2D
k1+OfSiUtGzvVjttEqzaafUNix3hOyEQJ4P82HG+9D8bQa4PJE5FbN3OT8cpOzT/
IWUxMLErlJaYsxUSSu1q289ZfZKDq2PW0aFgm1Ty0Yj9inmD16jBnAGqJEl1Q1gI
fDgHCo0dVwYDAKDwChcfd3wy1M+7XQIEjwzRJuR4XOzO3s0P0r2joqQtYn1+kVHQ
s1ogMRx2qkjv4mimzfjk6Sq1PWE0hR7o5fyb2+jH5lK03iSJc1RjaagepMX82BgL
ku0S390WI7jLs+HxIyNO3kUNYE3PIAvW0n18tgjudP0spR0TuX4p/sNiKm86zAGz
Eiu4jwRw8DTJz0wH2t2fXKPR7kbQWwdkBycNqboQhBy8GRG4LaQzDsLbRfKNFdLq
iQzqo18BLw85SNGaWmVOvjTYXAjZtiwkMKU4vEKw++9pZI+YGwZ8F2GBgMoxuJ0O
5HgsDvCfVmnN7K/6Vv1DSI14nTlEhFyD5BvBlMlir9s=
`protect END_PROTECTED
