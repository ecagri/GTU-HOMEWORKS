`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8RGvtFgh2UMpczy+sMauTHMgAEMh0qMOFDO+RnwETsl2TcNQyeTF+hZEn5BLeh5q
Con6m+UUtkVsaDzKZppj8KbNi8U5l5B6vI5b1xqBkIUERN0UZeREweG7SBnW65FT
aScPS7tnpRvy463SS4DYJ9Lvv2a1fmIL1PTNT3+psypq6enaC55tBsVxkYojx3sh
fNfJYZ79CCCC+s0AkEedQ3HMS9qSB52Opt3ZdjW7UBoRw3mExpfOPlc9abve/9XC
isB8EjaTASldnAqqgNWTne67dQZwdPKON0SVZ+9zSFhvb5nzk4LiYdH39ehko4Jr
lQHANRNMWVqNBjqdIykCsTVyUok9l24ylFLTe3FWlXWBqp1DpdeDJAWRB3mDbCrn
jh46MWHbzsVpPG73wwFUOQIRNtwT0B4Bm1UCfGx6lLKZYsL8thCfiPmfuU7QtPX4
2c+/wJRMyvsykEW2Ecwz7QJBQLUqKX6s6WgbsOzF/QQ=
`protect END_PROTECTED
