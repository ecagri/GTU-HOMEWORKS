`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
33PqaCTEElMHLfzWLpSnxj/HHyhzPd82AVhiypfx+hjFoDhMQvGjnEbtonFzw9Wi
Mu37TwAfP5UVn+kVRGfM6Jyx8g+oCZA+3BEmeX2p5wflJcwFU9lQt6Dg7TJ250sH
U9r/UR0/VZYGwMfqv4Hfs+3p6fksi4FqzH2VlPHd3t6mvPmpWvABWaNl3iyRn6X9
jaL+isK1/285kSvMu9st+Zwl7r7D7reHergEgS7nOzQSOt2c4iePXOuBXZNbbk21
rDA2/RFlI3mZ5qPOJ/HtrUFQZwj3/OodXIv+87PAmf2YhMCaApwgbFk0nn4GPJSa
jnAMa2LV/FYSmO7MMMNU4tudoDt0SsVsi/hXRgLkOt0EPknvYfcUjrHDQvp0OIJW
EGCuhzoK98CpuIrzK9jkuAH0AvS2XwdvgvewFrxxtDJ1bjeqfqGJFnkOARjfDett
plxeZrWWeWzQk+StaPyB0IvL4R4AC7eD1O7d+QSGJOPiCdYe9/ZR9bXO3SObraqc
5PT16ceu1EkQEc0zi3efzL6awFojNxXz3d8mgU8asekCtQpxNkaMy2vd43Mh0saN
tb7RZXQooTEYmhSJEo6Tv/H5tG3yPLY68QfgBJrjtVkuuPnKTgacTZXpYSvuqZSe
kxRJEhZ9JYN9+O2kz1xRCFQWybZwMjO4wfH7NwEkr8UrzB1mgDRjTn3ItjRQYZmp
6q9K9RdGGh1eic7iwC6V3qEPF8PHWimk1yTxXW0UHLlvprVIHocoCk+/aJpebKAd
vBi/vS5ORtOZ30FI/IYC8sNyODOaurhefGbhoweflIvWfvYBHYAdyBInAS60ee2G
dBPj0zAfKa6isFVVc4O2HhufzoNSouDCjFG6U/MsrfwJFnnqeiembiPrEb+4VLvI
4+/CGZ1DhDoKMhsfsEvzzrZ3jCfD8/hdmYRlRFlj8oTps1yBQyE9DtGN6SZO2bqi
VW+h0Yqn8+xoDadu1ErCHxjfYNUcYx1yQiVrKgNIiquQY8c4RqSRM9DA0/Fx0cvA
TgrTLt4CgOwE5P85jQz/KUmOwcWv4THYIi5OF4FkpbIfw1dCOjDk4k81i+Fqd0Jy
ryMll6o3IvM2LczWboDJDfUIf0eUbv2Ajhmzx3RQnF2JlEgXsVI9MMLj9ymnWT39
QMNE61a/ZVmv1UUvNJOw92fbGOdhb5bD7iSKaeaAFhQg/D+PvwXPLJYayDx7PaLM
9qyD6IPPWbuY1xidap5XJKKSbWwz3NN5diVmvKVDeCb5Hm1c70rUGLGhqa9fNGyC
1JcseXnQqjMV8F51ceEyyXSX26iskbgqKk4OfitIe5IzpaHyD9kzWFwXijrXHjof
ZRnp+B1GoXJFSCUzJMtr8NiRpqYQ+5oikZhG3QCuN8B0kkN6MeUEAZCY+dWqde2v
Z2yHuq5luwiBN8xkHGg0symXt6cBX4icP465GW1COg3aNcog8BRcT2xOhp23GD+P
cx15z7kYhl+LoNbWNf3HCwtjypjNASJUf/cRB7GapRh8W6+SJDw3kSW4H82TGu5H
0VpYVCOIIJRwOg6Glbudcw==
`protect END_PROTECTED
