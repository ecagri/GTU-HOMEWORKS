`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uupsVdJ/syrlKjWkE+lbW1F1MunSuYSkQU+5tKSGS3X9K6VRikty8l6H05Q0rxAd
JXmp4j4P14smPESKcDDSmPc1PKbb/8W1JmO/gWoP9r/NF7hiSzpNYbi76Ef+VoGp
AiNM/iMc1IAa4Ek3+uT1MUG6vt44P1YWdPjQJlt2Avyfyj+7BlW2qC4XcpAJ/Ipr
vdryqnXj3atJe3I5/IQ0klqTudA7EwXLIUj4Sb1WlKmGT6IOnaWGIqKmSTBAbuHr
fxpJq5aoyvQzjknPL2FeV6MiGWzOKZ6DO1wUnENjh6qTAVdsXgwmYHPPeTnzkTUL
H3+kcDh2r4qMXt0jKqAVdWrq0IV3wqbqTzIEYxpdG4aTW/g3vcEc99DHQw9Am9ez
h0MQmRIHyBZup2CZjkF/e3TprmtdPqkAGZ+EDAsPaJ154zEo4js3GsZU9zZSd+rO
P5xvXRWffLohccQjBd7LCvgnV0yLQqsHD1StxBiNX0ozHbMUn6tdFIOcdH9vFrKw
q7oU0ErvycEnwGFPUJvNaKJ3Hni/RkIquyIYQ+hYIbtKO4NEZhpxk35QSZzfEmqt
viqWVRP+tmldadgHL7D4dPntFD/aFcDbB/57Akw17J/SWD/BLrqyHSC89he1NwJv
jdbryrvRgribooJKKgRkbwMOyF+s0HBPBLyTrLL9meTpswOFtZD8Dd05Xm1dEjiB
iOvSlcB3vl6f8aVP0LufnoAlfoi8pwfEw+073gFahD5Rcnj9m/U0GwVGt7r+zvqQ
x2uFhkeUF7BXuABlUgqzinVWc5dt4zwC9Zy+yPnzEMSS3rqhIvzGU2miFoy8I0lN
xaln/LQZP5wPH9UtAEBR92lOmhCXQSj2B8NXKeHPSEz5B/Su5OtY9qziVI9kz8Wp
BRTNT87/pNpa8aaJsEGTIwEhOz3pvf61VdHj7ExM4LL3C9U3T+kA+Pz1fHA8NqhR
QN4h93mfR/rKKIoN9Y569AcrE5xfK8vqpGkVOpffQFMzvu0/TDVM2+1y42t2Fl9H
61a+NCfYTlR56KME2QC+xOVhtbTNVOcN8SK9yJP4rkcB0TEeh3MYjOQk5R82B3mp
ZanEZynK1NoBsVngLHPdNgCwXJcQxJK+VYTYJ61AXnamB9JDVqHyVdT/LOLQAlSC
SsDlvg34vplV6fpjf1eG8aJSHLTSaY244OX1dKGjMOiojeKCN+ypf9UIApWKrmoZ
bRODq0Ud4GU6ge/S0Wc8HDK7xi300OgP3Rg0YS/gPKlCOYGScEDMZEQjWsQv4SEV
RZUa3Ob+pDjm69cliWLiuEpwT/RWtY7ofb9Y8i7Xm+oB7B5dUoJSvqNgJUNVAW58
Z5Tlov7GtqOxU4/lDiIrqg5kPFdgqeb0J+OQGNS7Hpoijg6GLF/9BAMPZlx0nVQE
vhWs7xTIKlhlwztF3jvdpGC0FXZdV4K6DItsFMrWPUm3K+KiQqw2tRaXGsRYe9+H
87t5CacU5fg7ThLqBEC0K4Nsrj1vq4URmV/76sgb5UYCJNM5h+tN+xMylbLxllWG
IRaHheK4W9Cy9wI324hsmosDzx9Q2pteLj0AQEFUc2gBI9jQJNdNG0a6VXNln5h0
1Q9OlMmtJC8iPBFmUohGduqgRm0mUWLdT10YOgGKBuTdLsd8MylrAr56hErOdZTg
I+Hz9J7VwUig4Z3AQTsyiebxtXBX2hKk+5QAL5OXFZRN01gb9VNIBw/DCcAe78dB
D1BjpyHIWUMavhDiU7ltPpNik8fXcJyU0WuYB6sy56qZZwzc/sI+wM0EvPC5+RSw
ZArRLTZOsT01i2LcSvSwSkGGYmqq/5LZj/1TZE426zMzZvgKKcwOOhNTAs6SpB/3
XEJI/vf5iqkedzbqcmDwKCTraPWYeS+wcIfrQ2Pq5Nrh8hMFLUtJLPjkUOSTIDq1
xVjeYfQyv/1oUyRNwB2h/Jw0RLgHJrNz2hcSNSNN1XD/0MQxP6HOQXoxWGWQ2K1b
KIrxRF+jOYrRUXejp4YNLyLTKgpRVqAv9QPtuEc2ivcI4vQkcQ0Z33FiY+nyObmQ
MUETNhwBoHCs9QYisd0B0LeMBl6mj5OvylyAXzIpIgSnc4Pl5sqB+R2hvGRUyVBv
bqFoQJlhYWpQMrOBmYd6L8p4MpHOfItLvggUupm2C/AiSTKOdLZfkSGm0hqSEnvR
mfrhztJoIa5v+hNChP38xMXH+hqNQrfS/1Xrdrwgast82m4x1M/995kvVHcZ/uWo
TXRLSxaDQL3jrE1QzRgnPDKB1yyR2gW4EK77Ny0RDJtm0QkCjIheo4X/04p6xXFo
V94wlYgvWLyHtb97i7XOcDmQnnv0BPXSyUT/UD68mbVrdj4fdf4udzdeG/6IC2rU
8ZtWSB9n5Ba6pETdkDVHhtkhvThrc1ipFLIlzTuO26sLJQS+u7KwdlWk/RhkDCd/
NnlrQaFScJCftmEVJsYzfvhg63Cvv3URFCsQDEHY834dwNaV5it7k/jON4vXnEVr
mvdSvA9IqKlK90vYt4EKhA==
`protect END_PROTECTED
