`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gQh5HXEMvwUE/DvybnPRf/ghpR9P7eeXztyR+J+ORd86byct3OE3kq8OgWoPnun9
7913XFRG0aP6el80lziCe9UqYAxbLzzLIEU8ZgW+sgJ4EbKxXWQTtFoIKzbl4e9p
R5cj3ledtJlMIj3FT1B6hRNzZfuBy8I/pbGFKd4fb+99RLRQqLPSnHYeBA8Etz1x
vCIOqSVbezdq+9myLHFC9WFg7Clq55ZzUNW19fA+QJxB1GBEQuH0mbh5kR263MO8
HfLgzYT2jQiJMoHzSX48Z3CQxSfwpL93G8edfRUkg0d5vUZLBRuIIx0QkjDDuPf6
1oR6HUo4/adL3ppoWcxDWCH8ufsSbT6uPO1YKrdJAVA=
`protect END_PROTECTED
