`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IGzvDc/9jvRs7rq+SDjLYuhQdRAGDbLxuLvvhrPNJWyqJdnOXa2QzYwxFHwYWQu+
KMBG7Zi+pmUuc3h//1qnMF8lp22KNxHJJzEZXLS+9PVC6Pb+bpVCM+p/e20AwCGW
/zeFQepTnXz6282bpZ4K4OtzWuiESz30IfTQh1W4eyctpuCZ0caRxYPaND7YOe2R
+DXqVNe+ig9QAcGhbhY0Yo2aTqz+KvJAt3teMGXeMvvaSWR4XLtDyeI5PTc8L+H/
fr+09nHRAAekaa1ntJ3/VWJGOg6jiBX0F40W0F4oMpNL7aC9E7cyUJd/sO5fEyt0
EiMXEWiNZ7SBhujBlNWXIbaM2S5VghPFsaAiZ6BIcbD6OttEwvKQxsLgc0VJwqq3
mQpb1chfWHOFXgou9lwRVF8A0chN2PvI6EXlPcxL/umAEEABpOTo1GWR1RuGOetr
qNhEV9ywQ7pGOaXGyPYPGrW2HCB5T2Q4vizH/+irU83yPzA9IGCvBHtbCd1rM11m
cfqEw7f66II39HpuwSd6HoGlwTmHK3lE65etWvNPr0uTDgbWN3R5XWKiQtK8aTBp
Wr4fhbUvlJFM8/JyASJukKfE5zsG2rBEl89zEjT6L9hEZF4bA3X8mpGhg5m8tTIz
yrc6fd0UEgwH4IPjZL1Y1kSSPZAb2GMvrTX5ns1D/LpzBnJSkMU6zYC/w9fbFY4+
VGzC+aiNdw297cSWNH2M7Qsusa/Ng2crDcnjmgFGuOCrenqWkumcHAz8lJ5VBdAf
XcStntg6SCZ9DQrPVHyDsuxTq+w9PxLYPuEPUc48J31Q6dwqc4OCtAs4MyXpFGHi
/ec8It2i0v+CrrlPo7XQ70Uw6DRts8Lp3ySelwPohJw=
`protect END_PROTECTED
