`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kJwqTqNzHFYweBMOPecRiXbkQwxbq9Wv1K+MFBe0g6JhOH9uYpx47qIbdosR/Bq6
P9+yjZKCH3No+it3aUZbMzIanGBmpoS30OU2V2uqqm+1zwlZb2/X6XTWuJiha3oQ
DEj+6B+Lv4VFCN2KwuAXdyeSE3TvRoI21VfS78F23FV9+EEbOTp8HhBHCxDy9TrS
NrxfiE1qT498clPuK5wsI7VRjmHacYQSg7heZ07hopJ+I5lKjFMkcu9/zxdjI7hl
e1hr+6wDYyIJ9juDNVW0AvMz1P31EQa5Jo79KF01W8pZuk0qgav1br5d2f9i2DZV
6iuui7If/MKs/vrjJFjRtD8JEexH//oS5AdoxkKVDgYTRzEInJrJ4j4Eo0dqNnoi
Sst4XHY62hSXg7bUhCjPqRS7TJmSC7eYGswamkiEN3lXKkZ7jpXHDjqJ2/rRk0JC
JyMmwlwiVaquYoEmlcBBMPSqD55LXoaIem0Ccx43Y7BjqbvLsR9dzl1tvA3e8CGi
6n7UCK92b6aEsigSGU+IqqPb4SHzDk2++Fuk2IWq5d4=
`protect END_PROTECTED
