`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
en03lwAK7/Wn6Vzs6NScBOJ/QWngibOlVN3PA9izMwCW/1HZ4AowCMDQS9uHxWYv
NaPwI33dndkwdcSqqcW9kAm4helcRP1VxpqG68T/FgNQyfyFR51On3kUHzpIhfSd
HErCWFi9ETjIsUA7bg1G9ca+DmMBb1fa6nNSWhd1QBcrLdZKwUPJq9JJ5KUNMr5a
XTa9Nw9r8G0G5PPpgONS/8aOYafzv1KypExbRuaBiF8rcjIEvRE6UbCHoiK79ZSp
ml+5mtwj/gUNljIvUje2iKs1/1XWT3YQuiG8hkMpG22lh1WH9isFq1fVtAD6SsqO
lGS2NUfSoJZu6XBVtrd5wQ5yoyPMzHVUxT5j24S2Ea/PUHfafV+LLJJ//T9KmfEq
wX3RkgDmUFR9P8AxjQ0NoXBI56yO4iWwbkPdZVBkhVnrgErVTTmgAezj+2vPpYKM
f+IvYfUipooLMXeNqCpf8uzkV2KE2KqPmfU/vKS0KUEFrJzAl5COkpiPvy5Lsua5
CWWMhOOL6GyvjmkBSi00DiG3ODR3nRI7xOk8a4sEjT0avhXkQisy7ToaLZOBZYcF
FqNAkTpqCMHndJqlTVs3VGS2XZLjXZ1MuZ6RsDNIvzqbZJn1MdOf7mhWiBLfWnU4
5JNzQ5g7t3IEU7K4NRwOo/NXmU3uCC5Q9ex17/LGdf8jcDn+4lYcpjjcQUSzWOmV
gdorLM40xQuFa1SHKAtT7Ed2oYPjN1B/XxQSwwfxjsg9hNJ0fPvwxFsBlFC7RmWm
rj/L9yv+O/MBUd5KRCFAO2HrN78SWwBdpuW0kWt8eCW3G0fTdbrpNvnIhmPibIYr
CeXVWlz/GtlaN+bCchCkPpiL9SXhLb3+OSUba23WsrOdfORpJoDE3BVSc4JeGVbO
kyRdNBCmJsUX2vXkha5oyTnryBdJ45BiYas0H8uBmmpWIEDWwAZvzEIZtro3mPL+
O5243gcMU4NYuhit9yvFKvS9v3mjDvF/u2bZWufOh4LJOTPjCWacHv+d6GndFG23
7qizljJ4rS1BDhY9n/vPCAuzDMGi01v/TE/C5ZXyj3cOOjmcTK6UtEEQ0eHMgS13
wqfd6q1pyD5RvqfJG2hEbPtK6ltqgD+EY9xOI/7YbYigHi/NT27+ox0r91pnowAD
FiKmJqIFx8IWHyML7PneQO+PTbqDQO/OMRhZ8tbDhEVJdXP/qO66idGypj7paAs/
mEfd7MLj1hKX+5zEg0XZCg0QytyZTN8VoEWMVriMDHyR927oZuVyJqTrezqUOnUC
bQo0y+3c1a7yYpqEyjly9K5W34YT2tEKgqOFtOBxy0OgWsJ22aQH5zuyJoDDBJEO
TViHDqsSW6bAEGHQk9xr0DzoVcIGiaHd+5BXh6TsdT1q+mUn511tYiusUSllzwxX
K6ohdpj8VmRNSVC55deaoWABzpbMRUxolZR3djLc635cbq4owZkXlRBFoAiLHgW2
D79hOPJXPFQ/QbJ6wZRMgbE2pix9tY8OjSx922DaN1DK3ZqFVGds/6++UZCD7wSH
LjhMta+yLlUQLQZroxmpBKW4F0ZqyRgpGhebAYFgLPLv7rk4BF4uGHHDWp8CHKaf
w+OLNtOUvgdfX/QvK6OiA5mDPuacUIjx7YVzoJdCAeKmYMqMV3RdnoVV5lm1gD69
QAUYTsoR8HE/8z/7SXACH0fVDVgkHcDlq2Y/hZHs6BiSorubGkhuvtJ0eSTM7Dwm
OaPH5tuTT/sjgJkMm9zz+eHsoEqJ+T6LCE0HGOpc/syxtsTMLSQFRKGaEkY8xOKn
QbC274Y9hD9nhYbut3htzqge+z0yQlrP/lXWD4GuPZGdtabFA3ep4DlmQE4rCYbR
XgZHER3mW6zhV5szeJ6BWQ==
`protect END_PROTECTED
