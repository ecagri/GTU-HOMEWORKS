`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9a6FaCACrHcM6CRb477yKyKxp6zo2mslB3MQlyDac4azdfTnxjskbwmKVyiQVl6B
lMy2up7Tb2dMKICBM5sFdky/sF8zb5KysNjmoevsFiaP6AoYUVbWULuBFmbKY+Y4
goiSlLgC1doXkmY8n1LJZs+ll86lAacORpz/oWWZtTSbPjcJFBFOdBdDcLyBPk8Q
T4pmHwgLtfn5BC4beatnExdPiCYwb6O2yDJVgNg6yx3pTcfl24Gya1pbFlI0Ko5p
SLmyDum178eVqYaVmRTpwL6a3FYOBjgRq5twohJjl00oJSF31ZMKynHGO7e8DJ9e
gZqGutTPyewOIq12M8UHDx6uc4ATrWmouPqH42zliYtul8gEUokPcCRoZyUw8nf/
qCj4Gt3GfcEJQhsFtu3Mq4WccQHVR2XiUZOV+9lbLOYc1+L1RdmeFc1gzt2GcbdX
5gtoVQyfQvc4pFbJs1wTd/lSN81Rq6UFzFJoAcj1r9PEKoBmeyYqqXzckUpzwyjx
E0EMAYoNR//Bo7Q0nd7EIz1ZQysblQzNKSqrF5mmyFH/3kzz7LFA7DtFJP1QoiC8
XXe8OW5K/19BH/ezgXoolCXEqkGueFb6KJKvRVD/V/kwmNIyiSG/pMHxIB3OLSer
WcnlpoYoAm48s27XbJplh7CdftNPavzQXPvCA0ho+ZHB6g9QtxcQAjLLs2WhMAeO
i8t9MXcxauA1F5PfLf69+Z5DWarBAmmiZ6Fou2Dup9dseecE3cF+P6z8E/aA+QLl
AKSMnJRwmojK21PMmp6KLxdwlck3jR66J8k5VPNMjhO6AdU0JOpJC9YuNgHuL+p4
zz61ljyt9+4uFubx1OPgPWIPY9sDaPM7xBmJ4f1SYkMQLZPjjVcUbHdzGU+itiEf
Ff8YUfJ7mE0NWQ0ORfEDgBj7jcLZs4U2QTi+Ye7XOOU=
`protect END_PROTECTED
