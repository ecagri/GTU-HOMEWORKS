`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U1wohbSFHJT6V7S8Li5bfiSpq2n0NkRdk09wCUesZNek4Yac9W0+YcODSFY3S0Jw
D/1jTtCvudqRmKiTYLXP4ownWlpSeuWWtn7DZr5wgUejwTg+G9gWizq+iQ4hjpmf
C3IbbT/JfRZT6ikHsprzKbPtuLP4+0Fit4KJWwjqpvEoXhe+8OXrSqmg9Z/hEHBE
6Gq1rRpuYG21iCaCgdg3bqJB1kHnybmWN3ZOldzekNAwCuHrmURsyN0XFGCX+tbT
PBWedOLC/aO7HndtRLtmCnIXhmRBxvOVkjiM93nozu47+h36f/K2/WAyEZCzRNz6
DQClLfSok1YhKtcsPWlk9xeCRD7MMtW8n2IxINPw8nAbjjztnwpdBBJhmkbpNDvQ
NUwOUBykrxrTPQlJmOzYv3IqIKXcjPjHOvy/X8MuwsZFkcQyHF/CdbdK9Z1SXtrJ
78vCnhOvfN8fZEyZvJl08jnQCMUkX4jaF7kGqKfKV3WBXoKAHE2cCsFQiwrKkd0U
Do/f7mruKxTaED+T6zQn/XtL1CdKlHI5AAyY63TmobekRg9LtNwEpog6sVdjH/VZ
YxcfWwC+jWAHqb390AP+x7cykq4eBifVPJh3egpXLueS3/LTHfs1f4sXYujnJT5b
XJGRQAw+0XovmrS5fo3cV2aczCMlrKi+PQ7+wPdoy/jAmQG6WYVS7iDYU2kh6nqe
Y9fRYQwZ/xjqBOJkGGCSkXUD+ld91395ln0uP3hNQaGkpjB41lfu0O0gI5s2CWxp
WtYYO2VcyvpAYN+x8b090Q==
`protect END_PROTECTED
