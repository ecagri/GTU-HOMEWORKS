`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BJLkeQvLL6w27CNBZbQnwmW8f5J6ulC1J3bw8/qEZdxwUFkv8oWrguc9kpIEM50S
jkXO5P2Tgx/TBoXpdlvpm7Q54/feokTtHaPo1ldhUflYFcjeMpOy4A3eJFSfPfVA
tSzyOhYJiaXzjbtSS4lSD6IUgShBrFv9i+AXhOU0Hjvj7TFnvc0uDcVLEg0bTyQW
h/VLgvlsQKH+ZcTPEzTkHDEJXHR6hN36xD3zTv/1CXpEIX2Ro21uKPMFRNAb40Ei
uDwPkyUt21Q1xgIJ/en1nrW89nLhOe1Hrgnz3zp8CHiWagAmQG5OTyRPCzUPpFZb
K9xi+zirsh7FB2wOcio1SAOoZJp03wV7xo3fmRsvFbYkif5rZgtCUV/pvX4BiDGM
pYvi4+ZxfVyisuvfqhdeR/Dn6YwgKIoVCwwHVIke5yahHzdL6scF68ycRgxm7RfK
4UAyADl9fqWUnhTcb2rVbRAIzqMGuWMTZ9xxI2pY98C0H43PsSewGfScwXhgf8bX
ul0+wP6YBaMVLGvgxpIAvQOwZ86WuEn3367kKmUr9uEkJlo40m/2D1IJ7IEYQ0q4
c9uR3Kx5LBPFV1gClaOaniuEXXwgnIHqOb26JAOSq14Z2V8efptdmGzN8v0J5/LI
LPmqD+9J5LXhsDgQ1Dyp1DYixVH3vSJRqYBYmZhU1qlybIeB0PYVnWd8JUlicQq2
THQa7B5tBGjAwYmaMh6wqyTPVpdmNRUFEQl1zeA8IdZ597ksK5YL6fPUBqM76iwa
MpYJ7rIhx+YVi3EbaZZ6pNGoEcWvraAFUCZz9ZZBIIHKETvieXGJVsV+jYuUHfyS
K6zWPw3BHpwKjhisg9mvUllHevoOTgwZuWF7zdaoxzz8DloLbYBOGZNFB7lzelLD
aRS9fY3C59TMnQGlaHwLl60EKjq58j+iGWdsAQa4prBosi0Cw5x3Hx23lVnqs+e1
QzAx3zg9ORXWDa1dKHRxHmN0gy9PABPgyoGXL1A+n/NkUwdfcm5Rf6/LZlKCGNBy
lKNspJaDd+Qa/6RYOjAqXi9sXZKp9ipGdke0eE4G9+bH7oZ2Hk6uZTwBKwabSmyD
KXyDucOwnRtwpUm/bdXj/rwIHLtpFnYImH2apKlhhf8cP4nTwVPla2c8UqNa5IWq
GaVHpSqzdjrxLqb6puPvgv2sD8R0m+KOljgS7llkirTEdIZx4se0gS2famqI40RR
6eE4WROyHFxpUq1pN2gxrFV+n/csCIz3oImll9MUlgeyEaZMJjpI5hQY8usLwWhC
HA9/94VMmk+GN073QzjdeEq9unwR4KTFCfEdkxGrP8YJM2cBZAPIbxoLOz1gGwve
9rie66Rf151874yRdBvEmES+U4wD6riEn9yYdQKWcNrnG2iewMMAAzAVft25SlkW
6YhqKnFEibTsg4ksb4ZH6ZNDYEXGGWx+v6MMljHsIfQh6WrYGcF+pSsiXan1ctwe
Zb5+/jj/eWoQ02F2NJY4s5hwz11Lr4AppaJGfEjW4sihnxyhxAG3n/z0FzLZRcRn
b0kJ+Vue2a/0R6breX7ducKbvVslH1K98vYQEct0BB5NpWc5RY8B8cT1OCyJZsW3
Fb89vTMsbc2AAAiiVKvDQhwy+vpAsJi/0TKPIJg19yi8/zMn+NI+PKLWpLgJ8ces
qh45qf8ElhcHK9UMn8Jbm3z2cypBOBblUhqBE/Mm7JamxCWtJW7GYaycdPybbq+g
oAg9CylGq4pIO496Zw9dRVT1FxejE23EoLRLfnPUXqxotW8zBHz2YW8Hgv6BJ1RR
tIXxnoHfydYW9gOQiQLi/Jb9uMQjWEO2mpBtYSs0nmVQe+ql5WKLm4FNq0cu5v+c
jlgf1o4wrmW67yURDk/J1CnrnXtTpNGEfS1O2uUcVuXADvYxdM+bsQNBojeTbzms
6dNaESC9c3rFWTrFyP6xiXBFfL8g0OiiCxfE6bUsaXqRiAfwxL+VwrNk6q4qSykV
LohUwELSonuQ/wl9wYDAcym9LYxDA8ApRZgxjsYOo870ied9UMyBPd5pU1/nkGxz
Clv6xago809ne5w3aS1bYPLx6vukWyozZD1d/mazxeAUfd0YD3EjDvsjxZAiwlbI
gOjYAaToSPa8zJE/mqKGes/4j4z1kUvMJO+cxkbLsbWpSTdAIRM7XW6MmAqI6Ylg
ozpqSr+avT97v5WVdPDA+bCn5Kaxd4P88+OBGUONJfd+RrGqjastNbvL99saUycH
ghdJNajpz8ofp0T6Mq1LjR299dVF+xST28qqEEwx7EXdqqI9pRyRS11+F/0ILQyF
7+UZjv7QmyD3tmbPQdZD3+Rdvt41cye74zitddmmGP+1AXK8v7+M/8HoqtOl+lqK
DH11srji2inzNp6gWMgJXG48FyI0jgn89VQXlN2/+EL7V/xWzzhfI6Mael/f05bo
VldN6UV4I649N8yyHy+qE22/uk1LZ2onC3snblQSzZjNLbi7DXhaMBq4mETGkEvr
I6Zw6VO+8NMn9cfoIM+KBwuFCQqOpZ4h8hgxJgLL2Mo0pnAUSf1UrpwG5tQDk9A8
TTvMAteuPWKN7Icy4aXawAlgsR7hDjLa8K2wCDIh6c8pmyafW84WQbrqrQkBAOTB
5/Ba5jsG8Czatr3PJi0V8KAwA6jlvwEPPNRny+MQxPd2MubqNjr6MDsIu3ZDu2IJ
FhD/a2EeE7PL8W4ao1X4SiRAg7o0S0d+GfCFklDcEF1b2IK0qmi5mLRsaOMvl39f
EcaYL07sQikOhZPfmQE0GlGE1PDPr02TY7mzunVE4X3aNRdPOT1MvrqI/MxLw8Hb
DLQzDGRlJn+qYjZOv7h+DBbRxrz1lC3tds5Zc2h72U9tQWMhZg7/9yme1zqCCMcH
/2tOqT6tH+f6ROaSXdLz/0kJRzEuf4v168sElObj97EuW6WUgGxra0+8K87vb/mb
qm4ndtBIqYgnp0l0UQo5lO/3GH3C7HDaaDEy3G44FrZAsx9RE8cypjqpn0YwEw32
5ghBkBI/5BP3iPBjY6MzoF6DJip0DXGpJD/ZNRkaEpqZ9Z4dV6WPKP5SBr/ZUcyk
kMZQceu+e9ZWBOz9C4yIcK4Vz0ItzW60oiKxEYpxxsyVs4zM6QnI1v8wKscc0/wN
tdQT5gVRzbWmRWkSTqryPA1a+d5QlhjE1Meut+myqYpWLZmxUlQMxBIxYPeXX5yL
gLu6uIELrWDs/uSzksFcIb6VSUop3fae9kcwXLYrBa13jCdQoCs5Bl7PzQSxRGJS
7DO1mm79INKrjHZEj5WumeuVu4JO/ysy5KUG1jlg+usvLIxOSj5wf9vPq2k/FG3c
GPzMZGeiqEyWTr+Sl14UxkrBHo1ktdWm756gBPacRnh91fRzS/QmLvuyIeaRrbXr
slW8pSFKSAe1lIPj95bQO/S9TvQoJg5INf0yqIEeryccXwJSPlS6bi21ahWm3YSz
QK4WqC79n3O6+r9oZhSsa0Wh8HDDc/fmDnxx15/K4Uxch8hqFedIbtruilie1oK3
i5jwnMmEC+r3bSlZheDNa0Y4AFnH+hpraGp4++e24otgWTrpOZd8JApqWJqlvbyJ
iOikRZT5VV23KJVaAz2cAziiFAYQCbWgpkpNUsR1xQF/NTk5OCkC+UbE40GceTxK
fHPnkPd8Zl9SFngwKp+8UXQmIwRhnxU5bPKxmtRn2TuBpDYIZCkx5iGi2DQ25UDq
kUKYiZpY8gsz1H7wKFJArlcVn32SVqa/a3StA0HZaW3WwuHNsBM63J74vClpHBl9
kNuTqaFeYp/ntOMFyjw9H0biN6gXQ9hH1yrS/U0NJ9aoVwGPqNSUEQJhX3rxTblT
vlLO5jLp8GixoiEQhU7jaOvut+371sTgvm+6YxA8JnyWu+OMutcUJs/WtbyJECGT
gADUXOPqt///BPVfuqg28GgYN4eu+1MZ/YZMQBvygeulzEXBlM3LRtUC71D5lJ4w
zThojTtsRvF4pigLRs0qiOWWR56RYbMiagzwH/oheDu0taP+J5L4kAxkoy+htdHI
fx044MRQ1gVZRvdDK/oHLvpv3apv+giezY6tmGzLBKiL/akPtrPQtTtqLB6sLaRd
SVuWzkFMPCsXSutErec2FySJTqTNXfdueBxNXIplFfbZ32uOMPWzpep84T6lVju2
nbcxEZ8pY0+d6shhlXN7PPlm5Bf61xfo+WeSTkZd0CCppcLGt2PYfjWn8Rbdry49
G5YlTs4fgoAlWSjedBP4Eobghe+wOxoPdUeJWJfUlCmi4xCGEfmbjGX0kOHxIkcI
mxqJ3k7MwKtg+kmbxEeJFzkRtGOj6XNyEaqbrh05m6w/V7e5alciJpEnS/y4Aqom
hzxYrIOamLt/zs6WFxiztqne/D89NHmlPMz/r84LodRv+yjBfM+F7sfT1Z2IYu8N
q7PYPkHf9LOb3gsPTv6wUnbD2+U/utk6mCX1ltgGjJ2IVPIuknSsVCvCqrjzFlaS
Jbecc64ws5E0DRiqCSVJ6aab8aHq7DzDjutfsZBXLUzjSLv2mYvRZoC4/G2/TwjB
FJBvMEe6cCBzz6iG71CeifkqmXntiHx/awvHAyyl7HQGr8N65HS1jDRGZ9ETTcxH
OrqSSZUKvONuu+u2y1KdLIr94WzxkO81boOSgtD3H1CoYkZ3FNj79000y+KGvVFk
YLDuUDhcg2Bx+5NaQYl3wjKCxizl0ynA2xe/HtDB7Jz+vqbqac0nG1xS4sljDFUS
VxZYxCSX3cNxJO+JXl7vy/fAjn11BqAd12CqSwFKjSajLYnDszXpScg+b/l/JiC4
s2XqwzVzDDoC69sbTqah8qxzLqpg//GYADhKIdloMP+Ds9FrmBWDkhqEPHzlIBXK
mNz6b2YmJBj8xfU3jNJRxvl9bJlNNaqbuCSKkdLsKylG6IR/QmaR0wbwYAwA5kBF
nQ8dN9d+TdrGAVgkAc/sP3dkg3TvuZ7nWLUDT3S/GVPKAuJFPq6kIoyo6I8vfNsu
mfSYUQQff6jOZMaGb2MGafkrwP4vSxvaXts0gIc09UnNCotp/5ssHCuMRVDFNaL+
pht/RTTOMiLEMkOwMVhlHWCMwYCOAPB7YvT5UucYuFrX93V9QCeePaND++xEBz0H
scfulT8C38uMx2aMsqyjOY4xJs/Hsp88j+QTDRV+VWIKrYXWiqz3AwDclxYbaB7x
KeTfGF4K3Iza2P5kaksLvDjRqSy2V4lwifqitjDPzhBk/MIQ/2pZWGfDSl4LF30Q
hZmz3uD53Jn+S30BxtzPJ2J/X6rucfFkAW4YuRUrJ4dViDvTCoMmvbtUZVKd0ZEg
1NvFFQ/IYHEE2yZof+lddBq50LqwGDzA3i8ikEUNt8P7qlKcsNUDSNZg2VbsiGI0
6Wamo4zIeAqhQWt3knXb0mN+l/g+D6qm5TS1hTyetDPHSotDh46moznEMShdj330
EIIWfqOtbXuuD0k+60OP/0pWl6nLVRaVGT1fr3hgtnuWXgn611Jx8bMrCMyLDQjr
JXEHcO9kWBSfTuSfwEIEly3cPX/D9TGURJc629gquMF0tm4x4nXZP9y+NIQ4IJUq
L0NfOA/tRn+KxO5IZcxvZ/uz8cIpIVv5aZaOtXXXJl1SfUct4/XOscGXkC4fwb0+
0kC6EEmNGFXu2GbTB+gMplLDYPJxaoux1a4YH6Yr5AbHXpqjt/GPOoSNqvG7arQA
RAg+MO8H92DYozcFyCRpUIYmVsQj3W5YJzujqM/Em1I9IEI4n2qijFyFm9x+KYbb
VWmsBtis1q7ElK5ELbD4sGHyFDvhqv5VvSgeWH3Kjia+dXPuuyjfAl8RNScm6QVZ
48QIUUc/9omxX76XyKDkP4Fz2UJNBc88t7ZGm7y0YLFEpRu+RtU8ysNiAZS/gmJS
9uJzIsvAMtLrOIRs72CjTlyzrIQk4tYtxEq/u9cZKgz8eQeOwIjAIwYgIz0+J/at
wzPXWzkquUHW6BpLJ6Al6HpbRXJGyE+gErJw0npAajvzhAO7Oo8toA5ZfWHyOiMl
qiCLAwzNa4fRqn6+gklBESExLmk67p43cRw3yCGHZSJIq1dsOdLRn73yJ/5fOdW8
foYs92migvcAzwzuNwEqgjWUfapxbtKSmpCqU0h9gjm30lzZLth6CLsbMChh5wKM
ggd5AukngIwyqsO5YXOy1YPmnlz9aCg3AzFhNp8z0F+39Xaxa88t7AKCk2KdWt+h
TbemY5A9xunsTxUkDr0Vr8hh669qVQBCSC8ZDddMKD2hAnDcK5kH8HP1zIFrzCpU
FhRx4mnTgAfWd8+pOO3v7aSlaCZTt2V0HrEFE8WFKoNuU4FxkqcMJGexAPOcIOl+
aPjmXs7r8FMHkHpXzkL0WFk2UCNJF7nJ1IERC8D/LqAMybp85L3llH7BLqXdL+Zd
/cw1vLc8iJa+975Y/mclMMnxjuf8kAB/tuZR9SZBl2+CJh9B7Xj0eYi0VcsBz79g
mtFMbCKJRyg3KeTTHHMB+3tbM2Aw5QEy19MKq4slx26oRvj+1zw9RrPX19HmCG4j
MRBX/J8OMb53iagDee54iIhFS7IpdjNdxFLECpvroW/wwG+fAproJRaOqUNRZUmJ
juk9aVJQ3BdaLPyi7i0u039XvhdfTgPC+vl2SPJVQBpZpkEfA6nXYxcOab/J0HQb
xDXAr8it9KQyvyIALSa3q126WZE19/vKybT7wahqtuY752UtBZN57atiJubrtW60
FEgKXKWKJVkuNRe8SVqLp4HxBKuO9HrEHxaLdoaOAv9ZI53rCIHwHtxOMD3VwZiA
VN+lk9nMQQUxnxCqCc+Pa1/9E3XnUvG1CUyddyhtDXN+Wq8xW+VeauDv/7gRpJ0X
1AtUDjzA5fY3diR1pvrZCF38yBoK2yKB3sg47RDmLZlqiXNbXqK8oWVY71KjqNFB
niX7lQHJG8j5B2dAr3bSYG8pMDn+wsJIPVMhgklEhQxKsMsdifmy4iQKC2na55YT
s/88z9uIreC6f7IbL6kbpYxsSGZuVJfLr1szpuU0tf1khMOJdp0vMhYSWi+NXe0f
yO9v95fAs9O0yIZcSUKb0qS9LTOI6BbiaSEfJlV0YDqKRg4yiJGjedVMEsu+xeIs
apcJ2CUDv5CtBkIDkAir7BXh5m+QZum5n+896RE/3IelVvic7WhKJlrNnLz6Qn9O
s6ojOIAq8gqx93Ibgj1GRgWc4zLhc31kriISPfaPpyvuLYcJCHzHIJGUnYUUcmR+
P3IPnkOAcl5PZhhwiGJxqz2RV6v3iDXUbmzrE27VAWIcxl3s9e9fii4JZqRuLJbd
BCzkUro1BVOJ4+MlIOn4t9t495pVDl6+sVLjNw7FCV3jlqRZi/Voap9j+IB60D4d
t+ML86xh5cyF/f6j3r0AHtqb74o3orIrZRLZOZSus7DKhJ+TSByclgHzBsEB/L+I
Py03HPs8uIGloHHU9XLc7i1Q7zwppuRC855AoZci0HcUzEpXFxX5rwNbIiGkIsV+
2PkNyJBrEdmVXBdSsAd/NUtkKBY7oJI1Vu2JrFX2NgycqmkigOQvqlEg1OraL08N
OvFjmNYwVopApIfJVhrLkhCgASazyvvQ2LFPFpBvu0jThyQZgSZv2Ii6cnB8uALy
FZB/o0c+ytZd8+SgEaUWrXORs0R/F+Yp33CLZ4lmUV+PqjkVlovefdacocGXXveD
lmmO1fnt+q9pLVlBCMk2wo7ZaRjEPiDVObOZ71QXvUQ0Uec2IanDmkzCXzGA8DnE
0+HYRvoetvzuEEQMRAzHNsx67/fcdiny/CmN/eLrZ0qabGC60xqfw4Scpi9DgBpt
28OYGVf52xkTmT2cC1yAi6Q40FMsjBCB7Q1yzmvAs5dUXfIMadU2IJhgvv+yZOTy
teFN+ZK0Lr8fB/pVvxnw+8ETwZ6U1o1oXsYxPGC+4D5sRW5w8JLIsRtKlee6mWkC
NXbWQfWvrqS4av601duHd/o5yl7a6It5BkpRtqyEWN9kZ42PPIkTmPdPiyP5prN9
FVYeCBMyMR1cdb4kmbqOqe5qI7GoWzRBJVL9d2i3BQMKblR8aBGXw7v9HScxRwUn
2Rpjc4TxTEQd8FWMcjWc+l4SuqqCXtdEGMdq+0+yYeN2MLiTnpUlYWZHGzQLwjwY
t2gd6UO+p4fzP0L4pjfDqyB0HQJI4u1rzeGHEbryFdWYe/igIkVHdrhbXjpjGETY
cmW/TrB+uR/2neIIh5S2JngdRXAZigfHrFapZsoPpz4IeIEbjJgJ9kL7P+j/PCTd
Io8HHxB8ehLHxrvlqdCoXRMhIBt3bkR7yC9NSeEGcm72AuyL9ECaZV4FfGJLDucn
WLwVVCTL3AO2DbF/1jgonpstasfN4P2RotoXHQDoIEAXnDKyvRidEqiv3MgVH1sB
P7V4BR+dS6Alqgi1p0i6UULbz3KjSqt2aKbeZbgAhaidyaiqosmiZF4yF8V4Z0H9
fZSsQtuNUh0K7ZwoMsRYzPHKaYFAOiJl11fBgHvbe3j3r9r0XDTCgo+KlmIvd1uN
ZxCqbnoYfEtMdJEME5/Ej/JYPTAJtRyDb4Zn/KNQYvTBSt1wpIhYJ9eq96eHak9I
I0euHn3J7v8OFk2L/2FSUFhQPvXZozCCoTim2jaHrtFkCYu2HQcuzGKrWTNKuIV/
X728WILqqD9XbReoqG0XNWPluNG6qCQfxtGJB6Ctp8SjUka0G8VogRqtGlFtO3qy
45gBEaFyKEbnQjd0k8tSE9EU+ALAgUSBvfVn3BnnzxmPXLUeN4pBrbVWhcz+LR2l
XQePeN8AHP05lwoFM3KEx9XBPiWVJR7vfjvOAIHY+Uw/jHoKd5OKt2XTXkXsRIoE
NgyHGXIRQLwqbmUzPO9vrU6yYkD/TOx7f4dXrceJAkMVMU6sE1dyByakHs9s+M/X
E1TpqeR3H4bGED4BkAExzrbVBGxYsKW2tR9Ms9l45zHjO1IaH3VRSJrjl8Ebbei3
euAR77Q2xY2+DA1h/PLah9aXsrHFAFHzLSiGujLorZRnHInuwlQuXv2N+IfrcKXY
VBPpI9xcRXL2rQtvDDaFAGf7N55t/D1xexbUpW0sGxtCDVDROiQR5Sdt5ZPpe6y1
wMod56BvJbTD4GVU5FZY4vYmyxVFursrvJsj9AEDpIa46urF611APwlClJYPAD0H
pL+bvPC5ZWPr0JjK7y6piq9AbkigngQvuUidibAoCvKNNT5bufjGfQqqyxZR3nCE
1JyakIPcc9qL5Duw1dN3a75bHjM3j1In9LQx038HBZ8tvA6jAXpgHUD9DgY7ppuV
qm1C9haMNafs3bP/jh4V2a7mf4Bf6s2Zio2Dqufz3Ecv8K+7VBo8/7/0EPxkEKUW
swqewdiGFCP1BK0ek+n7rbTgRSKEbTtZ2Sz6LXqNIwvnTa2fuDk0rL6yrwS+cS5C
5U4EicdUIbaLIBlEozs9ocJX1kBIWK/Iey7RNePMGIsxuQ625MM2uL6N7yw2GdRd
/xTvcp+nTTgqjWmLizi17LigrjqKunEGbb1lNSEO0KCx5SP1ybgopZAD951mE6cs
4nCHo5O7ryRLQtqZwoI/ELxKCybF/CFr5pLXeXvk6lX0I8AUflXoyxcyvjIhs0Ma
Kykn9jPdYDdVHkQrKFZfIjtaSs0/F6oZ3jTKXdRxQi9AwbX3vtMHBbCY+93Y6nj9
WbLgzyY3NX+p/O2OiJa7U9AO3FZfzRTgghubW8ZiLRvesJ/QtWCkS3T7I2mUGP58
CcIRAmq6j6rQqN0OZxVTS0gCsps6QQ2eLFGj1i160TMIwCx3sPXIU3rk/Wj87n+z
h+kirLfDfJx6xngTOz+JNFYxRBXC3edOdNGXmMNdDK4=
`protect END_PROTECTED
