`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J3Fus2OaITCLtoO+EumghcktZ7Z+vekX3+TZu0AUCbBD4EBcqA4BuT28NqyFCGm8
AhTpbbG370YPhNZS5UsuODtqLYWsgjTX8ERfoApIGZpoxhZZCstIw6zFtH1udWn3
drSC8f22tdMZDQjRYuIiKRv62qTEV3m2lXt8IRzXk6tXxIJ/hBTaRPYUtb/8nCt5
qDDDdgo4nRgg+IptOXK2flK8gZuycZFq80JHIZX5jDtSq0Kizn2waP6A91OqZOB3
u90CwSMEG6ok6xVb/at3S79OLd84fUCb23c2xr/MIEDHm3+/WGTRQ+uWgbzRz52p
I+Koa2NCYbNb7tuBGcsKZv2p3B9YLSWoJv00hpin5Lgg7pUMjzuyRHGF1MTcKb42
PGkCMZMsBTIj7svax20Uyg3NEpvS/o74XFGsdsEuYcr+619RnjHZrUBzsUzgdvJ/
4SZUx9WV0qDXE/+3NGPNOEFLKQnpJdy/+7HtA0Vz7nobor67wGKJbmW2iRLiY2yM
wD/TiVSs2LChngLIgliACdHDAHtrJVbEheeiSBAQWrlGoD+ZhUh6BAIXwUeDQ0SK
OI+VqjpUNwe/vE1x5ZFQoYTysPIFUEdpZPJWcvzgkovBU8DS0We+tFKsIXdaWe/7
+ZTEMTyLyhK0zEqAISn+2DQtJCpjc149TEMdoqQW+LG7YiNzISiMutIFZ6tj2krl
a6DwG4jDYxfvvgfRHSw6IsNcDcm7GC38z9Ic8IbpHStCAeE/2dJ+i0Wf7AWNKLRA
piAgzD9mowJufC0afFbwpg4BhWSAflSmOYYdaXmrKPG+MuA2vT5uTAebkc7rxshw
U21G8+a+30mF8i6ikptQsGt8pcFUwWhJJokO4LZW3gMuv1jjHcX5EO31N3Ea7puO
HL2bcgeHL/W35V/4OcDy4Sg+PqdpRrR99uTEtJY03SuT34QRvShqzjMA/GQ1jOYj
`protect END_PROTECTED
