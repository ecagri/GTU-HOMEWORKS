`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U40rHrRCi5trCATMS5IYEkolnVElmlM0R8mSYvo6l3efQBbRbShzpNCLuGiMs8nn
Db/4oDjWw5SHqnaBmaaT7SwHtnHyXKVlsu4/eeGz94ozLhp2vXEQsednmi8g+eZk
KztrubrcWdne247zpDHFgrK4c7kpmU5RzYE+TRwjRrvdFHsVgl+FF45PY5+S5j6j
2XvvDEQMWuYZwICvjnfx5Za8E1EDIiFSVjQiiaExfjPVG+sO5gn4NFQcvBdyatWQ
VcLNbHaEIx2Nz9hQ+sGyEgKoodPhHPZxMQZJzgPrCpKltyvDdl0rAOdPy/0BWDAC
l3EWtSUpgX03kcz8EeYw5afqRI4beWE6rT5uvjNbL/fTwZTt15vLQAl4tHVtqp46
GyiwtZ0yOS0PFAxZGVcqzJ5kPdNienL08wQTpL2pMRHGk5JQ5iYVQPfQ7RmWyuh8
nTJu3ejltz2JsowzIH0bvrZzvpM9N44Rxu+PM8sf3U2CRGWE4xav1VLnB+UKlcab
H2OasDl/Dz3RHt3vxDyUDIweNw4ZFWGivZIFaYFK/rYy+DPTUPN0x3x5rPo3RRF7
rXVxrow9OsKhKpXtS5q3Ghc0NDi34RF5smx8oZBPsujPeFliVAJxDs/ScJuDlDc4
HuWq953DxDvv83GOELvbiPXxtYjJgK0is78g4q9ljty/4t8U6jQ9aQKeW98pDzcO
N3pXVMLXcXcKotru0vG0RjcmutleB989Xq5MGXdTvG6lWCSVlqRuDKFDoAj3mVds
ko9Nfng1Z956jacgx50B/FvMO+Q/AnDOoT0oyVB+qijFRxCaX8lHiyWz2AczicFh
IjVCGxLSKDDfGEvPO6kSeE9VS7F4x9Sl5/vWc6e+0n3EoK0zArlLusrjMqCEV8LJ
VzgXVH3uA4VTtoA+D8Pn7UIW87JfEppZA2C9caM4/MX1INmTfnF6eh8RTfpN87Zp
AXxVD8ovYgIT/vcq14mrDDCMDXCyU/PkFpI3RWvlRoAmsLzyxgI6c+x6KmCTGJDY
v5B+93d0+ueDJ/Hr4OE76Zj0gEj4l7T4ySJa2YESM2ATRIf+K8iNENosnno93ud4
VMPrOTM3PNdy2FlMjXqW3TicccrlPxeLVkoHoQSfWpEcOsvdqEsbqL6Qwjr/assb
dXq2y8pUXwpEysOH3lIA5OV411Zb6x+TQyeqUGVGE5GX/ZnBsM3iYIqlqeIbTs1J
3hypQPRwO+yTApyTgROp5zG0asjY8RffX774dBBGBHA7yopFWPP2a6x9BDUfMMHR
/L9WRPV2WuIUwE7lbE7UrC10z6q+ceqwmMy5y38vusMJuh8bcQKLq8JjIIxitPZV
xYPTbl/U8OtEHbR9xrw11eECKRJSA135+LAEySmasXUACmDVBpwUY/3jdybHiEOT
3VwOxk3ZhGe7vBzP+7xvwBAuYANnp82Wuc9/w8rcdnTo4HjrQzDJr64QRa6njFLs
`protect END_PROTECTED
