`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NDK1J2x8Zhk/EZYVxiy3dGL3DmXglsvU8SB+TULodyz70TVJm2cnENrJ8ZeR5z4d
HLKE72HCf+iALgp1dJ8ngXPNSYE94QhmI0k7z6Kjd4k+3ZS6Ba47phNagLx4a3Ma
wUdIfhz3b/ltjBEsB4ipsWKyiBQ3bcdNfs6KvGhtXuOHjgB8q8lwhUNr0SjEvPP+
fVzk3Qpaoe8U8vIw44g6Unsp0HFCZmcYRnf8X/mu++uRJZLlWmUXZq3RCr1d5YvT
jaUvMdySgIJTyCOCj6m6uJ6kDy/lOvU9tYckeFvf0eOMt9sY6O4Fbyhujhld2X9W
njFCcNpBLUMLM/Mc1yo9KmmR1Eziihd2CrDCiD52XxSNpcLQMfTScc679qlAwPcG
7VxVDpyPBOqr/PGG+LWUPAfXnzTJoNHS3ikkYsm/iOAFWstxa9zWA6mHs+8lfcbx
gz2SxUbhVCjr2QNbsgiqBnYuVXX65NgRPXfnh0ZtxmjvrcGt8UIgEw99/MkB6OVW
cIH8dYOFoFg9JVXtHSDlqKEcLIyZGfaEaerUmHnAhjjE/1atZ62VgKJpKPUJ9fgi
7jzrc7aTi/1HXYHggubcuR3OgVsTEUAj5j8B2IQ/3Dle3/rStgVPwNm336Nj6pq2
JZr1xiyoFnI5vPH4J+xOuwq4VtBhSdMYMNzUsGWv8+U3ToU63mYtzH25zevvk2fm
84YIGLjOhjszLSG9YEJSAAik/ZUCXQos2nAFOVGV+suvXVaXVEvH4bE/vzXGuGm+
FOL6bS/L9iqE72BQnQYOYMvjgEMvVJx9hTfVTSO3pZ2vqQn+f+NjtQouGTrxyg/b
JCZBIeH7NxEN8D7tptjQ+Gc/F6sM/taFCyGqQdCwIZ8We+LwVgvDjok55gUHoWR7
kRTdFAoT8anW5stlSmLMyGZU/5QYtmOTShdSUNvy1K6uNy4XEieYITlfQOleBUu7
BNf+Xo+y5V2eHqeQURmRQWoPqKbrU14P+QeR5Ujrkvu7aWT9PvAN/VIXkzVisY2V
GaNXNMUfm2/lFlnflkuT9mmKBBLlQMkOMi88975S7vU7oQ44RRZ7Kf7avjZjrwOO
xizfCn581ImTqGLtJrUHxDo07AOHx6djn76wF2Qew3gQFYER/6qUiI/HVO7YuJOM
sSlDXF9MjjduJ57GHwq4VI+oeyC+DvS21138p+RHUAUxGl+pEqSDa5VVPMg6x2uG
nmGDdRB37UIAw3wFGPgBOmiYctiodkx2+atj3BVZPfH8CLgYQy0oHy3kKjJ46Ddt
/htSVNUDaFUYvg9rpMExlPXZIU49e/PSzw0m2lzYwT6HNeG8n5HRVdryoXfGMyHP
gPzH6FVfhyEScHCmDxcZZIROFv/IFcJCsriFUju5TqgB64JpBoReXVMUJPDx1FxT
y2cRwNqFWPKO+HSDK+nlp5mI91WJyol+M6XTfepMWmPptLrd7vmcDS2Avz35+wif
7oR2TMEhv0peJONaZbqAE53KD9ZKk4Erq7sS2dL8PPSR9mDvFIIggRGMOLDfluYQ
Gbw7ixgtzkdqyPcSmcCZ/lGlHdhwWWGZqGORGVrm7q82tsYcbl5g4dPpj8tjoH+X
Iu3UU2GDaRWqESmkTy/pv0pgsUE2MxyMB7DyhghX1nrDtBfPIw/dHbvki2abLYR2
qqajYA4CpkDwp22o452ar7RNjH2ogr/ag9rLOLPcVWekx7+dhCYokeK+7V9aDf7V
so37+Fi1mAf+marLyyOqSQRbFR6x/3vkgLFteMceZxIwXDPxwHAi600r9pWRJr6u
H02IsnDirCAY/aNnQQmM6LfG+BZsLnDNys7gPrQKlrtxnFhfF1HOU5tBDKqpgZY+
u75mDNIeUYb6IV9bddRyJeIk61xD7kx9jOd2pLyD8t98mKg9ujpxE2/xmP36H7OC
iUeT/wsWAAvG1ENCYbocPSAimcZCDHXv4cYJYoUgLF9isnFmkIx8jy8+dNKUOv/e
ymmvJ5gVqpsEjP6lUgPlCbIQxsfMpEopT1zO5nusZZCGG1xzfXyV1VchCEbntMf7
APtH+2O89pD1xhvUTreo7efEZHTVElG5XTLdHVJsGR0A+c54s9OXmCGNQCoxiFwT
aHsZJdovvHlONAqkjg5Q+bfzFG9tags7+nIQsJFpiDq5PWE3CfqQLCkzxTBEhCUR
yVhZhIqS4FYVRef0Af8rfsaSa5pN4Av+oAYe0ckvw0NfxLAchzCC/j2XB+CmGWKk
omxsNVSrZmzQ1Ycq0wWLAzzv9OiKEe6VJ0derBGcIR5tcTG/hqeXvC0Bo/CmftpV
zV5g9cy1bg1EZ11tnTbYf+Y9u8PPfaWIGqp+81kMAGN4O7QgHNPov3gKFpa5Bnag
+G6w00MKRLO1FYNRLjxh2bOVTCNaoVwsk/zWIrxPtNhT0OVqksURMApDK+bCziqi
pbHMeGzZnx+SiXLsDCKNdfD4uzdtLI9VgG97GiZgkWqODtXuBG1wKY65yu28aV7j
4tQSstXSsR7lRsd2SH8f778v0tLvPJcM9mwNdYTDnZhvTodVco0kPyqh5ZNtraeD
vITCGatQQbapebk5CbR6tIKFdEHSRyyOucbbCa6VYn2zs86Wbu3xTQ4wSwH7wiEC
7JXd7PvEYOW7fLo9U9m0qJXrXj5wBWof74tGKVm4hQsyCohcSCkBnJF07Dv4o8pY
a13+dQ/reLfK2RL6zMRbYRFvcI1iC/gxfbtTpjuj2f7GxNLu/ZwA50TkTO8Tscdd
pUiIT6sWdN575YHNBzpcWx/rMR7IYWwCGvOGpnslAWpQmIT1IgpjgheW/JiIADoe
H/8mCsOp3rCiT8LTJHPzJPW0DDFPbG7jcAF7pQsuNnFgnhPFMtj57T7/+40zCoXO
JehzLiH90CM9tqwNXltFQaRXM10JzEMka+TFV2ZlKCXEiE9qIt/a8qYCbroUJMku
R2Yv80V6zGc7+5Zfjp2rqvNSKLRjAXFhCF9H1FLsdtyjxhBHn+HzulYhgeoTGTru
`protect END_PROTECTED
