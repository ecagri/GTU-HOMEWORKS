`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5ZutG2zbuLQ07Q/16SPR69F6CeUFtsmKBL7WRF7ruNarmH9ADGYSRAfIGbKixiqc
p8S+rIot37APG6LavkHhhwCPHdhxv9ZFIPojPjbF/3jsS2sVW/7WvfiOPe4Nk6s7
L5kswUyrTxM6Y+Yni4tkTl2J5o25a2jRDfO7YBwPBxUQ+2br4ZMawjLmg2aZbS/g
xwmf3EHtJ/TMj/4FldtZyWIGZAcdrLktW2xaoL6CGh09Ta03/8ZZYDBNV1FBVLji
OkQa3MxMEyb9McEAowkBJaQpaMMRIlPsYPa7mEnRZ2dmYmK564X+aEDx+JYf8TgX
ZX9L3O7TcKBAQgHKgyvwbhausnEXHA2HglvOlCgPvB1pLy6n4jsRJmyuDpXoBgZS
UBxNZhF+6Q5taVrPGYxxpsOv9kU3MrhSIsH3jCwDTlLSYO77Bfdj1RQCFjelvbE+
q9w1JmMZyhZeh87XYGcw6IXwjLNp97a9uwwM4BtCGdSDeHjMLap3S2iYS0isC8g/
DgaC42CwJ86oDk1v5SgOco5ElEIyM995Zw2r9LWmlffuyKnyPnxRoMAviuWaodiB
QDrEiv/MxcriwXOGwpPFHGCF3XUrEi9fo0ILlBKOho4/0iDWTXTAdaT72EdIXy76
+4DtvYiAxq/kD2z3nT2H+wa3rj/A1mQvOrjWDoMlPdtOjStWt6UpPr3Sik4bOs43
b9TlKKF2B8PlbaAicAVfmPSSKcJqfKD251l2ZK++nLs=
`protect END_PROTECTED
