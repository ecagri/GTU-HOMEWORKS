`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rz1RQ1Xf0SFCsV5RFAUYMy8KnaBLE4qPVIvUCZylSzhXpfZ9ZMLs3Mx3NBtkz++/
cNNDLK+LYbAiO/7Ep4npsZnwuMcQupcd+QHOPVkrcaCLyAW6E/eBxHFWe+VChBN2
OBdI4Fx+AO1CS3E3JtEN+FzlGa2jmlEz6PtyFTyxNkozgW80kjM3HOuE9orqIFfB
gl9xRqOLvAN5lkk/c8JfOp4L3o50V0TzHSgjqXODLenqeCKs6vyMuk0i4vx4dUTh
1vfJKy8xERV1lO61SKBdj4L2sPOeUVESJZ0s9c6ujr99jOackcfDghQaEDp81aBs
Ab2mBSDZuBWhcw9B8cFLKCvKMCRbF3CUvYmpbk6kaW3hyZx13BIcT6qKQL/FoIll
yab+OHaTQ9vyryqalYYgpahy+HkgW6A8Zlmgstt1aji93turG+xBSLIfaSpVN9PB
YxwDin9Mtkr+fBQDy38PNlIeh+bPNKoMhrjALWTQREI=
`protect END_PROTECTED
