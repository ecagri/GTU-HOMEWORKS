`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kT+owvt60OuCdgYdCKlTqxbBZEfv8IT+4Z0ny2vetiaRzFNWojzm6BEVBcnwnWcM
nmA2z7xp5u2Ka/k/lSJnhIQXeQmy0WP1ihtQ2T5OFSyLNq+Zdyp1j253eMFNpvg9
PNMt2nay/ZT9DbBgzfNQlmFGBGIMZD0++8ULBWw6Qr7Ghrq15XIkEhHAGbUE098Y
4dzhmEBmki4QUHJ8VXaxAFJaocq3S4urMPdXorJhqH7R5QJh3I02uhl5kObwRiq/
znw9271S/etIJjK4u6uX0+9qSxZBAG/F45/hI4mgnd3oKVmu/yB6v9Re8RL/km+w
WFI12RKGKmjtblmMFkVwKveEHD6Yd7uUfShgUhVa1zHWJ0gBjrUQdu73r+28m2zq
CCJCaVODRJfMv5e0vNGpK5Hn8gDyW/inArYFE4vYl+cWDx9jYI1ikCVEY/6LEwVJ
pU6nY2vessjLT889TR42K9226O+tAG93M2W46xWHmh4ADwOHDDMlULHvHcxR+p4d
Egz+ciBqHHCDJqBTPP7vn552De9QhBoiMWbL7UHCkSmDOj67prZQJpiB/HBDdldj
nVWOxPJDJWYWphQWQ4JoKMx1aeuvfxGyh8OOn2DCZkEW5xDr/HT+DEg6xKwEw+Hs
hMYtA8kgMM/PKi0CR5twrSahXgLtOG4oTCzAcuVFaB/N0hEohvLHsgr6ZlFyKkZ/
CrM8GZva36AFgvmMW1pcYp/wF6yZNoZ8HqKu5d5JVSRSzoI8b0XF8rL+61hjdDQH
akRObvM6Nf9JxoYOXureGivxNbLUcjaBpzx3uOkGUUsqPnHyM4GHem3ww2EKrCQu
X65RmDMFoHzPBzpAl6jpa05b9T0OI5wNdjBRxD1hUnMmZFtQtqRgjrOdzzihqOwp
7aqEG2q9wC7U4X4eZOw3VErDpdNfTCNfSGSHYYG5O7+z+2V74VV6X4DId3jioOtH
1ZW7fVwvxWVeaSu/e0omok8v1jT9hk6hhpBlOyTCTkoX8Y5OV0TqJI0H2ta+Fsj8
sclbIqeTqRCet/xFtg1Kj1j2pbkhxsE09R8vtso2H88K5NpWf2EPVeQkJD4fwTl+
Gtf+71EHSvlmPM7GhWyk3xpyM+NpCKbL2D7t3ume3oJxUpYpxDQttGyrLRBv0amm
HkI7VZX/67ZhMEAMVBbfrwY0fZD0qKKos2my1hvio/GDzhD1KdIvLEYyoUdPg22j
eOjLAWRDc2HL946ONGo/gxQUguVXLGSI4Uhv1DDGsqVifmDwURhHiAF19ZKbZ5gr
SLA7SoLyyG6+JaVXeiFcd06fql7je7Rt9F7OyIkQrOabn55tthaj1GN2OkTzSglH
UOxLRL7fIES2IRv5ZBhtv1UaYVjl/7KY71aI2yDPzhXzVrpQJRVjX4ylkfCyStZg
f5VfzHDXdG6p8AYnHa87XMFfxST8RHpbFkAGwf20LAB97EY/GtNSsa/thjfPe+aP
GBRdx1gELAMeyMLMyTQibw==
`protect END_PROTECTED
