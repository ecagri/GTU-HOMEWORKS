`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jierkh3fhlNC2/u79GrurkB4Yt4kOOF7ruI9zszFSrx9837FpKMF+whgIRQ09jpB
ZBHaRUr9EtKWbivxNTXVi7e/K0+ISWGdxvLF4gzkpDstzb4/SJZHa+LgpVzM3N5R
jfw6sxI09uDz2t1g8k8H4sJysoj1NR2okq/ofGziB8fJAo+h3x6E37xETVCEgRmB
v59fENPelPK3ETjN55xCkrBjIN8YdSAazPPpBJ7mMtrSssYAbCU1wMiDifdDj+CF
xW/OIlTJdipU4NcV/XE45OBFm4KZr7WuDjgmiM0Mo5a1JM0bCK0WBsiw+4u8g/c+
XL6gsPbDEO3dLHmwA40kfiideUa6epqDHL40Es4cUYojXni+Q6xS6bJekZxoQI6D
CvVa0S2y1/LoAMIXQuxY5BMoVAj3xh6uIxzCgpBD0fW/zYGx48biWZHwKlxU6KH7
P6u8BKFFaC2tYN1DVFjYsnGv+AKk2fxKFVtagLqQwoAWDofVzfs5DKr9D4PmQqyE
LATxXea2Q/QiiCBhZ5mORhwQ4ab7UIcbpwhyvKQNn3jZEpPXfpGfThGqtmLTOAs6
HU6tR96stVjZR+8RHRVdCVuBcdz5++cm+YIeInM0nVyC+lJGsGWRVLgvfKDU9j1w
5wXJz8hGDJXhdDYLmKLpS+GVZkU1lV7jbyFWLg+QjRqIoef8dCLO1RiHjCWUaIlS
DhAdiwh5RwynG/FzRpchwgRufBhB7FYyqW4iBeqxnyHh9puwVFjeBKdE4wR8h66s
kPWb6iDjOsHEnPYgWOAkZjr2BjQsoBtBCDPz4sBkJb55NtDtfPyguGFltcB6H52w
JYfUHRepU6LWzssodJYzpuEvt9f//g7LM6AtaTQ46gfWgdz5SFGFgBp9jwf7TmG1
YWwPrDTMIT0/+/9XJqzl7EJlHsUD2FVK7Rg08+NtJ6aBl9CqG0irMzjl/Pwr8/Xg
KGypSRGmxtU0IYmcEYH99aKGfU9ismv3YYx4K1dL3ebQPvxUlARwpVM06yAo/TPy
tVJwI8bo2fpC6lVsVF6LW06Ydw3ZvwCZevBE8FIjkBAFO53PRRKLU9SQJXWywnPx
HPycynxvdJHiDMsxQ7Wb32g0SQJBCYX2BmlfFFx7FLbsSlMvNjNfh91FizSkRYYL
+AtbM+52J4/kpJmUZyGxuYjnVolAdXorg7weTykEyuZ6P/8KbiWiW5z6YW5TBpwA
cvK88ihihNchJz4OZgki4vyTENn2ecZi73iaovKQCtzrq2OaILN3uEB/sU+oS31p
4fn2n/d+9nWLRjm9vBvwpcCh+rWd5VnNQVv2XozOtfssxPzmjkgQeaBVOOEXxt6P
2+XCFTdW6IVlX9CFhRxU4j6+BY1jZqVHVecwQe5vzrmqMf1kZ1edkcd6LCCrbjto
AmJg8EwoySedFcDSbHNZIm5tO87jujhFoB5ZlMD7B34T27QA2nZWjc3fIL26L67v
sG3gVbyJlXXVv8ssYSWigZm3Nl2tVuIZYvW3JtBmPlhBR9cnWpZTF0Hu5IS2l+F/
JSblEy69MxRCDfbVgmh7ScMgwNIjvqxd2PKSghB6w9UzSMPtzSdOT8AhIDm8nNXV
8iS1tM8j7GtERFRuCe3ShdMORmtrxF7QF+OLN3f3bRPKWkaPJXG5cPcdzm1FCxEH
cB0DrsJeQMZDj26jJ9xBzfYLqAd5LthVPXPU6W4GNduLmoLb60cxERoeYk1sjEBi
N0o4bax8pMENPdi9n1iO+DjaGB00H0PkNMq3mCkynWduB+VcCd4HYJ307G2r2HfW
rGML+HPtWt6zU/qq60tW0OLOgHeIJ3IjLwXIL2gcK/u+YvBjEUck6HTJ9sPv0nOb
EgFsFee2sdbYIdztaa61uiDiPpg7pCo67sB/61osoG4EOSt5roeFo6sdd3+X+kSP
HZCp2MUGd3RsPukDEDEc1lPsdTfDwtn6iJm0IH9ixJ9AE3Z1LSnKLLcYNMJd4XJx
Oesk7yAhpwSR3WaNZVsymw9y9l3LDvekLRboJq5+OjWY9W3++ctI5JeyK6O1GvIX
EGmJb53MYs/PrPT0I+4N6gqcbOtqRDLvxbAVzijm+YRIhzpqqGT/EVfKlszLDkTu
rTjjOtsXnfxWEKpe8Gk0XAp6EExZlDAzzt6kkAPMdn40LHaEUTfH03mH/E0JJuwo
WT5hXq+5AfJLewDOhfMrp5GL7fD8p0R5CH+6MLXzqKn3g0UJfcNe6HQl8m1rsHZT
yaayuBMjRAKFWbNGW0JRLD8daWipQ+UH3YCivc+QDy0tNHuZpSc0/P87yc7g9CUq
EEDZTxmi0Gh2MqgMyf2xk8qjRKTAlATpOEeV/9VLjaw+glxoL1hAFi4zDGmU9kPO
835QR8vVVCStvIHCiGTumHsXrHKRwkbeFhOUCGbxbBEkjtChujTFWwi8oOLHbH6T
7Z/DY4xaGAUh9vj1qjKbMhe63ZRHpSipOV4kGW2aiZbfVXCcxm7sdiCKYJUYBBca
uqQaQgYPuiPL54uqCrBuPJUpI0Hr3IHQRpSxKz5IWWCUY8pc2nJIyD/e4SlXWz2V
OJo3Eo7fmsrDS1wJqPPPNwDMRwym7rzFSK4E4SR1kHyUJYiCFTqvZXI54PMtaajC
u3Q5XRH9hYdUtT8btQHWIqNgSMehirK5kl0Yr7k9Np5orcigpOyVFAmVbkEjNdb/
StYsSy8+ull2hikhCGjgoNbOidH38fNP9CAqVL/X7xjzGZYj01B2ESqQ2NaNepBz
YkZtgOmB6p7VqkJwtGUYJb1kwJp3/tUwcQGE4isKn1dl84jmy/Ur4BaCY1oyQd0j
fPHrA0u7QizJVKDuIcTZB12t1xLHq8of5Z9Qwm34sNiCEF6gcENGxfL6rJfJ8een
hb2SMVoJgTbmLSIQvCFl315EGjkUMBtgUvJ+ojxOHMSav9KHyK8uBHbw2ma75BKw
Li8R6lmc8cTW12M2EuEKT6LbmRglgrKbIl3IA4CRPMhl6/MUcUJV3heAEIhsRWw7
bnemyA1UkOQWvW0Ofs734IfmLkuuEekwOkcdWiU3ax4kGIswIWnx3LPVoBfGLc8Y
TEUXV8rZXxtIzzXteAjBr7XacJ1d7ZTr0/Rcm+lG5JntNZX5/+dwQZF8LIeuXNlP
UneESgbuxD9dD1A/TCOWWRuya9Q4oZnu1sfT3Dx1fKE67wWvfX6Vu7qqvvYVho2x
PqbtMWg0k4XEs+dIkx7AsOMVbbrN+stjtfMVw7DfsH7F3zSMsZer7oYTCAIcLxl2
/K4LRxPGCWLCJXJFmYTiHIJF3vkJgtQ+OZKCtOBKCf+f/VIGbbwz0H0Nu5us73m1
t3kKnAqm+Phg8ZulhyWw6bok3JFWAJ6B9yL1FUCfzPx+fauxIikx6iy1Z38WFcca
trU2gUUI6jKSeQreGgpVP2Nr/Z1LwlVL23PamCSA55v+GJ1YADfINm4+VIn0iQq6
7yjaoEpQWS8uvkg+xJyawiOkOQQURWOSKsd1HWQ/I+4jQ8fMnZ6sh/hm68sxc7ML
dWFyek2XypMiT3A6iPFTv5KXQxLwykhUOiNzT+uKt0WMqL3rWtl9u9yRxaRzB4ba
F0jURt4ixaN69zWWa2DgXgCkPxEM1UOMUzaoPEDcc52QK+Mk6BiTeDj1VgxkQ0hb
e8W7sM+q+CR4GH7hTSiT1sMXc1d+Je8zYcYW0pnmKYNhf1Ov9asW5wb3vw3tmnfO
ANAgG3JAuM9X6Rz8P6XTYuGZypX4lStfUWRI/Znox7QXQCYgRrpBNLf/Rcjd1dUZ
tjs0zH+TvdtuHBrNA2MugnFYWkzFIPXZtOfiopokNfdB2KbuZLDONbIypwJJU8vA
0S/c2zWduw/dLT22lQlJZxc5lMW06TG0fik3iE4dXtI+oo4t0gg7rP3x2PeFoVaW
PLgbyPDKt1fIbgtEdAvqjdyMID5S4MRsj/EJoFR7cd6PnLWdfVfCpS/xtPtFDkVN
kt7jSwzXRgpcqb+tDm4xpnxgH+rM0rMkP4QBet+S2UsVeoHwtIbkgZDiEThOdJx/
kA/FgsjHWdOgWFGFTsGu3k8eaMj+Cn99wC1iq+LGGM2gWo0fHL+r2xeqaVpctQgg
YKsUv6TZe5whhpMuVJVS6R8eareRh9kkrZ+Wm+haXflxby3OWrI1bNCheDeDL/mf
iLizzrCPE5gMyVUvCXXn7PAKNC2fLGc4RibKt5DPjfd1EnKDFEBFY5JgVVaUWNI1
bIHj+0hIPup9rQNLIG5aWYWrEe/nmG4nnA/wbxfGTG0XQESZw3nAoL1iF+bHQ2VT
rekzP3TfrYEFLQlE9JF5k8Z6RKPfRoI1uu8i8J2H84AwP+QEonvKjUqbXUyHYyzD
gHMpt/RZIJlcqGoV4sdiRhxu15vyKIxmDaCNYHhoCPQSllENuUjFIRT6YgKSgCyg
LNEhe0SU8uYnjd+CLolZHf7ANgUrKEgRBQwPdSzDScam3gej/IIxxkRahQpkulnP
7/aMzM7bluES461pHV0roKUle58Cj5CVd0a3H686oA97vGJ38EBXm2BDNkLxU0NR
S2v+CqHdr8+RSaufY96KrJJ+fMu77lEwdbMPOIaFwqOc0IP6Rv/r4sP2IHPGDNvT
jd9y6g5Tq2CwjhT1xcedm4+XGuURwHdYoixnepvpjp2bKnz8kJXIAWvLzqYSC/bg
GLnECNItk/kNIHF8Jdrf3B3pEUO05ixX9g0OZGLmvVhGHIydg7q2JUa+XLK2uurB
TObBHYILrhCNzXnhggaGRqlms9yo5qvkImIPo+V58XTPTXAsHIFdgiz0aiP+q3kT
MkLh1gFBEztYPm9yQmKcrhasqeLLYhZrA2//b5b3Lazz1yw2CTHdAA4VRnhG1avs
hmC8cRC/VQSXcQZ6lNctLxniQb14FVSF9NpSLFVWHjTHXJ4bU+EhEZvpG3PXTHSq
afOy3uw/BL41TuvRCDWogzyNvj1l7JO02D7Q1cgdZsA2vU7tCvdGMAjxdaGJlfJk
ZxIoMajMdgrVu4v2bYr75St8J6C0btrDuf4WW3GmnAH8GbwqXJ0Yp3WvwRh9upjP
QKzleAdWqw72WjEFjOFCSCslxz5cPPE7ernyeDMg8F52RPV/TmxeTQWGmUnY4tRu
n9lMvc1cnGaqlyu3AB4ww48QqPpWJmHo3N5efK1TWGev51ZklO18EUoL0r4M5rTn
9jY+BtZp4ysyIGjNCDuS/VqYlqRW9zeWJ45mGSH8YqDbRmfOBX1eqEV8RC1YphLR
VQ0xuHzuYRjeSr/FBAwyaF5aiWbZrk1Uar6vsee37Ms9eKb7gsCBa1aP8GRHICt2
YcFN7KAkYs9g4mY1OjVQ0+bEu2qzytNmHfo/d2Ghh9usnkg07A6s9lTyuJ0Gghl/
hYB2opucCGMIpcw7gAYOMoJIYBa4AJJ1MvOOiG0MwXY1qVKAyp0PzQgmXYGlyTpI
+plg38LawyYnunRH5Ny8xA==
`protect END_PROTECTED
