`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3baSrp9/78FHrRvpWd3YXByEcPT8Plxg7fwlheCCWBTGK6B5/nAIWdoVk07Uuvzu
ZZci5G2g+80+0unhjwTC/zTxXIp7hQe+TfjruLOehw1NAHzsx6W6jDn+pOMtiOZr
mvjnatuTxGu1vmGoymyq9ArvsRNzjqxXwMyjqXmEntILcj8AHEkEmiA8hspu6aus
Jbfbo7hDE+K+Tgg6GrpkKmBXoBfVNj3T0IVw1Jm35YIHLizH5vkwGdV5KoEwwm/a
MaZf+UG1SJx9a6d8f5nTZyF/de4WMt9cs6/etuuSgfCFZYl/aPzqVi4ttxUAaFEh
nXipZY5k6w8u/rvR9Hc5j7sDZjNmtG44Vjjnig4F4K9epLaUD8ir9mMp9U94Su/Y
Ey5rlIFDpDB3JZrC99XjbvInECNYdiZ6xTZhOtyo9WjVSeiCxikwMs5r811Tj4iN
zRKPZLUi9CvnRSytxF94zgGxY9L21WUrL4+/ytxPG/AIfc320PWGB0KylCaknT0Z
z679V7Hcbp3JtfZWGIWYNcgEJ2AHZuhLh8el0+BwnrzPweFwtNZGJS/6MZ83uIIW
mt1PRanRO69ckarYaugHNfyygOAExBQaOHaDNCe1AuO7ETJjsx1aGKgBeD9QYHG/
Tcwb+IhU8wUhKsQNiqrJGP6XCnz4f1D1NoU3Tn/bftcFNKeZWgjbsCri5Uv8ybjb
cpLXaY0cptRqsIfAVMO/OAusrSJI3w2mx23cEcN1JYPe1IEY6C0DwADa5V+fdYJJ
xmr1nU920fNsTsHTA7ytGHGBN108oijOMI8X8Ajs9tXz178Whot6O4Yy7L2NK1E4
uwRyvod5DG/yQkX+bNI1ZPlb0aGojXEkBHHtacuyNQPdtlpOFqNDgYsEqToVLxbu
bakuHRf/Qql/FZVIsF7E6z6A9ckmtntnPO/+yHB6wqzoQVoiyRin1uIab+zav8sR
Qx4oZh4MX5ybguPgVcasy/YhPrB+s8g2ERQJV0qg7A3Yz8DYHQbo4T9gTeSM7MWM
BFgoEt/2sdcbgw9jzLig2ERDXyPZyhhlQleAp8TX1IEWbeqvRpCUhIeqVHA93u1M
DKmQ2FNeJtusptsdSPtPCg==
`protect END_PROTECTED
