`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vUu2O5Fif4bqBXVepham2p8bZ70ZozVqfvbcqfNELtZd81a5xEnOZfegiR6+kW/7
5tIfARquCIS2WJHsDXPHPN0vPc+eB16mRHbrMhbkwnMjYGeRfqTTJS22b5aSAveZ
9/1bCBZAwqHN1OA7n33jvM5IEcnpbjK2NV0B768kCbTxX2SiNQlyIPeqwqa/Gxqt
x5QenW6rWjt3moqOJspy4oAm6OrjWwMsrqVeVQ3Mf5VXRlbROQBkmEhaoBqkxB4g
9BtO9qeSMsMcsevZXbEgifNtC0xewNJOPUE0hrkgzFDwBbEZ4gFcEfqiC97XmDNJ
VeKxdz/3PoAYlSo0pw3fKYtrp5JvbGX2KUw2i0bY2a0QvHhx7CF+nIdsPXlni4P0
oR84XRQDp66TSu2pucCWfkOkvArcPrICkbiBLLe0BDddORajwG+wsyuvsuN36ZAI
DsXN8OS/9OJTEOT8rftc5aR2vYsMYnzDr1NvoeqaWGR33qxSxdPGC9yx66PtecTp
QnkCGVEfuVIPnGhB88bkMsE60mFNN5p0uNYvU3U708TLEuAfhJsD6ntFtGB2RiT0
jTj+HuzOh19KGsufoaWl2frLIpG9UYqN3R00rLqMIvL/tWgft2Dmii9jSqOrp07s
NvT/zZ1+EWOqAAsw+2DJypvED7GeWZKyW9SiovI1fAeuCXXzmqsN87pGJOdbzktB
sDiIjt5p9gOhYe4MAz1mVVUq/3CpOwiZ93qC2GLsPj16JjL2EmBScX5D0siNMXqR
48hJd0P0rYBtIozBZ0m0GjEosSEfYlkZRpIr2xpR/MUnFwpSSL2bFNeq4yxO3xNI
fGDqmcztU98e/KC6gkUofmMXobOvo6KNWdYrRfs6HzUy5VVN9KRThOYhnrxUfsJk
BtTbrK6tLN5DR6lY+VBOulyBsS2jEcewVpFCv1EdEZCGY1gETLxnFjGt72d/A8sC
cqMHyQKN9FPrnODPx8PADPgCDboydhA/Cq03l2dGgIPcm2g+RsBB7BMG2AeT/N4f
Z74KIqcBcofbJJvbRsR/gxEzZaHN0AuW6Oc7Zqzg4LjlnUINsSFJdhRV186/e3bq
bBbdDU0Y25N1VhT3VUXUoVJtt+4gde1hCmh5PyFOyxzzroXCPVYSZY2b48GV1d0N
hx8Q38O2jVDwjeCdzrRdbMGi6m4WR+5QQ2T2hM6hDLiiJup/1z1qnO9lqCwQsUvN
2sZRKVa+WugXg3rr6DZn29QNh1RZESzOyfsjyALXosxO7R3kjLm6b4wVPaAL09l+
Z9KoM1C0vqgr3ykAywGf0xNuvlq2afa6bMuyoLJv2e7sFBZYu7KV7wJwZnYPZk5J
HMZ8tyf3TdtOJP+qMmekP8TbR1l11VVLhFDJhSO5rcGzIETUkOhGWmLH2iWSaMIY
Q7Os6od2ZGF6SMXbgXxLG5B5A0ORIxyYB7f89wjgVKaX8eae/MfzjKIMqeS46KyA
IMDMfTi0FMCcd1XW3W6yI59gvhOr/6smUUCd7rIUBKR72ufm5AZSncujHo7yTST8
sSMGVlJvRqbLTve2Jkj5m05QTGmRRwI5lVnobH9FKor0K5n8LUD0quEfJi78Hgqg
bbt9DPvp1jgT8lSWk/R4VAMQUm/TVaCW0i+F1sCDHCyId9ZwYuN8NShu5Nn5+md5
b+UUmLiMDgvmnyqmcglmYJIACb37z3KCU1+8OaZKGM4T1GZs+PNiODFPFuGWwq+U
DDFQOHq2pKhf+gSt2GMEWKpJk32OaQp4fRx+5L1r50wOTusnWg/9Dzz8ytMGcfYc
h4lVPvdm9OtVCGtob5H5NBWpcBjjs0qyjlHZEDiiBwpT+sBiIGOPY7ZrxzEW7kWU
kE4dxhS5prggQYviQx3ocwionsfby6gSl3hmVUpt7wA3duTnWlD46V4hlJ2lmWtv
SxIcVDTGT0MDJLoN+1GvBQ==
`protect END_PROTECTED
