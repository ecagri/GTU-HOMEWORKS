`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8ZpmfpXCOQboRfCPSlx5bmoqo90XySRxx/PY3+VyjoUd7btYcZ6GXZPot5CdIlEs
VYK/1ySSyAW69FKwnVYSzs5nxGXH4zDUgcBMGmc7LK81B4Db7B7Us9wYcEyVKZJB
ZeDK5Gui4lt6zgoGyy9bPvBNXcszuW/s3M2rhGjeJVbeiyqiAGAan4a1dwbLkFG7
AiRX0I4uLjtNYshBPI6RzXEEy02TtL+uRXUq4mCGtjOs8CnsxQhiizvJMYooSH/V
m2TigwriRtx/IWHWsTJSTOrdZec3MfITHFwc80pf5TwCMW89UCRqRdjskoRZbXFZ
voqgQ7U6VnVn9BcaCobmEsZ2yW3Abr2Lt2t/V45z5X7NOfwZtMwFR5aRpdhQrw3u
/hwHltB5HPZFQsIb3MDo2fZttxmSauVr1rxppWNQyzS9hLucIQJr1mFilei4W2QU
Hr0hdHB7HhOi5hPZOTy/E1xvHbgZn3GhA/iLQqnuB54Bqdt7axW0/5QOGE5Gd4ZY
IZ3rhA8Vc2KgBddYyM3lbHZV314fzsos1dUsV8XhvCnnqLKBKqvBfLa4jdLb7hH6
MbioEXEWmBIxArS7VEzS9FBNJMm7DF50Hacj6Se/mW/39hRnHONhVt3aclaNVjQT
vbtNIWH51888oZ2/ZvlaVQ/7/FlgaPbmmP35LEmyh4FDEeVY1vFLE7OG4kXxl1+6
7+Mod0aJSlzarWaFZmHa2ZXoE3RVCm+h5QlTxbWCVImqpRZAImwwhkIZsOO3tzuK
oY/xziCIPKYfaU19W0ppIMk+jH3nCkKYZLvanET7ln0on69iNCbxCdNk12dqYgTR
RNIC2RjlZmmUxjwJzqOklWMIfmbCwAHKt+sGeE0t1Rpd3NXfnrbsmJPZ/g4n3Ua+
kd8BXQk0CzoVDdc8cdn+1j21vYaxbT7PR3frAV5oeeVm2zEQ/rWr6Mv6OnNu6lsP
2+L59N2kkNzWQTw6pgEmyDdZSg80GW3yo480WKKWWBPXYGLQWrPne7bRWdVfZ1mO
ZokCkew8d2VhKYa7Di9p05n1pte46JIPWXWU4mQfxpV64TP9GlFj2t+8e28UzLWz
B7yvlTEVWS79KVw+lqsjSJSP8+b/2xTTIz/C1d02YIHe6pF8VCzZc6thnVN666Kp
KzuiqjR4p3H4Hl0RAci/ivpEuPAzsdUL0kcgNb7PWJBFaTIzgL3d+p81X+43CEb7
l+Yl23QqjH7RCoov2BVqwIyITIl2Wq3nR484JQafdiADsvBn2jDishl4b5E3UXGC
7VJ+mTghZnB/anxyi6Hs88EsHzZW+taBiM1388aYFSkyvRirXaIrGfiIN2YrusA6
dma4lGssrbV50gOyIvTSbMcdJEe0Uu+sRjDjhe6i2kwA+k/gy7LTubzC8OEOGs+a
jltseaqUMV2PuY4lrD3wYQ==
`protect END_PROTECTED
