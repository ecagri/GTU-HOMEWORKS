`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nvZGFMs6y7kfcnnqH/ZDX9Z5UwQKwOHK5gu3dcw4ZFS9tjsIaIO90h9LrhCKw56B
65N46VoJCiV/GthbJYJtZLbpYaQQqo9gx1WRNNKfvfhXBIuOc4Ft8xll1l9i2Zkh
NEL/zCwubcOqZl3nv6h4dd9jdPBlq2I45DoWpmWLA1jJs6llT90n2c4ZgKCJzxXl
oZTjPu0CZBvF8oDwxQ64Bf0wXQ5+YyYpiU45vQI3/gI6wyWx2en+wEy6+8QDxTK5
lG7sS4gO4HsoY74A6GXaR165V+6RRefSLOpfZOrl/JfbB2xq6p8pJFghO/ndJZPD
Z+D0+xZWosh9y3pwex5NgnEn25qSqX/W9QXlPOD0hM64NGS01TClT/84dQDASIgt
l5SPOMuqkS7w0AgGpbx2ChbVRRsDmR6bUtRpi2kVP4P2xBwtU9roZ47vfHhmdOCS
TEK4AwQhQQV61ZKhua6YNnh1kK88SNWvDfuPmqZNlxRHZdO39Z/BVVchDXptAsmw
zrqgmPM9a87dZsP6tRTAAgyhQ9wBcNZ7VeGbBI9bHnSlDIy25ZAf0WuP7Le67lag
PQAcZTh5y/6xK9HdzOLam/gtA/WA8RKFrML5/h0+44zilhAffwtJs2qpQe0qnUMZ
SMSCc6YEp26HARn3QEHEpk3QvqL2dnxHyWazbvLrN/dowe3nqaNX8uGToaWYBMNO
yGGyCphZPJs/EKDM4Oiag+ApCCWgq/FirjXIY2uI0VCFPMsobxFq05QETBfz9xQu
WoeUEFUShGumNmL8oCiACeR3lnQY48LTdg1vH8pOLu7IbqTq1SplBw5W4T8yZXiV
x+dNUnDWmjhUwoJSMON31Y6kR0sDdcG86bSNR8rc43fvYUwrXy5wj6P6Id7SgL6k
+SDyWQdUuZwgXQeR2auZzMNx3MBeTplDlfAPBB9nc2rv0SPhGAlGGjmk+sX3HjX9
b/8SUK98QO2eB5llpgutlNNXVLOBC/Se0UzTBt2UQO/JtHsIunXsyQWKbm9Zb3cO
zz+bQ0pC3bHbK50jiWCZWJ+SnELrrtZZxZncINklIqSds4X7GrIGuMPFQyW29thM
0tEDGzRNnFBDl1J3PtO7suveZkAixHCb+nUVvlgUa4w78mQ3yUdCGaJjALrBLhm+
eN+ANucfAhE/V6NGq1nSS1P5ZTuXj7p69m0QfJNghVFUS563zwQ6/8KJZ0T1Dq4K
Wjm+9j/8TeVEKekkOPSTZIDlYk6jNY/OVYvEQ3psBnTsSJR0Mtcl10NbnfWW99DG
xhlrZggFuJK3ICUJ0F+2zaFulYI2Nu7Ktu6GspkE4SfBjEzHN7/4ayYYL5WatDUL
A8+SgldGsdgdDU0RTKarHmz1Dr95ceYmOkB/plfiGS3pNw12UhGFEjuyMBl+38+K
FuDfsD4J7Srqqssx/FRG6zT0WZfk/qCOMYE4zizAk1ix97Zq2k7gN97fJgEPhOet
rKkcnqWr2kdomRXvEYOjgMGinVpKv3fg+JwKJ4dVFG+kxHczaO7qIThwBAo/1qh/
dePVNboOIhWUeC6sHYUfSBJB3aXZodxpeezEtNP/ou76jLymuwxiVdvCfHL51q9G
1lt4x/HOV4ErFOx2KSn/3VxKdB3lPExUk8puku3Vcyu/43kFqFYAnx+cMbK1zknH
SPhfm2TfhZbDMuDSSn1r/nKYyVJ1fl5XBSRbkrEYOaH3emYskzV3HwsTlWBSoG9c
fkxPIqslv54kQifRHRyAyNfO9GuavsnngbjdgBThlRvjljyrG+V5uNLRyEOVjEQq
IaD7of7EiPbZMeMsMfekrDSYBKqXLZFwHWsYTLqa3yquZ6wD9buvJsAPCpe4VM8Y
D2AppsWm5LyM91NUw/BWSceyetysNykfxtMGRDJ/AcWg/8sKObXallu0jgpSJ8Zz
IRRzOlMe97SWPp3FGovta3i6Y155+ZJvnFocZPANb4Fc+ZlnBFa60qoorSzqxS8+
IZp2clYyYIPB6P5J49MGEGf7fZjfUQOLVnWXP3OKGOWSQHC/Cr8VbedWap/dq5c3
x8Sjr8jcAzUrPcH2MjB6iPL0CoFlDR5JrKFW9c9DSKfj1tc8evyb41qBq7iWrxPx
6XfYEsmzZ29WcnjHLz0VADNUzXk/E27jVWJwIek8K4fp488po0omyiJ2TQPwpI6U
IXTkVpQtobVg6ygSFHlC2DsMxz8tD86CozIiA3swjMpkeF22ZkLcujDzCbwGF3hf
VDbazGjrKYbkqMxUcIBgLecoxl3Neapz8hXpdRUAsBZhtaunyfqr1HstQ0jRFHw0
kirN+UhqXZe/2ENEyh8pMEKGq9VpYLA9JECeTmq3yjIO0teV2yZyDhTJ54DT9MSC
JRzyU6v7Vw45+Ce0XsgoxwSuFpvi4eSoSbtUiGOsZdANptfaF6Nkv2M8OdvPbNm0
vGHF+HvFGKyKnJ3GrND8vLlOL5Ibc8Dl4j0586bx67E1NolHJFHG94xzSZQt4VSm
AmEyWp4CS7M+xpB7pMBg0MHXkl6jlTi9tLcTeLFAIE2JfZ2Ea+qQAlRmBwt6WG9R
Dd2vfQSn8kOrRzF3Yzw58y5jsoDwTKtbqCwu+rGINk3LGI+oAmGuGYhhWg2mhE1/
QfifXIjT/4xaFnN53KOXZ020gxm2JMPhXynHHOmNpqc3PPhMYav/kFcMLHV3IaIN
VEeBpasmUF+EjgZeR4UDOcdqwuMghBoMay4L5n9pIvTWCOSk8/vD9sDOk2MzLIIS
sGlH4B/wXTYZXZuvIxEnshTBp9ifmW/AnWbCHDaT45jgcvu/E65OPepX/wDQBxXO
ZRuZ3xWv6NgD0q7p2natWMF6zUb1NHFC48YsoX+bsJ7apUn6zA0lc/hp5uXlWjxg
yD7CM+PcdGk6ApMjzquOZOqFHl6pNc/Nh11sZhs3AspFdb2ZCoE4QehygMu9z03f
nezxJJgDGR3ouDmTunACFfqACJtdjucvSdLtH8w1pcfZ24WZ8JeIy7pdz9MRxhOg
4bsauTvWW1SFZnzOlU2gN5P3x1SldgjvOeH7mODBoufyvUUABxBqb8kSBzlOpTcw
LWSFqeIZ9hTcuUGs2ZgAIRwJY4zn26naJmFc+c7jw2+9WiLEH4AYvB6kjU0O9pC+
eD1jwg7FVzxjx+cQ49kGwhOy6xpOhXamGAHhv91KD93q5kUVHzlRBnqIh//9sFWF
GK+tD0+76oZOfPKGddKetXGX4cUJztw5pfJH4lv+cnC+tMosrqPh9SGff15r5O67
hWKng/2M/smqFMa9BZp6gvOPDwHIkIkvhGs0D7WM0YOzn93lB509iFROPAkfa3Te
iJ0/hcZBkEuxSJglA7cY2bJHw4UhNmcBFXyJd2Rz3aYrKqwnFealpyRomHdvBziN
xHuHjRZa/KqqUmtnwFaVlHrcX6426fkdCxVoF2FGLHoIlpXtQN/x2MX17xlmz9HG
p1bR8etd+jVzH2LHp2evSBnj/OrHFXLlWUDESj7BbeWFZFMJ7Ju9B8xuSMulRfm+
37ZKmqxoMuxVmSS7pET4rV9FWwZHCy6qKLjF0JTSxfyUZn9m0m4Gu4SwCPtPQza5
uR/fRNAs+73rCLRr4R+G1XPei3MYC7Aqxd9spyMq5drX23pbysXrbGhyVoZRX1NZ
16wEmcZ7A9wVN9/r454St8hSHbSM2ELTDw+Sagdk9CkORk6e00DVYn6jVaKzNicU
Ekj2z7WM0tvTkHKiNgopl61R6oqgtK7VQq/gT00Aq5zKxnJHOJI0qy/HJTsEBfRR
6g/ufhGaLz4e1fWy3UHhVLm0iHtQEc9K7D3kdHoENotNjzC2E+eXuURTACDyfD2C
B852xVbByyk2Q1sOGdKcK0TX9G4xHHP2H3kn2sMw6+7z6cu1AtPobF7ON/+hi5Om
PYbancuUEQC99ZC7u5w+wq2SUYysp9ttFnsKJxOz9PhMiYkVCpEec8TGg1/dOmWc
oK7YS9z3sXpuMaqo/tf39nEH+MSq73b85LCfqOfYHlC5hmIi/L5KhnCtWI0Wkfd3
+6ePGAzpuT8YQyOMCicFaab8Zh6YGvPbpmXevZ+y5IF12VeDgjFrmYnHHR+VT1jS
C5XAwJF7m+wdaMGHpAeq9dbM1MC6Kkbas44K4opu2qWLtR8V6JTYQgvhrvZefmQj
Y9eedH+Rn7WhVJHF9A+5ZuR3gpo0iG1+JxaJ291HgtCA/Z5//grqwN9DhVPLAvzh
IghXIz63R5YP5PAKLRovIu2kNDRRVTtW3rlg9167bAngfqgMkjDMN/86HyzVLhAL
L5q8jNEoCu3daYs+pwf7ccK37LChsBt0vTtPeEqjZWU8KoPG8DAxUkt/IynAcLTa
G2SlQKZC1GE0Z8C/b7LTGaNItCmLwTGW2twdsz1v8/mMIQxXmohrmaNIzvRQZhHz
I1Hs1GzLItYcnYThB2IaPhef9qw5y3q1zzCpoOhl01hsMQ5e6aZSOoVBKEkE3DsH
DL4ZJkrGLJC00rB5oiv72bPLmCOphbkGp97RPOZCEE7dWuccUvUE/cQGFgqbtB/L
lk0wa6llKgFNcw5yh73noRD6yv3xoDT93CDEj9MLrrahXRg3PH/wQDTpmUHf2ise
5rfxRvRQiEjAcTYJr9OL8mqjeiTYWOF8QU8dw62Ymc2pZ8fz1Og7DsxmXn8SY36F
+U1hmgFfL6HlFPhw3pDGri8D/rY4Y2Ap9todMgJNrT8a/kVGfGgIoyq1Jeo7qOWj
q1+oPGUV2cd0+6zf2WlsvNBnH5irV/ViHnzr74V+oKDpia1JeUUvmIXihlteLuqh
UPIx2RPpGrXFQpfWUOZIaPthrucCP71PPMvQ07+B5d21edQtt2PdZlD58b2nv7Sj
0VIYoNofeKSKxKCXiorCLvyJMm1Cyp4QC2wgVEdoAjImOgKvhiO13lynfKPsBngi
1ADozWBawqwqBqtRnuQgnLldJcuPto5TqpDSj6HHGPSMV6roYIrFw8C0cgBAWts4
63IQrROYYpUcQi2c4mZDeAN10ZMGb+hnf1rQzDm883Y+9VunGyA2xBDjyQfXNsbk
gEME8fdmHQrNo+xTYnuN0PfDOEwwCskYqRuZ78K9eY0oc5fdq7b2H5/t5wzl4rJS
1ZajmcYJJOoo2hjqB1mIAf03PhUYvpasxkgaEmVwk89Agy5LlumxlYmhCFpDPxSl
gcbXYtqv24WsB4a/iv/xrUB9fkBWAvAU4zz5IJ5/RAwFdpNaRxnIHsKDbYYAMZ0/
AA0XVRXc1mtucLyFV1y6cqt0IGkHUNrN6VErA6Zcw/NIHGxnKfoJVVcxrWgyAl9m
BSMl0q5xVOb4oIqIzIkGBCsVIfqCniZP6MRQ95JA83IeRcnWBNZ+J0ixcHdDDbhV
84mBPHKu6jlRCyAZSsIuhNFTcAlgLGfDVS4rYWnBzbu00Z22t7OzKpKyakA6KZJj
x+pLEQNWm1cPULqal48DL1Qw7lkq0tszbjFqgaObXPSkAlcls6SieeJmqCp59riS
HtE91J9SgHssq4jyXnZIJNNT6PdR8ThSyPpEdng6a2KQqATROJ7ciXxX0y8D4bKz
aOCQ24rrQ+6CO8EsRE/ciKFmx7E38jdhtbbLySzeYedJD2vhaBv+oU3VNt1gZZSy
IAhhRr57No21e1n67lvxoyb1cQKth2VUej061SLW72f1nOznl8brws5QHpZ7HEa6
k/s23CTAqG3DE2Wdp23sazfWbsH3rIP11nuAP+cmopWql3ahRTvBfPOeeIVhoGxA
zA3VJONtDZfIst/OvKAPcRT3U4mE4dNV/ohpB3wB8z51/aeMrS4g1lislwU6nWSc
mHKVfH6hSIyp25HzYBFjPY2pzZLJxsJiyXyZ2SLl8VlljnYAzD8aJoRMih5/k9Cc
YFA3O0LR9Zs0xAIGO5lzMarKYsN1BZuUrjEOSaS/KUm4pcB/bD+9Rh9PM/ty8qkQ
EVVN6eZSqT8U8zSOMWTNeOWYRbssVG114vZr+Je4PoOTdb+of8f/PjswRCKSreIm
OtIVZ3mYYbdmUdErGq25S/PIjxWC0UtKVYsWwDpEzz7puKNf2yV8+N6IAoFbacRO
e0LPoi6k3NWL1IIvV2IdpmizY/C75EqIsoZsarV/H1GHbn94gBIWBH/kMbklL5w9
asc4K0ReDZSu5c1rmX/kPay8kubAhR6iDbZE1V5VsYtV2f7KJfA289K5pARfiL9r
R0O+9inHaDkSGHpJKiuAVvx3WNkDOAm59yPNGteA38p7M/152iW/1N6UdQmwa+6O
L3TOIsszf3BmaUy7RhxCYgFm/tX720ivoUDpAfoxH9xncNK2fE6hGpLch8s9blrC
0McErtUqStGwMRNR2/RSBvdUkkb1ciMH20w/pfQcRdE2dtJLqF/LWhn5H/x4WUZA
fMFflPGUCr+SrQmbcCQ7LS8YjUxvhwPIsWpNxYoklG6Pf1b4dfT+/CbVkYLvzCSS
bM1kpkRxacR9xyvCqTWYaQlA3A7f1RfrdO5cKkR5Fau1DBt29GXoRduuFBn1Lcsb
LQ9EP3vjG+ULfUPatlimBY9zl1PppULZVluDOVA1zsNiZMYsRA+ALIe/WaP5LIlp
y/WINo3VR5KM4L3wRStNr8iBDHnyxFc/yfLvtTyrM2hkRcuas5NSIW+4kKrycs+5
19CODiBeNqrS/gpUCepPaIxXlKAvIKoRjl7+vukpko7ncsaHZ7+ePaR4IeGRdXlr
FzKC8oyx4FhyTib+eQ2Rfk7uJpoQrQjQeSmFmWDhkvizNH7ceZRrMUtZvlM0iG53
UESYO9yK94KUoAtzmItgLQ8gL7kQObr60UDSX8qctuYMu+ZSrg7wCtR6egbgnpK/
6ijgOm3+nDuTfWNsO+tEqH5Zq/Jr1U6jkBTHv/jhSS9zPpSNjqFo6IZNiNw+nLbM
SIylGpStzx7j7nF5gz8pOYDryTtU8BTb5TLlAU+WTvi/6y3P9RufsxJrth4LhWsa
AWj4FbktVzNyecShcLoquCrU5MXEUkK1VH+5FEMLBlw7CcyCdMsNA1qRQyyiaYeN
e9Pdn70142T5DG1SN5brPIl5F5Rlhk4neRlPE0KND7oNPLYJ6cKR6450WTLGenro
nwV/Xyd1uWXArYAuAxAe71ksUrU5jOzsxvENQHAoCSvItPPW2gJ/Dg5rucpDobPH
pI67Rx2j0qMAJustg4iL+SAyhgMTQpbbYYrYBRCEvY0ANK0xtQEA+yLte8dUlsIP
ZtQ4Qd1RYp6eXR73HIBoq+1CFM80uNMS7V1fb5K0+FLAbDVsDsp2/Kn5PRSOZUL+
WUgBUkS40baMDIbBkniUl1gYUz/32hRspmZSZpcGTWuWw2aI6tAiMLJ5PAajS8Go
blCPyp+UUPxs75VCtg3rJf8dzY5VQ/H8/p9IqfONaMJiwe7MPGiU/FiCdQu0MxBJ
3hKBtRIBYK2Y8nhOWJkiS+NurS3RAiXMEnVdy69IaY1XCn+NFZhc8FKmpxZ4PI5G
Wq7z01piS3zrstO905VoVUoHOUNCxvWganHXO7xf/KB9zzRNYj2J/ERVPR0tjXY8
Yz3yTlQapBW/vRAsRo3kQJRAJewQEjZ72MRejsnmzngvUA4Xj0oVc5bCMIRbSNwN
RJLYJDA45ueszXA3YbCdETkNlVCoBIQXRp33kPb05bYj7iCKBcKlazREuSNpZTx/
Di9CaFuhZQ2x+VahHwDHgabK7ffnbcyUzuCa+wzbQdbuxbj0i0BDgyXhlnRMr0rN
rjGS3bgPqO3nzPqvLe95ySzgK1JFUB86a527gg7T9Kyu8LvVa+eYP94meVof7ic7
/IBS8WyIw6vIVfyMNioz0AzAH4Qk4BDrUaWH1RzmTjUI2jDr8OK9zJZnJ091rPFK
BiBzEaqETAfS0kcGvXpuo/09u43ANGuWOS672rsGJJon5A5cfqJMR+mbg0h4/bq1
D1NsSzkex7Gan2KPauKbv8f3L3F9sZcty4KjR9BInC7fQw6LlQ2cA+63JAL7+YSE
R2vsNSzByGSJg7HSwUi2zss+7MCGGEloKobDNirdh2Q/vJ8jA51hCsSBPoX2CvT2
cjbHLMhFI2kh+x+hlvKLx8B8vNnlr5mNwYttNFfMf7wDy86cz9pKJr5mFcHrZpBe
qNNgYHbAr3hqt9yL8vRLq5ppOHv37PdS7YuZvlq1qWqojtiDU01MrkxnHNhD50zN
d86RIeR+d6h8nNJvxjHCPVu3FYbb4gXMVh5VnQiF3KRqMlIdTXABr02BNjE7wlEG
CHd5GgLvqS4AoHsN5sqbZbDZm7vOKng/oFgFRoNjpT9yXoQUIru6nGkXuPBW73OO
exIWF2t3nscJHmWvqu9jQpJp92ASNi8AKAXi9bCoZobhfbAtpizmw/p5wtUuP5FX
UiRy7P4SFJqKOPh9QiqpuK7W6dUgPUmclIgJfFmTlVi3QuX84Uo89jqm3O07wo48
+cDWkMY8a0HkwAxg39UzMfdrA5aelwEl6z4J/dj6MQuh41hHREwBvQvQ75L3xynT
Gf42x2HMpCehp1OZqQ3LpPqC3Y3NsTDxZX9N3zZJHBkz2hZfVU97Y4LZP/gdXBwP
6Zw33WtBddW7tPI8tLDOw2HdykYBXodFaMGJgbs0nhQQPQIfli/u6B8s9bXTTQ9N
FUf002geXTw2bya6jpqHWVd1cBzbxjrsGYIpOvP94JDbfTdzdT6muYaBRzkxxLgN
xOefEyr6nTLr+O9apINRte52UfYrrVO1QvoTvrfJIN98B1TEYdyjYgrsoQzrb4gR
3J0w1wl3Avt4lYSenUU30iW/yLGJRvZ7bAtf5u5AgLPZ+nt/QxV2MIFCpWqxxAI5
4ojRYPRW37N9pYtsX5GUhDfaNp3R4qhi6B5/eKgHlB2nWr+wkqoz1eMtobvlYlUy
sV5FC08jkTZ2dULcIcJ+s/pxoYsxSt+uW9QA7fAM5IfRxvR5vGWsBrXpkSwo4uWf
j2Ybp5thwFi8VYVRF9Xd36M4hhL+01PI9F+PERxp84Kl6iPAHDDR6xlFWlw0VCPJ
wFJFb0US4t1nvtibJnWs8MYyzsj/t0U5llsYVVBlRtz82sSPYfmwy0U7Szqpe7Pv
s3oTKqMdEOATlTlCpXUEJ2J5w2rpL1Kk52ROyZLGtiEq7l77TjyZAc5l1LeaVDD3
SP1RMGYGnPcvN953gpUWij5M2NEyOxdaMC3boPBnyolMpYqdELxoQbjb+cChZLLB
woXQgAis/jwHUAq0Nj51tm6XAjganbWUZRwGCa9z9nr3A2MpaZmjOh4iOrOtnXBP
6vJ3zeQSSBTPNYgKe8pU5ak78WxoHRQxxMzsDnTRbJBr3VfHrqTqhh3jztdz007A
y0nuvvJqjP2oLGniMnfI6HCtniZCXjqJggCth2YEtgJGMhVQs9k+kKTR+MUx2+MV
nYXPihhuL0o40qWp7lP5M7NS1SOhFpOejPoDUjSYNB3hFJuynj4za+69AjhbvtGk
tsBjlJOmXUv7uDJZ2uGdox+liAEdfzpMbJDcZ5L5I0O+WaqPOjAxaEeNUKKcZoiO
ijLKMhGZ23gJ4phcbpIj5NyAieZ6VjqWZOmEgo/nys1kgYwFDiHYmrT3Z7HXwtAT
dsR4+4rsMi3I78HC6nR9NffxDxTlCGntTu1mi84o/0WKCWFoywQWTRYNlfndqHxf
ZTixc7y5etl6tpGvYeqOv8ui1U1TskE2ooLmM8bWoImH9o/QRIZEjdETV7pp26nX
xLr1ZuOs9TjeDjHXijSGHYUVjFcuNdLUrVZf6Gs32rjf8Yz+nLqc0DSq8oP1Br5U
98DDW5VncZlafN6prt0qiuwJYPx3gUWekY+d5itrcguzv16IvVdq7pYrFE0naxKf
XzTNcUkhYhR0I/lYMuh8MO5SyYv0STsIHvO0LxMOAvb6zHtXay5zVgmHnPO2ljlw
gnhGEIG8vfRpK645IX2cOUErdryJFRUHdBHV9OFX/IZjU07Fm2lXS8glXCDWRc9V
9YzvhfJ7T4HkPWdOHPthRgB1XjlMZz9o45EelS/n0wnPfOf2yw2lZqGqzLGQZTdx
WBfwo3iWWsyAbuBXdCFTwts+phkhLrkTK5P5wzvZdndcezbSL1eOwZ0ijP+ERr+H
sPQgmnwuICp20SqFz5WQl0LkeDM4rAJ4vyL+WRBgbed2vkRToeKsVln52YqWM/RT
qMe2vwKx8FocQHx9nh34FTcuRbfbzY+vJ71b5Jt87KJcnrdaGWeOKoS3XsGdTEFW
5QoAH8vSZ0hfw3sBZOJwSjGDLaE5APs6XLNKQ6TIQztSWU26FZDCJZo+anjDCeJA
WPqRzvkGj27P2v4D4ezSgZ6s95CbaMGQ1czk/GksAe0w/baALypS+Rz2gEzTMEgH
EoajlPXXR8kvJO/CpnCirQBe+1OVAHZmtju0WVUQV8208MIE/q1LWmeP861MKkaJ
sjLgb1u8tzcJD3lUQKm+1GWkgC++Ofhv0z0XRatvFXvshtS+Xcu71EcYHHHhKVae
xB/T01s9ihzsRW1XPqZcBvDSXqeGwmza+Orjo0qgVYJSFuKaNpOw1sjiGaDc9Wv0
e9TM6d0TmXEhTNXJ6RqjZTymuyXx5wNFUsDPtv57vdgQl8h6zU3WDQE0TxXV0V7l
B5nOIzLDw0TYIQXwoOqFTEffpdiNFLdeOCsOSCxq3UqBN6Sdi5IcDYOIB5C0vwC+
LBrtcmQ/GkeHED7s+5cu7i8lH4qlD2sSCSOIk0bHzP8yJ2h+BODwX66/zSz/kVfS
elVB2W6jGpWRTLqH6BKac6SCPYPHSC/vO0M8DdX0OfBwqRWvJLNm1rqk6XEzpVQ0
wpfWrnevR1H/WFXHMt3BPIeMo4TxyNvNJ1KUoM4GqWrNm9xg670ZWIuHJmvTEMQO
hKM72HmnguzWvSOr/kVjEAnjNNEh8TkSCg6/THha8UNZguDJ9mC3uNT9E2a0S4LU
8Jq/pHcOpHIURFKXN2Oejrc2zOQOVl2kWv73Ri6/+kZNM6kxQ9OYbXo2/2xi6YY1
IGRwnt8ea+dPS3gNImB0hibjrZbb2IW/isBQ1myZ3NfdeuebK5YVPDvdagNYaCpy
JtS18pZSC+boDur3sj4guIZZMgBlMfQ5QSelsLXRVeZGgmBUq9l68/1T2ZML8eTD
RgPoYnNgq8dqOf4UDw2uknZhe3fazP3wrRxLCzrFudc9srdJ8dhUhKCpRn0MounB
rCNao74yyRaS/rMVlKLqJZNCTA9j36XynDKW7xSsO+XXVS/dfAU79oQqNwUu2vdt
kk3owv4Ib7PxgVRdfaLtQGjAyvjjfdVY+LXmTAXP7Y8C6igmMuGc2vgt20jzw9SK
M5LadvdnLpfG/WS61ac7t0nTTIDX4dcsQJEaLJoWvuKeLuzaxf/bNYjEf2KCGiAv
i1MwP6OkfL4jaEzaYLNQFQr+IJHkuAjAACSQCm3edMxjFW7R3I4cs8NaxZcKY/am
lCkXHGBnDXURsXAGdAhSfDWXzkfDgAD8PZbzrNR6dupsyP6kzhsQ0RwFbKycfRuE
43UgtaClPr32wHGqsqNNnXZBcG4hRsO9BkohTEJPtkLSo/w66YB8Z8GNB1a2GIzp
LBRcSVMx3awd70Z5LTc6E3oOp1/aF7xWs4kVVcF3T9hfjUSleffldsYmUTb/tWQL
lIxzXyHBXrbwY5OcWampkzaruzlEjBbtT6I72PRr5taNhSVKKG52TFSUKShMpFYU
4joGBixT4x4CgivGj2FtR2GiTcZbuc9fshOruXOgYcPuMPpMktmil6XfcB2VzpgN
Cjzjkw2Dg3jQ/Agd7eVIEGiSc3TKBQmePn9s6JWkBvUicNs2JnA1bIEYqh5L8sBJ
Pb9gSTUBZjtMXNLoIZKXvy7BzZglnDefTOOyMMCJEDbxzvq0j3qbJCnuFpsco0uK
RUW0rUCAVvsD4I4mpPfmNIh8mRjnStH7G69r1oYw/WxEZ4OzFVKGefIhkrTCeaLI
g2F1EaH7T0drf5CmALyllifcqI9EXxjEJ49eO5eFiROKnRz+dK6ev9QeEqToCH2s
GJ9JoOK/w4XThphZM2FTPlSBeD0xuTd3Dw2VD0/T52CUZJ3AjKD7WAdW6CvO0n2X
QxmB5+IMcfEFT0TwD6ij+q8MFXT5DNVUYToLs8KcuVT98qQZ0GVOt3PcQFMt9jVI
GV/50IyWFP+NeV2rJAtMSgLsysA6cuCmSo7Lr3ycVbwEd9Mn+zZIcUjsBtDWd9al
Tel73pofJbRTZ5d+g47f/dkpG6+hP36V+qc1WPT9RPZVVn0AFEJ44D5FyhecvJQt
TMPJYoniOsP7Y2xTb4iVV9a+OrPXTuG1oUe7D6eoM+UkRbfk0YTWgn8a7BEMvBug
nSNBvzXDXnMRrasoKG+lH/kDwJ7DwP9qxMKZtBMhIZWqZU317g53d/B5KhVLnSbU
ZWKJL1USXStAfVa4UlPqfDEayWzwui6DiM/dRVwooDJZ2NWl6ZYIF32PefJss1h2
Z7opvgkSKJoefwrGMZrBznXBHEDl/qfozrmEv0ucu3yHytN3bMwO995UutqnHRTc
NuodxzMpppDD1HpD2VXQ58T6sPK4SihZaltsZvSMd9IEgDQ4/20ZaeM3jLIeoFVe
yaMUMTELgnTB45p8+lAZAs5GtzMu1YWjx8OUalXNCfUcrYVSLf/dKruUKy45kq3F
PI8Ad429N+6cxrAnb/9CCMvBtSzWzNEYX2OJtj/7jsqJ+Ax2YUC2PLPJK3KSM3y9
FjSQzbdKVLBySjV75YnZDUOjT4A7gk4oeviO7S+aiq5kz+KjUDG4HPvaIsxguSiX
hDKtD82cfKaM7XSE20dfG4UbVMvIWw9546NIhthD+suZuT3H//P/d0CQIRUsX+vK
QXjYtxNqxRfYj49+U2i0o2GeIRhvsbWmGoZgSrMWLogjSNipawO48YibMsyiLZr+
Yop3dzlJ3sc9RUg7BixSBI5fFq7VNL7RZ+9GasVunxUnBcGLLJJJeUykfwPzIYUK
i1PSC6SI3W2thoFCIn0jBBjADYwQNTijGVUZVywLTZKLJXCpN8wG/XU4pjSuEe8F
/dE3yBkn4WN0xWD3RGBe+jWOYFkK48egfReAk3wh1mfHzFnIGa/+ESWmBT8jOd9M
/dTYOdTIiv7aKb+aQNLebRe5hnsZTWKj7ijnfqJb98SPAEuUZps/9vKcMwSMOcIA
EyG2tfviQmSLfg8Lnq+nipRnxWfmntnKCdurF538DrkkzNCVUTGgNhXT0aKKPg92
snRKbPS5F344Iuxk3mD7zy8q0N4U9c+EoxGY+GE8xSzC+VEWKBJdhCLsIW2hIof6
FsB4DjzKyD+SFHN8bmVLsRaN4kdpUjG2Xc7N6c28X8QF6VeznqHPk/SuIZKZoG0M
HWNn///x4fIPZHEqolKx2suxHfR6yQshK4HO5mS0ed6R2JAYmgxWIeEvDsFmmXUn
MJYq+2Z3fDg88kEJ1DT5AO4xtBwWrDnLQyk6hYnrwNnzZUP5SNyoElsgAcwf8oMl
kING4Eg7hiXgOTSPXWqk3/4nAzHHgITPGeaa6fT78W0afGEbnCOrUr4xM9yojK8j
JUqAyIij+eXolhUdvNClMFhzO6RNWpSVpy+AaFgxeDBzg2hIP1qQ+AYTYWE1V+SV
dqsrkSJilrcGNwlLxCczjG74LyhRO/OCVasNYZx18OJaELIDpyjl5wfCu6OAtIaU
adW5JFA6gmeW9OXaacg2BcYshUPaEtlIjr8yztxYmmRvxj1h2N2daC8vX6vxJPqX
103Mov1a74bKpvZAdbzGGPfvqYRQm/OdXIe/0BjQeVHcxhJuLRE56HyY4m43ccQ/
egB5Hb61+hPRhtlVQfVV1hld4zvuR279/Gx8x9cTtpXa40hWIyiB2QlWzOgB3Jx7
g65/91os94CvKjKYTVn4aE79bvj2d4zFmWKlM5BP/oMf2jS51ifmyBjFrpSnBaXd
m+3bzi1Vq6IQfsahyiYE6Fajzyc5bbbmr22tY1vzq8oN/n3INtvrpSBPE/8S+9Jy
1ruMGwM28dsoxcYbzsHDys5i7Vv4a5iXd/qUTjdQLTAQFZoSXka7DIeeuzsVCsIT
e1Ww/nfkUD4mejkbINB6aLDMfVfRkntLn+YNmwi/F0oj1acg46dN0kW2JaiI4dFv
iWpbC/jxzPRIiREimwgOWj3n2OYUmdyqvOVu5e1WUiKEYumpnFUM6XnCN2rYBIUy
oY/kRJm6U9sTRo45uKoRJwaNTvcy0/9hgSJD1OPoenmjlUxh7gqC2gEWRzWNboyG
cIymT3RM0WWQFJOp53BEKMGEWs+FaijCI0oDZurE69x518QFEZN0pJPxCpHmgkZU
iDoRqC5QUg/ow/kFnbReLyABFUL2B5bi+x5+COaz1/gMoEwDT5xbKdJN1HhVO0Uy
zK7TY3RbiMJUOh8OHJZA1HDaXGVCGOqctyeoC/DSOTv2SqLMkeo8WjnYjLCvCn2/
Jzqssuac3ktG4KYjvTFICrHY7dQ/SSSrMpxCEsrOqdw9YyKejsHCtLTgJIXsmNiP
e3DkpKjAAtjyG0+gTjVizRYBgHUH5NPyOwssmoSspBxfPgPlEfdN5vSfpjZ6NzHL
5jrPeRaOACez6VDPWhC9BYcUrILpBhLgPpLr87Ghvoayrqpz9K0IX8lCuSoCyVlS
ee0nCx88gIZe/AMF3fA8XTYPw9iPGCTG7Q2lxs8sXfLnLTlVVlxv/TfgPjPNgBr/
+odvzrKJMZ4+/B3WE0A+FODUtMgY5JU08lBz/It0AaJcXStQBIeEYefU7e1cKhOa
VqZB45SDSuHh3107jSAibjzA1fZo2pq0yCUI6Qi9tcV/2+hgCA7KKcJtaUt9wOF/
O+BA7XNvdm1N9LH/U9UdEf1Z7OF+CH5EtfHlQT4yeRwm9TLfX9whxfKkoaWo5U/x
WHGQ+At96FCixirzmqM4KuDFjHK4FWvwVMrN9OFHjswYgyOCZfMM40dsQQcsaeNh
5Beaikzka+SSwUodYpMms3mTbqPGGwfTdTZ7V1++Nvs1LNVzBJE7+TVz5ocgkFzP
GcAbg5NLPsohJU8DLURQ73WpJ3y6zjqpI0uGvTmr9TU0dqjuLTIZmCQr7BxUGBTx
wwQP7a4w9A5YzjHvca+kdK68BTUaa31QeiIf2NsuvHTSiL+KE+nrzK7WvJhuO9F8
09+UWHI1Lyod02T1K460uIbpATUZd12k3V0kaZnPxUFrhvTZB3GBSf4+z41DjHZ7
KhhfVzrEkGND8Q2cwEBox/uBSmqJblTr6FMRrsfZ6vb3b8HTQRdwjzOAYmiLj3If
ZEwCJIgbeezKWtqT1a9F6p+Hoeh4Cn3oSn6BVe2kh7tu6K8ujVlJhpozYuttXmpJ
VsVKIPAx5+McCCCFYIJPmbD9K2eX2wqoWsOyzHYaMd95+T66w73XkFesyhxeyipR
P/9mpnlfdsYySYnI+sH/XWEAoc7VfLjQclHlykETNDeWfTgG3OaHS/BepgF7z7xb
kZ8C0ECthVfyFIWa6Ee/MVNAgsSIGfOanbaA9/GiMhtKfvqGP23AMDLHNauUnggd
gYwE4eVQ4eOj7ijLUd+GIwDn7KMOjUryZOb9mTjMI/7V/IxCKkATNGON2Nus0JZJ
9fMiJqBAz59E3L/XEbRVu/WtlfPlyT+6GFRUgSQHNAwW2A338UnIAO0r3o4nQS71
6jhfLxY8H0Yatqcn018oLTt1j2AOsbDsixQBIRERazsUfzAGC5i3yVLkCecZ1nRK
q0plokLIJN3CH0FT66xmcETRkmd4FUqLFxwerU5nlsr1z7Z6pSXL6qjxyh9mmCfv
z3nOD2ZK5YqhQVwKybkMr365n4AhkCrmu+bnHtE/I5GzWojMPybnRB+46SEgYmzM
QtpCm+TmhsXMLeTl6mp73FYnEwZy7AfBVi8COmJ/AkHvUzIrKsXtSVqEl0Ms8NtZ
ZOal3QrdIHGF58xON9ehYEc9lxcrVQTlvE9OKsX+hdWaa8T5orUvyWRsGgNFkhap
L2QYBiFGWqI7+ScRR460xtAib6apnN3WXr090M0e7Uzm9DhPnkfdeFUf/2shr7+d
sng6TH1CPD0E25bKOfaR1rDxx7Aqz5JvLB544TblYFegLydyd5rRnjw74u5PJp/1
ZM60kAwzmgSz61Vi3Zj2uzVcDE8UurZ22qqp9e/lxU+JJsg62DTuuO4o3VmGuAp4
g2Nexfl7UItOJ6nnCFZOS8SqxTNZfwpGmPl3EiOztejK4qyJE0tToWnyv/b2QjwO
TVgNZ7+yZ25BXn3z9ickUxZhtVqGq70w9rDg68BCxtzKQ3iUGIXOMh4scFPZAvaP
NpU2k2AJkPnDwWfjey3CVIzhquWU9POtMWHt6vMmqIgYjr9ERnBbbZlpCia3igIh
Avyjq1zrrKYK0olxljV5mJ7a/am2k0ScbjufxcyBgaINYXy+KYG9rtYgQpwrhDfG
A1QnCKV9lBkSWu+BlGcCnXNpk/GC4DTwWY8EGvGFttYynGtsgwdABLD7rAurVcNd
IZJb1YoZxr+rPhOBoUUBh5xv+ZoewNJ+sFcLRE0mS20CE807QBCERv/cIgLbwfgH
LCZ+gwPYyc0vpfdfhdgt5TpeMMAudJoYsvebhPwRgzmkongfAdnEZbFrnC98/YQ9
gGzzlcwzlIZM1EzxazyZZKHo36qQDzQzjd4aHX7wLx4N7rIpk7w1zNEOqQCBH4Uf
KmmAxJ2UWNrmL+u2f6gfO7ZTeTmKS1jHWWvGdkSMyfMENW4a5QcEkDMQiE4iXJ7c
pWx1XftYyYG8R+X1V9TFoy/NNDvsSOuP/aGxVWAXr3A81JZ1FO7T6pi9XM4ubzKG
CsPbaQlVzkQ+iju9JtR5y9xFx5WbTlivA4JQPinYRF5ueEy5JgKbsgPCxFSDsmP0
RE9aUdSNHeyw4KFzgHx3B1zhbvqAQ0D8I/PuZxqnFPU/2/+HLwGKDTvsp8ANh0T6
bPyhBZ+rdsRcrUA4ase6fojQJz5WpnTCF3zmLlUrlC4SXYVYKCtLWGXhLMHuV7e4
4LeibVElgKRA3QbPkyoS5UbOfN5qugbNP7JPeDrqZrBV0MYVfMPDBG4p1YJM+CsX
WdoGNw9xBb5mnbVgMV/hz17ykDdgFJyftPuPBOWr1GY4Ofnntj0zBaqc5L8KrucE
cDHL77EHjRJiOPMxR2kBOvFPgX/FSybnMUpRSUCfhX29+Vh2SyF8G9kptxLmkzUY
yBX+/zFB20Zv/+P7T6+7Mrjgoas97WMD+EyBxI/hvQnH0pY8mxfqypzjn0B5yPr3
bLyH/3GPLSlaisuvagiQjAmyCK+sjLCVtL3BeFebdmW90qIaTqWyhE+m6eMC170H
KGTXLbqVaIw++YhUlhCTonNFwSia6oichxudjHudx4Gvja6+fNmJACDNnwYDFKSF
FcFRZfRZa6jyDH/mpDOuFT4acXBt1Y89jygimM4a0L6nyZnWTX3h5FJ7r5BDhQTE
j1HNj1w4DVROdEgZI/yyhFe8aKDwuN3Ud0WT/d4l+3fA3xPinwvrijI64caV/iJd
S/u3oqoIPLCGe4EaBKzTsBCGbgLq0pqp8Nbmf05Chhu8XYWHBVbL8XZ8qmjSTKMt
10zGrt30DseKVlUlgNLCMSNQv8YJHyiwWV4k857WbIFTOO/qETcXebGJeXpnwwgp
qmItiVhxrQvJsaQbe+8zQ7N4QfiI9ws+ff9c1XnrniH2ur4HxEn6WOG0Jlq32Kr5
ly6QwMLrqiy7Cc6J9SkJhVTTX225FFEDi+saAmKvlQ+cXONyZtcBKosBEM2Pi52N
5vJ5se0aw5ZETLfL6IPsX2jYdmLtwn3ntBOBykRxacNpQ2wEBraHutO73pN81Bpx
9pMJLszFM6IVG+/JBXCSyZC6t9fdYOuaG2m4OwKO2grr+09vlCa+LM/r5oZe+fd3
exJnynXTaNZTRVBNmM1AvKcjqPXDL0jnoyh3gVVfh5IRlAycPhxTiL9rkm1gjO0B
wT33tQdCHcBXj5hAB2a/TgRlhaCnxl0+HNY+QNgqv6qs12oSqVOmF7eiq0MdWuLs
oEZjJeOfai9Sb5/PkFolEX7g9jKRgqBHGO6O47/L4oJ7UJrgadYo0DeyYPMQr21g
1qRS1ubtt3fVSJgVKHYt6mhWeN9FDToHe80OlDBUxnTJxO57jNKTyekevTC6fnLj
wl2JBgNHwpTJg8IWLEBaK8M+lvD6M//9vJ5Mw+DMbWeepIM4Dq6YqOqkznRaUWHQ
f7c3KJVa15OJV4gNI1aWXeJomEue/p7ADQtHpqA0MPq1mGJx3HhQwF0b/7xly0C2
bnXjFGKCo9MZWcGUHgWnEhrb4C/ciPPSk7c8WG0ZHuTGEbkpH872auZR2zkomvHu
I3PWRP8i8mh9kC+lMigYxGKq3F8wgkOi2RCzDID1tyWvVQte5zXzTQwN900K+DMC
NrtzoDquMySBr7OncatOVIGncL03Hj78VgKT60W7bMnBKMXx0/n64eI6UTH/2NfM
+7HRctHZNGaIvj2tTujXCrolB0e77zCHXDw9rZFZa8CMyzE7XK8wvpkqst04WJgc
Zg/zRyrq5Ef98sP675tfQxgKLsd3lueOnm3FJ2I20pkW0K+RuKn9QJplCGYAyIQ/
rksZW4DFKznfxriz73gcZSHCB+flAZDKJCeDTBctvSM+oz4c8tH0ftlv+mAhX/06
lBz9cXeAsGruKLAOELXXeLbNv6wmIKkQFZtIcEUyprJyOcB+ugwTAXNEKg/MlUK+
UL4b+77j/dpPrrIm/XVup75x6YsFIv+VY5CSHgXeSSD6JRJj3ntRTogJknJQkPVc
nS7whaakj/XxKZaYAKwVvrQ+qFMx0UTLtFg6z1Y9H4dw7Erm+SEQs+1dnh32qp6o
2qwxBUycHxoCCIz3SpXSFi5+rGXb8ERgQuUMDflkA0HVw/so4ASFRV3DH2P+F0jK
x0SramW779gpn9U70DEuTK95ZzcPE+kcMCfhYlmJOLc4z3VExYZjlhnZ/jfnCbhi
mcQX4QDAW9FQVXepEVVua1b5vMJ7ndUkKkofGhmrhfV+BqZMw4/XKM+/zhX2BdbH
4Hz/d80vvLMDnjYc1kUeMW163wleM9wdNLZfz7gTUYWHwqAeGC/R7kqOY/Kn3qeb
PkC7wRZ4GOAFbVnrG2QVeAqmclJa5XcoesFc280eVKqhUwhDlmC+Up80LN0p9Ued
4XTksHiOjIfA8Z7I8mC4Q//AmnIbJpMPtWo0h0lQ0xsWp4SWeUlDxRM8omsjy389
NJ5lSaHJDCKTEwo+5FidVAYTBLOJ9qVIISWoNa4PggpakPe8XwhrzoM+ruziwRhU
UErKGJyPElMLu+J9rXI0/2TTg+Or9uDGpP9FkHr82XNPFD/zEiFsk3MiK6KG8453
u6WnTvDNnP6NnSrjEp1BAs4xUazscZOZEeUahGMd/oRRGdG1DzAUdIzjl9/EHqPo
Y3LK3Ctx3/SwvxmVwYMVugBxHYs/4IDHUQ0z7g4ECv1N0r8wAHjvXSxKy0tA9Gzl
f3XV1f5dNumBUvYyW4oZRJu0DMiZbdPO+QqqYm20i6dYlY0vi+MLurir8o6B1lQ4
U2TqBFg5QwV55/W/9aVWHct0WtEQz4r0cEHXUxOx6a58z6Jh4L52DM7fnXXUnOsp
uyxh1wpWQmrniUC5IT4ptqolR+X/skcHDbWuSD9nkXoB7m7B2BxBRe//1//tGYj/
5yfQeAT10pU9ewJ2n0LMis1LkK6QWLiJZGNgUGaEmwUQT9um9nSpkACGBPECF5RV
lkfDVwaN4OEf/977Kor17fRTwqs33z0Z1+utw+hEZoheblpvqU6vyAoCYlKViys8
pPowsFjpDM03cEQwlTsenpSojka5Ld9wbVr7VC1879Ine9dDeUpQADnpf/tYvROt
WmAYnJlG3gxsuiIkaYdzjJlXTM5lLupMXst9FfpS6LjHQPxhaFSRwhbQCzCiw1/s
ZXhiiNl+5uBPCJsHw+S89YxJNfLJ/f8Aj+MRwvKeSY7Q79I93oU25fY2RTYTm+Kx
UgsLbDhvqYikBB/83B5b40refzWz7qGW/U6xZuXfkeVE3pYR2irQK1bhGozLl5tP
9h2o2iFfxg5Ojsne2pl1NgxOvfT+HNXQP6gEz5kSuzPpdSOvdu3sEffBGlWGqxjX
PiEeDnWckzgub/EmeiPYQUWTZzuBboLCAXm/VkmjJuv9PEznZ1oN4MQOa4ZTc2Af
vapWrgNHYPQU5VdY86dozKSWXpZW0IC4X9RTRAzS8dl6NR/fCyiAm970450h3V1G
y0Bk+Hsoia7/zqi33mrDL5K/fOPBJbtN3odRcOEamPllGqFs14uytGySRz+d6fFH
IEJSXnUiownjeO/8tTcRKjqQofHjIuZuIU6wHcQAkAUdIYUGOpTPG5lG8+VuwQdh
Pvd7vL+C/bmmn7Hx45ZT7ebw81jtjmVxNqti+FTu1Yri47NrnqzjHhIdV5h/Zasl
6Up5zUDIll1HvcoDj4BkBBtIQJNAjDFlImB81XPF4Fol8Xn5LBrkb7fYz+7zeGe/
kYY9oUwF6B0b6mQtWl4014GiG+bvvBLfxGkMc67IvBse46cdCcTHcadFbm52K6kz
47reRiRsAt+lfgozAFL6pHz0l7HYoOwYYKK7Y9Ue/i1pXhpH9eLy+8GeR+wEwfTF
S/YWzOcFmlGg+YwHlV6dsabW7cW+rVWi4+Jo3Ia9fQW31RSsPAIpH6ocAAbqSJJA
T65R7k0Sy/M7iy9qSBBPypaZQfS4z5pNXlEnDpHXLb8RTUCLUeedNQnJIhXIazwf
3jhzdJk+mzhkV/61vJhVpfmgFvEwwyfBwQf/LTVmS+RWMVQmM1ItmYQ6+JbrKFa4
jI9uct42iFTCCRGY3YmxVKy3PLbRxF1IEnNb3L74Aof43Q7+N+ewzL+OoOFyJfss
SusHy9pVGquqL/qbFJia2Ck2/thTAuknE2F1zjh2ojaidTx5V8fDuzIEz+QtiJWY
WyG8whpewopGKvu0GVWs1ucJ7jq0Mmvt15GTxnbcPFaCv3JxHEO3q3Ao3hHPulhw
gMxSz67jQKl1XySnPFGTxuI+FZVJx/JU3lDiBqHU3+2rd9c/khRMLj9HJUf+3DLy
Xw2Zd0qdcXo2i4qNV1HX5y9RcfXxGBCWVub0BjloW5Ylrp8y+8lzmk/mIGVud0RT
3vps1QYnjfWFJQYVw476TMHzP9XnDSkGySiV71uEzmZ4/wGlFF9yaGE7r/ZbwGV8
+2+KiwB7gt/dJ5GDkJ5Y15/qy5AKAZNvXLE332CmwYdoSb418pvvo1C4VOQZJDRT
hT/+SgpDwVZmIaI5+AuSsJCouaeOWys1cMYJSZpNQaFdSWkQLuW0UiKjP2E/oCdo
A0rT0NGmBQ9J6s5MvyNZb85Qwno6CvkZGUTAJxPk/KxLniUXEFDitSKH80iTapNr
k76CJ6/2/NUtEzA7faxasPYZRkvSCXjIu/HFQ6j899Nlpn6nNqJrNIFtmyfmPaEv
VzrdVYXdR3kK5VFMwRyJ3alH/GADo59CWQ8XHccw/+kh0CgBkkJvF/Z5BMqsM+1Q
jtMJYtsMlmv0zK+jyUdr6sa8OXxbsSOQbnh1uQZk66Uo46+Ev2pqfLkeNhjdbfpk
ei5FIYj7E3Goan+e5Uw2FHOGvH5ecdOa9VUm5bpfaxKJVPuCTDt8AhSWU0hsT9+t
9mjQDIbP5rv4QUBje2XdHQMIaWl5BtJZmCrrkBQEGpeCObGma8mYDfDVgi5rkqgo
SUIC1f7GT5FdzyvSW9jkfmaQwCWLCQJEy3u8o1jpXWCqOTYNcWzdPuWTHNF4slZb
efKNTAWqV4cTJ3jy6wiXvZ+BYSAnQzcpKvcMAdL90MHN2IWKHRk1lxPXBu6n+r5S
FSA9qeAuncpS2kxrtQuITu+IVuKZyZzKf850HvWFVzUn1GX8ypvmnuV/lSS42Gkw
6hMkrrxNIdl5rVJis6fQGxNtXm5pa79I3zKuDu8cvnZOrNjRk6laZN56UfnOBaMh
zt6jeAle5ia1g8F/myaCyDWvxPOzKS4TNk5GgwJMVbHwzPmVXeNtH9Q3yK5hAR3N
rnGStV/s2e9rjlvoEcfyeVBjOCyOPjCOahUEIPIJCPrlA0jl/YcLBQqc9JWwKfaa
jUnxDZJFdtcer4fSWxOYtZwQnu3yVnxedK4qArjZvQHHJBLlNSDyoeV9giuQqoOR
Bf+6TpdUqUTq72m04sOjUF50gfii4ovEBh4oLBFsXhZFfRUDBpNuoG4EN3EnwsSK
YpnrwVmz2fMt44a9BAa26i3nYVhxcILAVgvpIT0Sq/9Pb6j81blJ4oKcwuN3Tfcb
k6OPh5GjBvGUY31KVa8emfBxDexSuYpX3+c45Zfa/VxdhVGxdiVWGhYkrGPrLfsH
QOvexAUHL0WXtVuO9aL0bpgrWctCNPGpb70ayocGLHO19XFYxn7gtMZGbqP0r765
igIXxh/u41X15iYMNf2j2H82hf1ij1Fm+FJpQOBjgU6TrCEERZSALp/2msIp5JcW
IIGb3eI3m8Tt5ajF+1kA5P4zFozFMhduPQW8urZNw1uZHIy/DAUTnt+qB7tjaaFH
1jiru9Ug/f4q4f2BSpda6vTyPDVKu9grj7VIo3Fedc6o73APVBDyokrRdWCH5w6D
EYENn3MwCFJ7DIhd4tRwLl3ahyW9HKgWS9WMENs7iR0OaYcIdBBAEg+j0PQ5l1Qn
8ZOW2139XiTxpjUqPlQz4m2nqeyYT3J2N+bC5nxOaGD72hdyhpmTa1vVBe8T5N57
2rP+ArlNEGNeplLy9TJtRnaEIYrVlse8AGpueHJ2HKzbfEBIGfLfeHgqTkcM4SDk
CXOKvwzV7Cr1PTuX3rITT5tCd45h91btwJ8hxQJe3sFbgqFbvlLE4HxU8fvwOx61
AaYC4EzYu5NtP2E0NDg+bmqKlMQ73wMdwSoVIUTKRwJbNeUTqaIPqD//JdXEenan
hO8U9Pa12bEDHxOdjHLiz+jwBplXiwiGMKTR7lY0U1nzMptU4J4SbevsIlfmi2Cm
fv0hIIjcpFSGu1iq5wZet/OHIKq7PJQpT52MQu08jG0/fYI1zgdRnNMSyM8tjT4t
AyCEJZ+Q0g4lqJjVyN4gtif2nLIYgz67AtjpjTmePTEWPXZldj3synzWz/+D6rM+
8zkCTtq1bi+rpzIEscYz1K/y02gMYy9mMazl9jO3+jlWtDMem1ff3AsuCkQiApIb
i3GcaNatn/VjTWWPmuEpw1Fa10CbwWY7i5BYNMQvp/NM0+J/VHjQVTlRLKRSTvt2
3+j5Uwg81EXTT8M+chaHvEScCnojjsp+WqgZYbnrvIZOD2+aZ0Kd8+5GGBnSWrSI
qfd/PSuic6OTFzq7O1juJy3BwWx2jOIMq0W7zyjoHwCOlEQYEL6JYlTw6VT1BDj5
KrAJ76FCuvPrKVPOPXZRUMduzD0Rs8tNuU9ippaj7wJdi19R67c+rXw7Vj8q5j0i
WEFJdu95kexgLmsgjbwt1ERsQ1IPxCQi0CEiLaZKl04tzHGJeyLDVLOZqwNGRzJO
RWm8heERguIpLaDD1m111eLag0jsTd7MReKT9n3W0s1JRWPBnFz0r6Ks9fjM5l+j
SHZWEvnh6qQ6poL+Wv2/QGMmpv79vtIYcuheayQN+j+lyE6RhFgRHAwvPrZVDfU2
lmd1S6AM3OcsK2o3+N7TXQVlSbj2v8uAwg454/69fGSQVQLyob9cLbXYlBa6PK2P
GHHGfVR+P+iY1i1NKc5rK4pk2329f/FJ7M1xH8Y5uFA52Jd1RMhxusdN0fu6GR7d
8E2g5L5JOyeo8PZIyE7L+q4sSuzqodnXNvUtqTz256GdqNlC2y320C4on7JZVPMO
IBXnIdfLYRd7UTNhy/4J9IGb1KvpDVhZKHdsGmSI/ltLLy1/j7JGHIlnC2WxwCa8
yjWCb7OeB5JBYzC8/hjUVPvp2LiYqUZbP2AdOI7ioCe2c3kRJAKv53ka41kse01W
R+5ti6D6V6M5fG6R41STBh36wd5YqmBj+z2DheugooXFB6euIOlU9kpK7BrbtaAr
F0ZV0RRDOiD/7rZg+BvVwr5KmNR/BBZAmoarmpaebcY05SZfLrDP98Qs/WZmrfij
SSDPFMPRYTB8BgDPu8WfDOespyGbu5U/UOCFT6W2Iz8esqtji0GzvSv11TMrL+JP
G3QG/Y4kfASnYvrjBLVdJwBFTrM6a8nCDYK1sUQuietwnGobEDvSBKPsI/pKvzhg
sza2PVhxpe1Lhy1AMSjLBFv2ICnpR+UAXELU9JuYAG1HgHBNJJiL8+0Q+nfD08a9
uP+2TnT6mMK4uFW94yH1B5IcLfaRU1vEA8zABeyOISCt7vv9k0870yvC7LWJeqrV
ECTV+xZy18wSItfThEDQWP1rAN9KexEPDevDWsJ9zr3Xv7piFYPwYiy0vhpTBdYu
T5F/5pooDm/UaOxE/7O+IQsAuhNvqK1oRgDfI3+NupiILy9sY/dDe9O4WXKttZro
n5DG914jwcVzjo+yWj48xUd8OdwJjSUAChF3vjqr9jJfZgqQSEPudfDEWuFz+j5d
s4q1pjln0F7m5a0KaUn+So8ij8QNvW+ak60Sxc3UIUlsnhR1dWvLc83B+jCifHTE
0RYvH6UnA1y4jUY0G2SP9lAShz5rGZvsBpZWDcjpep3sJ9o2q2Nqi+yNY7/0ehNd
vtgqMqRoCygCt/uwCeZSC3l4YxZMvaG5OAJ+3DCy6w3ELDUYVFNCkM0LICX5s4Hz
iYHxUVuR7irF6XVBxyKyb1ZUrW5d3P8gLM+RlFYLxjMGglUfzL7VYPUpubSTaehm
2sc+72FVA6QJqsj3xQqeVIqI6KB3vmAe63gvS5XgRQ+bIYrbyXiro7qyhoVu7aKD
jZ5rmfy1M9dqTz9AFqf2+uRHOww6n6xFuhZ4d241DuJOiq2yQ7VfYHjdCc+hy6T9
OO02d24olhbR+seM4l9hZT+4MVNUWuncYY4QvrInUbdk4FCN9ChbmJDcb1cJhEmz
/xFqYN+0WjpSEvnexKiCbzJKxdCkXFUPMuxHSSU++oc+got5XtWfmdhdAGgLBdJl
4KOcCfp+uYBKrcRwBeut2F3Z4ByX9AE1jRBXDTpHOFOiHtQ9aYADhwkZ/1GOg+vq
tIBe4f0OcDXTD3uaH60yZxHC6hHvX7ihXs2CRpfwT9CYS65kGqeZJ75PFSa7rjE/
Er702pk+2ICg4Xdga7CE+GT/8bkVG1vAc0TCup5J/pSHnZm56tQlEgwMi3lHMPHQ
M5+eCmP/JEr1g0aPxa4a3azXdyu/z73VMCwIU1nVGmLiU4sdSiZHSlgqI0HWSxfx
jCsbav73RXZwfQ+qFt02BmSqU0rI/nZwE9mEcrwLFFa/2C/4DzsgRFdHUKbISWcj
vocnFbQEMHyjv9l5eD0yQaMPpx1RCP1SCbS8BB6Thkc3hQ7sX0czNzOqH/TBQsV3
g+3ub6M5bM7OEfyzdU1AVMegNUt4Iatwrte5b6C/5GrRWr4CEhW5L89TphehdE0h
DoVWJAcnzvaXWLPQHeciFdmK91+3ekW074O/2oVBKDD/LIM/m6Je5mKjptvvZsLe
y5fvC/j/SuzbUAplOG603kw8VHvYQItxC2b9FSRffIt25Kco+L+W04/rJQswNhcH
m7rfcbzg9AX6gBjR8yqSirdQxkz6WXOz9qETceGENF411yZyThVoIUAQLldAvLN0
YWzD6o+JY/kWMi7lQ3xOO1lwF/Wo04jPxCDWL8Wm0Ha7lokvyM5iCnfGy/6L5yJN
g8aAOXQsXWIlSMzDr21dqw+E21iaDjWMzZ3/vHlQ8bsdaXlFxp7JN3syC8w8CJBU
Y/Sqx6BmBSQ7ISalHWomMXvO3HCkDTZWO1TKro/A6ZN0fseCsCJ58ru0+D8Qa82o
+OJVSBQPEiQQyhL5yOpmlCGrm/A8InxHTMK+QkIEUdv8OM65C3o1kea9iD4F7vK4
TAOm/YzBEsJE6jUfaWnENXAUxSJ00IMRSBqJMLbYLMrSm6D7GE8fTSIHcO9/xkKx
tyM9FA3X4u4eiAT6rWEkmQvljVtwnG9dGIkPlmrSHMkR5ZqWJHxmYacUEB7VIGZF
NANr/jtfl+1zq0rjqInbUW/qLzC+ZTZBlcCNLs90zvNo9mABrch/gJ5OKz/RbtzB
rUD0p0C4hgeETIqCGIFVXWpJDr0AVPXvkW4RQExqpLAtpx3+0vqR2qED8gK3b86T
366mZPI4XuCBizTCiulNlFlZIptWQe0ndbVfS4O5rI4hvWwIjW0yBiWvO3pw0TfV
kSEohLUxO4dVKcNABih9SwqzYf/C9TA3cKcI1Pw6Lh11zhgvoR+dMO8b/j3WTsw5
iPGmHY5rXR/Ij5pZo59osNds0ARd4hYhFqy5RakPgVBhlnWm+cutlFzVQTkdlRUu
nl3Bi/ZFwEksrNXAFD2lZGbWLOA4xFGk4d229s3qW9G3BfaGuLYxQVGAo5CIlTGf
o+Pp/UFRrSbydUd7gcYC5FMD0QQu8so7WiLjsBbsPWsM7ZW/0FG3985YBcToL4QD
x7QzquTwdSDyvLnA5cBcwUbiwSN7fsQ5U3ZHJ0c98SxWMI63MkEW3qvCJllPTR22
FeneNbNbV+bR4nwtuf5fGykjE9X9kM1Zuqwg/HmVj+XtIwZIZVGejciW8aLt4XJZ
XTAReTjyo3Zo8zkHP4ScoJ76PoreHTebWYTsN3h1+/NaFeeryhmkq9+MEXAriYv7
iT4FQVQj127En5Tf7EJlu7zy+5aM1EMdyGFHLq5GK5WMCvWydj+9EkdGlmgFRF/T
KctA8D77MBwIe4KilA0XV1BFRMQq3kx/Crg/d57i6MtNqsE9Kk41L9oBLARduCZZ
qp1+sykLz2iyjUemgZwPxbWCJjYl9so/BLO/xaxTdn9/lle44PaQib3tuNAdEBo8
lRY5gKqjuYB4J4UwYJrCpaTcHjSeGvAvvngDBkVweCCUen+p59dW/xmynONcrerS
YB75hjYBZ22htY+BadAmFVtmFnkNx1NpGQzmm97epPE73XCtQHVXIjyXRVUCJFuC
6SWm9vtWVCEvvztpuUCCC2xhqhVxjRQ6M8fU43gKjG8WwQqzRhQPtz3+u/MdDG7D
r/9m7pvKXLyXra6aRXw8i2cWhztVCYrZfS3H5dXU+AH9xNpE+1SXcwoHRMU/QfXR
Yp1co9eHZPz/GHhfh02U/jd38L7mJTzRkT8iOMsHY3eQ55hvO9yD3qmg9SqctgDt
ps3307tqb1YcUqFcyGtTZ+SNE0aLmo9tsmKb/jhydzBxdy++ulw7hPLdxh9YOnIE
/JF8hNUF1ITmCQoHCyv4NlLpOEMkekdbv5Ws+A7cRu9HCD3Ioo/8yv1jTQp2QC8s
YsJdJMM3dL7B+/9zYz37NNudeFy0UeFm9IYyHLEWxnpARqm5MEbNxSamf+x+yF2I
trF0lcPfbckTta028eHI2fYDTLS8g8iy5TTvxll5dXrNj5yXUdgnSFvj5dTqvlEU
UsfcbjgP8kTW7+ZMXv0RJQFVRJGeqxltZJxXeyHTcL12Ip+BzRDupXWjuv3dlUFZ
KFZ8C2vEED9mOg2d3KnhcNpOS7+HMmcTJ6VTdl9bauAEvwLTbi8A0dQHfAdUYROa
bcUq4F+XcoZhbUYZSux4U8EI6sH+fwFMLktg9NYBMXVy2KO/xAKDVwO50q9RSJDl
6QF7V0EC4SHEOThF2Cj+c3OfvkQfPZHmVDvQQKw81dCOORCTU1JOzc9rCmVPU3BU
pC9uOAOFcErKSXXarYeSY1/9tLSjb9fGAttliAPu0XJCVjz32wA+mxgo4zFYiesq
ywxYYn5vPeVCC7Cdds4u0CfqjmkzVcoUZ3TRc7ljlKd5qRleiaAwk070/bJib0Ui
fahStbYRJ9mt6ljdejaF03Yl77rZkRf1FHoitj/y9dLes0nabjcG6VYZP4K4cxUT
gehDWO9qpR0vCYBhb/mcOswR18GNZlf+wYLILiMQ6Cwbn8PLqts+PC0EMNA2VRnZ
Eb/AlwpWT/1R8wQGjGpudGaqTLi34TPe/nvnTyssgvw96eS5TNcxD5XsYTQJPoma
z5RKCXOKKpshRzOz8UniL5KXxM7OeVnhlImdw4kW7xlYmCJj4CIMrbbqnyxoQh1W
9XhyoADRSlsAEpl+1X0UkutXIeYhqlRZQgajPiULeGLqcJfv5Gupf2VRlRcRLp9s
62EoCywHFntnWwixuSlZwHlcgG8xbTngKQ2VAMNo/YlpaB1wPAp31LOMmSpK6pUx
L4n7/B1PoFGPn9GnOnqfAHJrxmBfR7A3o+ASd0k7lGk15IRgXIaVvq4k9y8BiJHx
0VZ4l62l2pqBi+KJHhbmy9Pi1GXg45s9omq5wytSkbjXh3FJiTvpHhWNWJdFJNtW
BTFgrVFCskZGGH3o5IUoZae5/8DMfkJ8laSkVVEQQPJxSrt1vC6Q6jJIb+mcUbyx
jbhjE8sXtKVSsmhiRmr0H3Mvx52G+REgbWXSWgFreGv4goBZp8zI82aerUanhwiQ
i9BJlFdEIW4QT1WnVHi1dUHrt/8uoIyzGQgrxDBEijHln+gt/8zDm8/KzN5jeTao
TYKXyk8ohSlM51D6AuNuAjTzQWc6/TWCAdssAGDQxBU164wOhWAkCJ+mvTnpxm9W
CUeSiBA8taIQpGxqQb5ubvMqcWOfRpNtP2J7Y+Vd+vgHamRFBOWuBP07PtcZk50I
bHJ3CpyIC+dJyP724J1KVHqqNhhfZa5ET+wH1e7XQypp40HdPwJNxk3g2htLMPLM
Eg37ozZ/xR2fc9r8SwmklMqPI07jrSg2hyDD4xa7u2NM9/hKxqBJwNEXaD6pJc/8
UfAb4v+dm26jmNychd5entXQ/bj/RRHvB8p1DbAaJu8voKWNt2BmX6I6VNFosxJ9
UDtNAZk4UpsDqE9oww4V8GMGxEDaXXJValE41V8AN50ooSaNHrXTAqiO+mQBZdX5
J/onQYiPF5dMEAHSTzfY9oTfgyTXkUVshtnZL4F5rj6k9UhTOAkZcK68JUKD00T0
CiPqNu9fkt+ULNq6JxlsnweL9HBjRxW3QzUgLoFdqQrzKFwMWp3epzKaUXM1wBG5
kbt5DasqDQ6q/oIGzQktA5x6a0gBhhUU0nIHNyrNoZ8+cK3VDceI2kIAY/zzvrrd
mKSS4Q2Zw1DvDJWykvHxytcU4KSkixiJRl/CuM1PDyxvr4nhS/4zEAB+7wnH34i0
4IgGcJMpgpMSVVfC71T7P7hPRRItQUwW0VkC1pdGB922WnQIFSTxQYVmzTEruvW7
bFpTf/4JKnwfOHo8kWxwUj79ABuAe/NCtyOzoPiCXD/ja21bNxJJ8ZhC+IYDIPOv
h7lQyl0hGVkJ+uNaLhUMQDJ3W6SeOtB5OLD7KG802JmUMcyagUpdWxnPrHWcdXO7
6ldhj1/rKD2zCxkpnRGKPXaIJaeaf9G14nBwbs0usoKocfvnx5yX3NYntVz3zgVJ
jOcoQY9PkqfSlHbJWgkc+0BNCjbMyj97mZ4VmCfMzemkLwTsIGa7w5+GiVK5lO/B
eE+XXvLGevTdZ6RSnjc7u2DJ3sxZyYNNtzCZqipNbUl51g5YWEcBg/JFKqwZrbrx
UgsH8k1MlpGaRoKLOTQ99d887SaqC8huQvTIfr6bTyjtn71/S1XU7pV+PYzWMX4W
M9+DoxM9DSFalmm9ve5m1O/pkjmaJej0mW+2v3IYcZo67z43QupGuzq+wfF2RkUQ
Pq4Mg5DIdQUvqgdhUhLA01JP/YDAcBaVkMi2DAmiUmPWc+byRLtlaDPwl7/poACz
kaOpqtFWCVSa+pIMJQamrYyxhykyxIxy/RLvKMFFmaQjnr5MoiETdXcqI4IS3qjW
qbpcCLMun2frsMf/9jPIXLpq/At//bD42L018Tr5uy39+gLqF5OH1/H6M/9cjnlH
N3i221u82LXwedf/ZMNEVaS2bF2EzWlRKs9+GtuxHCkzwY4t7gIj7U2vWG1N2Prr
wz4jwS1Y9DT5mVpxGoLyAWfzfTdKPfzuPU4X5AFvNbxxl9UTdg4PD9oXvPmODGf8
LNIdyYeKuZUMPxW8E8WOa2c9WIgRmX6cqve9cdbrZauYnfq6J8e2taSJcV0BvA2W
TmTIdEzswrd4l0vR8VBEz8F9OrUW5sC6/dycTamBdz6amCq7HPmUo+iYb/UsqZgr
fzCnZqWoU1XYXR++CWwC1CXyBLUL3fALLBsuVFFseQrAUbQwlfvYJOYaybMjPXZJ
4ytwYqBUX90vQBvXgv5ox5fq3qagJNGwaMhRlhLkGkHXVXQUDV5OzNZJNxr9mIHf
OsEV0U03Uerk/lzdyIZvPTStG8x4mSPw+yf49ONJTDX/PlQ6IrmMjWHYGDMasnh7
xcxlKAb0J4TmNA6RT1xrwcU4bNLnRkTX88jqJrZbXwln1flfBpmQKtAVDTt1roA2
yvKm+E4Kk3rDkAwrDAD/D/yl9P8xePik6fqGpw0OThO5y+1wUJdfcefkruDfmsvp
EkEDAU9/D74FSQB3g4Tq6gWlt3b/P36OD4TnHoHAPFvE9+p6VFleb+K6JJJQYQnq
+NJFvhqDfapQznUmo+BAAH0qzojl0KU4TevBSgHopYXX7HctCvMSBsCejUBixeQU
cAYFC1ZMnfNPs5VBk+GnDUcWuQV56tNoJfhv3UucUPsKN99WjIrpBhYxXRBmVlEV
u3LpA4ld2yHpia+n4Ny3xp+eG2asqx6eDRlfinPgPPXSqOb4Pt55bRPymXL4HbDt
wIYR2O5t2xatlgJGt7TO4AQkcrkFjcZKA/usQabh+5xfun7/Ky8IvO21aBXNMie0
CZk457HzmHVhOf7aC+vQfPqWgiyBYH/unVST5SxXcR01NFZJlYafD+mFy/r/fhOh
uCvqg73L1+iXbP6B4F4/IwizUOUwZWWamcZEdEz5eWBHNgGULW4KUJeYI7kpAsR8
+yGWMqqs9RglgQFvyXa6RCx1wautQJ8x+AHZLQ6FF5FmG+cfr104JxcDA+za3ZSq
RBdigySQDJCp7KxO3mRvfObeVJyks00pDDXW3e9KAohtoOLdHxtCO9aV0FuCaErK
49BFTIrEZt+yKpq2pZXas+9Ypl/WJjkj0NvyIu79+SLQjqJNhjKXEW062FSm/bDk
9OJ/wo6mxNe1zRpa9Ta6UzSQZptM38aTf3pA8w/CaaPdr17XL0EPPZeWDYVgCXt5
Wkx93JGnJoSkcCKn1ovhdKTjbfayt7TovFgXatY3AHrXRvnWfV+5WKV9gudsF07m
yILyuH9JXb6KsEvurRXcRLaI+HIzPqoSJWkYwd9ZSU42BaJikwDT69hIBWHNfa9s
LAMs6fcgJO+EPN9JZf52RZcqmD6OOUdl+UBXAUQ9zYdqdMbZdIz2LV095Ae1+bVt
M1VIhLzLhlm6MghsxzQ4RApCkwiKBA339pQwHhQwo+6L57fdGl29QCJh5UdZUz89
gCLoVwmhrBwNhcHWsmR8C4o5mi0aYX4RZjMWTmMQfzwfYqDZJUy04xvvCKiYMFTY
ImfnsGuFDSMQrODSHEYiAv4eKYxhCZx+aVRzwYJCilNXWbS3ka2/iHqIvcRkV54V
U18quKcLytR0zAYE7/lVQfie5CnmhW5v60sBV1T/EEE74Pn31J3LhUzyvoToTL3c
fsrpoS1bNqSyUKwzLyGxp44ZXrw8bbl84m4qXS1RvFA4iHrChkD2pMS+jfoJWR7e
EfFo21+Q4YfZlTLpw5kIK0AdwwLmKYDHmXCj84MSiKJGLliuiPrMdXmY9v2FEtbQ
Arqj+HxcicWGA9bm1ZzIxbJS+9hceBkm5UguAhrNimLoYWVxOMMWFxpkOX+U58dg
lDoOLXDOaKMGCBOCL9pKEGK98DeF8fYIMJXVRZDLzps=
`protect END_PROTECTED
