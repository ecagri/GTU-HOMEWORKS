`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0zTm//x2nEX5tu1N2+quLJNyfekF7HWSxot9PE4+b4kkOIgkJOhz6Uoz+eZ3qSxu
oKm7qFddKtQzs4S/PyttRYOc0mAFjnL5KwJr8MiSURsq94AhPrb/d4C6IqK0/wsz
OMf9ORVXv+E9zVUgqQcAOngFn2YIeSzdF3H3Lpzya17CWjuaKDlSym1Dry0gyy9E
UKBIC/zh4nYTKo5LIPOYcqi/ZP3cbKLwCtQstVkUNt+T2nTnoMNtrJJllo21pIRH
FrJxPo+1nG14kYwTM9t7RZ8s2KUWtdO8pzZyb/F3BciJfi41WixxWbolzUkOnfHz
FNjxUt6vbHVZfFGfIr8gmDJ17GyUNpXpbh8wPJ5GYiO0GXGIVsnQR5K40qhInkWT
UA0gktqB3RpNVkbbseBJqpPl700KmtsZj8vrV8ZBA8UgG6PqkjbcWZzyd/rHDQQ1
GDbUNBGQoj+TEfoCpm/6QzQ/veP3ATcdbN/WgqNW/2OCLbIOw3Yk5WSyMug3bb72
mz++mHDrX/IJiVZwNkH5Gfg3yTUbqdqCCMSn8IJuFzXyKFFbUKiXeKxaRpcCkc6z
ZU/9uo0rla5/0TAW3toogGzvQka8/nCv/hiOBZ4cPgMo3D+AMyxY+jLwtO2Onlon
06KFcCj5Whngr6IRvlB7nRbOz87CdLRFa0V7SuVl7a1DtOJf7U7cSJ20LzfBHjSB
Qq5/VE0h9D0GE1sHaYikduwynTIk7xKWEkS2nF8ymXcwTX6x36VLJj39MVqHIxF0
j+RPwg7TG8niR2JyuTrzoR48wueyMf5jEMLKeNyIiGCUtC2ZsRF+5Qe8w1cuFCY4
rHkM1Rzk7p2dBO1O+vkQCiZIQbmRdd7bj0f+txSmlkk9ElivlyzJv5AvkyA6zUna
mMOFfr0g4+43CsIGHPL585minF8t7j/wGdSb70+FMhzOnDI1jhe0lqzZKOx3MTfZ
m48c4zHFi7kj8CSa650Qm1PNDOkyUMWl3rXDliGFyQlMMwPZ8EKuYl0eL2efD8Kb
gjf52hr0+2ZuYYP8VLgIA0EC4+JYJJwV+X6W4ssHifTAiyjgfUb2njpokWLB+afd
FZgS+ovRcjw5Ybc9cPgA2H8o2P1/atzsyO/0pzE10uEy9gBHg7iEPB/QZLDTHNe4
rIlVL3orjDPSaT/fyKhouTh3yoMXAsq4DUuKz2paOiOfCqu5NDi5KG9i8pb8d4sI
rT2LzIOyp0ggw9Q4XFJLsNMG0d/WN9Md5LyFrQhqBc2GrQn6JwFBbHasWLoXXJzI
KFolA1uM4wvFc5S/tlR3ZsoZj/NKkeeL6glWPBJoZzgLsAYdF3lnrWABWQq8+62+
O9t+BnvQ7G6hmOoRJidagjquM65p+ya/yiJZ6cai1h7zmTZ7putcGv/SMtICuF2K
PEsGCjIehIsE3i8CHmuFuvc6pdNyFFP4b5IwNHR4uNTNXXdLvXwbagITM0aDwRqK
5Pu9mgS3Q9AExGaoBXk0OndSP8IhWrcD/JjA0shmkjoL0IJA9EsjNUrkOfY4BUkR
wg4DORKi3wiSjlL1KgrkuCvjem7EmlfLZeUsDbrPZPRXlixsn6r8wONLjUA7XQ2q
t7udpnWj8gThltpz7+BUCtKxjtnfjwdbh0FuGE0yY3hkljpZJPJldEMf1spARnTj
FGKAdR7M35Vb6wT/FItDS4UI85IX6AJvXFIBnwBe64Pcic7B/FG/x8gC9pwmyGGM
8w+PcFvr0FTsvC/M7uufyA5vwM9IqNNGnKIwPG0/q08/1czHqZBWroWb39G/Hn8d
tPLgD0SURIpRRcL9uKaxjHQ1giE1NvPxWY6nXBT2E5xKvFQes9OhWSYxffnhKrkt
uI1lcL1HF9E3IRpFh/U3glznafK/r4wEkV7Uz1x2XnAW9IcAYBWuLl4hrQUcsyBp
OgbCtF8jzxWadRlkzKn88h+aHKM40n78Bj9wx7IcnGix1cxbR4niVTAUw/QsvpO4
vOMg2121lMDgf6Xxjk5ROUArPOc6U99EZRg1YSCRGZy5QEla+eKY7WX083RMucyd
90bk2+BN78NgGPQGhZ2bZzLVnJe62bCx7rBEBY53FcKCwWKn+I3dbQz5IhdB7erj
Omr2cF5+FF5iSsIAVyEg6a7kVyZlf8WVwYSTsSTk3e1IYQwqdnF2o3S89tE5tx+F
4DhlXdvYzk2JTF+yU3VoYWYycsaZwWFdm9F7HKc2NE+EW+EgheLEK0e2W643nfNu
cBO7qdffNdnTc4s9Y+Q3kCJ/lPHQM1e19g3L+8jAFynPaeBkItX4hChWOu2My7/t
f0XbXithpnFqrRDu2TXSvT0aK/EMia0TUiP3eqT+YUC2R17YwoQNc3boCLpbumOn
2cVLV20bx2n7md7jYjxEO4eMb10FaTh95vAuFboHQsgXy8zymiO6eI0GZJL5hYHo
q65JqZi6GQyzvvnGgbYRdqyAfh3/cG+h5O3bIKqngJum2468V4cDbCkh3gU077Q6
GCzobQwZdmHabpM4JpA6sb0R/mH/jJvIPIeuqxqYVmWXufBE7/h97f4np0iZ4o2w
Zh3K+3/u9oO4LJ2jIo22iJrAVM4fz1hOJb5Ynes70H08E72tij2/qKcHVmrB6OEP
q827h3m7QuOrYwwoocuVWKY7y15tHZiahp6k1YunS73fM5o8KUW2ZCf4lVjZhdRR
BjmvPMXt03zWooJljywaMoyePOIfnQSqE9hJgYvPjbfybrqoIqv4QQuWe4K9ijcS
ctCjTFodTyLlv4darhrP4piPBWA8u1+DrnO/K6bcWch+OOSMpzrIA91nV2LKacQL
YNjp4lNchvn55iip8Jp6OwIvazQ0/XexACG4KNZRpeRioAnkoms2uXPRvlj4VGES
F03r079HtM2KxIUmP4MgLFT8sGGDSa/rPB7Z0c32Bic9LCAFxBCwju9K8XFF3COj
o3A+XR3qqqx3KKSVOiJ8f50NkUgYXLqFSoEitZpw98HvEDu701L7F2sZLjS1SixV
YfZPUdSlFoo5cGXKZrB0PiLghQXp3pXzJtTtL1a/RDROnYICQapnChd/wP06C+Wh
kBKW8/6Z6BHhWJ32NaA5znQ4YumCFKyep1WhLjW3e5QVR1OjHWm4TnRuBHBMCjyY
qqTV1W3SDARZ6gzMU81NPa+XOogk7S94tmHuxq1zl8gWVmqu+iF71faap/RwZGbL
iAXb48OIAjRb7+nRKixm4TV5OrSKjW7PlgzimaQ3R3lbe5vI7nFiSqqTqCHdkdbH
S0bNa98fgNWJoS763sPbZj//TysOTrB6CS+FHG2jQx/D1HxJ9l4opmA/SJCNytvI
1GligeBJCO9Ts/+LAgGgvulQm8XZMW8/SNqO9EJdZvm5VO5mmdyQnSk52XjAWX7e
d6WQPf/2axkUdtY7QBMFLkqkA3FwKcJRiFKmYTqHPnODO1e4ui5OaKu77XkQYIdX
Jz2kUHgfmbH48r4TSbZh/ph7W63V5Ivj5vHcOxanmAABPrByBfa71quYk6SptAts
EaWswDxHuFD/IgotDtTuhdKjSncYwVd9SDREeXpeaBZyBRFRYwDqYnHP5xX01H7Y
GV+uK2HiYrDuHp11sF52kSJzEpA9DA+08O0txM8HfoGlBuO2AHhzzGGvESIG5dP/
Za4LY+aLjTCR1BP0fmOk3DCXPlbfAts104A8G6mZQVFGR0MB+ZzBQR8nHpSVUuIJ
2m50ocknYWs63AN5a6lTKtlW0NpenKcppSichQHbYeaNdRqRxNdRBSkuQfSkHBVi
LWc3w+VX0L3++sQ5LcBv4V9O+fq6PZFp83uTyO7PSVjPI4PdiSAIFHvbrNgejCF6
Iz6pSYeNdGAD/njYpFQwU0FS4Ykg7ssyxZcsCX/vaWCNJ8N6be3aqcT7ckWaMv/p
qGmMbkeTSK7A1GrQDanKj0WHmCPf+PD+/RtHoIyPYudsPH1TmV9VA73Itp9Yfuji
T0/ZZtD+VYIDvDNVkzcvU9fuDvQaZNZ/YNuNDjuakI83kvQ0+ixYh7oDSCqcj0VL
Wep+sKcyrbOq+vy4FmujE6EuLL/pRJOE9CRj+QP+6hWtn5+CZ9oKMWqyeE+L0ZPJ
Sn5/IVaMTipgD6Lg0ShXiD/5ErjhKDp0Qp0qRfV+VAenckZpud/l4lwBAHd8Kb2b
wpuCNuM6jDSn+OM64Rj0oMTaTg7mfeOpAXLq7O2GAkN17nPI5YuQA6PQuKqQjzOZ
Rhh9xb+ckhIiruMXT7wG0S2zpbAy1ERm8fcv1fZv9SrpCi8gELy0rlh40LkHFJrA
BWEWbahbY8ZVTSU5ftCOsqLkMx07sFz7ky66SZk7HeYDMlEY5liBVxuRT2ERO+JK
T/QeJrh/gAoC4COG/roN4NGp/xDvI/GErH9hI6NUT3psU9pEuvf5Ycyx+Cs5L9Wd
rpEvEHsNQiSZPitLad8e+Wr3L1SydAldItm8/aTaJ7OhVw5l5cZLb5OMlFHYUKxA
j6pND4PZc+BwOeMzy3Eto0pUJO8wtUWuxad6w0oWkudecDEpitELz2qQdXygsRNd
+kp/rXCzUIskqu1d+nQXpiPhi8mBDQ29RhEI9/z7YDQytwEyAD7Runkw0EaC6MnK
rzX7UH/ePVZU/VsuOaxgLspjMAlsBU0Q9IuaFqpEIK1VY17M6lGF84eNqo50Gtsg
7n709f37nIpKieVzp2eFZ/PeK2Ldf+2qd2NgKmxN9mxMtv+FbH4B3mD3ADBTg0og
GM4/QwJzNVFNnFOUhm+rbiy8pdZxT1mWCdXjUFIb9HXoZKLeS+kcvauQcQrXmB8/
x+6J0LA+q/OjPp5JGezbQuF990sACAN43OSZo6KZSJCkq8cgblBPlCtMDlo5pFva
RAq0ueUhPwVX/YiJ0VKZNkMqwk6Rt3xPBbVkE+YRsgpwM0EEnAWxYmuSZVVZvBav
`protect END_PROTECTED
