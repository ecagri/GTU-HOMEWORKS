`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jB2OmQDWnUtrXy5OdyfTtFg6eTmTUtgWDtel9NYFbxIIZl1geBocyKoUPRSQI7oW
fLXirtTmnOfhY1/qWoxOFeVrdr+NrXGiEx/AZpx4VZnPo3KVuXkdVHeszJSLJ/gP
PwGk4lvv1jf4eH67u518JelQY6cu8d/0k4xfVPH3qg1Z9e1pfJcfhE4ZHqwp+OjL
UeRyDT3QtfoHgD0Bdl3mv7GStho40trOMPXfULkzg6LHXsFrFxbrVYYtsndEkzF4
HKjJome2eGlp6NCB0hG7cvTeNTwH+q2XlWefWp9ucyX9csYsnHCQRqbJAj+GAIMY
+tUnsXy+jFv63RBaIfk7QeNb1+DTT9oxpFuCC5JycMbCBrkIgsM4hDHLmXkENieZ
vbYTfoNYG0CINeHT1Ij630m/P+Z4tqI8/z7pWrgbZyJKcBuZ4iU1AyXc6l8KDHJE
dbFmuSoPh2hVO6keFHR8hPs0laMgAENROheUkcwrAm/sPXgb9FS5vUshPA5pTV3l
GDdU6Y9l2VmLkx+iN8FWueOev0ePcvluPoGoftwSx7OsLr+OiDBhlt59xxi1ahNd
5K1gbiXuNZOaXC6YtcuAU5FUiaHyo4QWDqtIqlJ0PEj6JTE/eEn02jhR2HWcgqlY
+xms7vQOKsHkDBLfiE9IfCJ1pJJ1YY6VAfn9/sZ+7JMmhB5y3EkjIEtvIeTAaGPY
TCpOrJmGNz3SEBR9KDkLPMbSGSmikGM/iJqkXGBJL8GjnBabebPkE/HL89SYDCEp
uOgnyUJWHxOTSWxRZYr9D4xHX5O4SA5EaJxa4lophXeWXRQj1wWhLK8QpU8N5reS
FVmc8/Yx5+lSDFtH24dwlBEXTrFwkgUkhaokAkaybfpgWaoybZ+Gz8zcP46jKzZc
DMqXGwC4zwt2pVMwdOCGjn4gPe/mUy1AviE7pJa2bR/oijVqBD9aCZS/P8Zr106H
vvxdqsAKv6+daTs+dJZ9F6BuArd3BOYvFNV58ydwapKJAiNmzIynGrFhYYiHNjoA
UxMBb+gPVdP2TMSaVfw3GmpsRvRlb3g+90wF7xutyeZ8Of4Z+XBoNZOabPG5paO0
8hovfj9VmjC2LZEWjNwsfpnpeTR3TeACiMkMwfeD2cWlFG8ujowCqYo8ZCnohBUV
steVmiHVM8iEKMH+HWzEZs1gSnJqxM9wZfLOmvoIP4D95takQDVSOvilWmFyDEss
nC1YQSUlBIYvPz5BLqLjRjfaUV1JPbrVkHY/THP7dDBiMPR8GIWBRoWOmoT3vHib
ZdncsshpJ3tviYf47F+mlk/xS8oMrM/xZlztEqol2xf0BdSj48wlC/EyHP3mzbJ8
koQTlTgOXmIL4IqEO9YeFNUppQrm/TYsHGsAbFmyJhh4hzMu7G//5i438rgP8KjA
x1wg7KeYnIYwOb3kcUHTby8ruXaW4abSbQ40ZDeY6JWbGdXthiTdfXo/qn3Q8vhd
WFlFNG01AS/WawiRz7LOPzVnAo5/+dcrMJgXc0NMOKuTSJP08xNjf367EpL6fMwx
IWqR+G7Hf+S52545+IPL5+IUdJt4zunHi7aku0ottudJPtYN8FNMCte3H3cvh0j+
BsuCuM4d66i+N/dpQNHZldUVWItRo/uu9OGxyj5OnivUvKv578mK8gF/iBhi3FOV
DGQCmsA1rkvTqbG12q31/ajCED+CijncB93iBLagRytdFqzVUZqdJD9JHYnCWgtM
v4k70l0fuh4Gqnod8bc4hSh2LvKwzV8b3AMAYgFkZ8nG6rUzuj86JOjCsIRoaBn9
LrxCzps/0R+G/y0O2ZhoZx4GWRAUvyVH96oDL5kh6zekfQK2iN+bIDZaIT0je/es
7VmFuLNy1VyuK9N/abihd7HSUaqyvOvxquNm9JwHpE/n2YITlJKsI646UzV+2pLM
dLqLBzAXCofQfmtnenD9C7Ri5I9TueXBbfz4r4uwbuz5CVYKQX8+XvLkknx2MRV0
KyKq7rdfoGVMSdcy4xQHcO7TgqsgCKY7hp1/bPmHCYI9OvAxkT/Rb9C/gp4BR/3k
JAaYWAk6daLrbrcQG0EoFGRskb1+33v20AtH1i+WWgoGQ1QVXl559CqqZtCXhfYG
rE4Rs7+v1HRP9X8OeAFrZh7i3t8Fo9Tx6ogYC37f6HCeRP51KfirFRJvW0H+EFMJ
K3mGkODn1YUgZU/FybQzwETkQn1Gab9N5UxuaE3dAVonIGWq/Of+c2zPHLFydP4Y
agyOyTrMDcLlJpZcFOi/2D2sAA5rGtyRh9Y+81/d/ey69huvv0mP+8c99vZgTxsd
G7lUnlwtxFvAU2Y33NPDCY9RjtprTyMYA4Xyw7T9o+7dKUsdurPjpdpCwSHJJPiW
xnm7mB5j3nVjEMDIvvBfBlN60a9IeD7kGn2XR7QBz1UGVBpbN5hdPfn1u8+1ccoZ
7QZBIW+hAEI3hT3fdgFygDlcFiyWaF7G6OABBTaGt5bewJQHSaaE2r0VQ4/S1Sa2
G0Rik+eKVEGn1egH+PRkps5z558UQMdq3aLjov+oobq8Ao6J9wK8LMaiYR/wswUX
MMayRoWxN8ma/Q6XjxgDgadJPzRo6Wg1ini/CJnpFbaxHpYMfPFwlPwLMexzXPNt
pneKdW120qirqbGzyqIc6v9ZYl9K8DX987QVWk5xNp8ag6NprnyA0DtcvW9mp7EN
UjdWj6ByB53PGSG+6wEyrfmcEymkOE811UQHpMPbz9ADTQb+EMgR/v9+f668z7Kx
HOjmuNrVApUdn4hGcVVuT06FhExE//SLs1RyasEvdZmEJVRwnMgbOfDlh5PkvJOZ
FxHcB0THuwSXaxFG1jJ1m1ZSyaPovggH1+DJ4qME6tQQiPhsHst1RO44B8pK9BIG
w9Di06XDcjiNEziaJm12VUr+g2CK5QEyZFroR2X3L9aLMzixqKIbjSJLhU+uq7Kz
xLHLEat8ARSOlt/WAt3GnwHJMVmqY57W7w4PUT/LXd3v0oZLpsXZoXV6g9kZ4+/w
KDwOt5poNPaU/URGmWV4mZ3evstcxJNjDugqdMUhOpcvFEFQ6rOnxPsql1n5YiJQ
0vkF+eWmhq7BlXx4ttMr/VmwC00/p+32ta6Yzizx/gOOG9argVmAx72qaZNhd6ED
LOcDIXncFQKufqLGkpjJKLEF8rICKMYmvktmTaQmhubNcx65nlYYjZGA02wlgkzI
EN4uJEFYowOayijeMDLOpValgxi15b86LDHv7fkUcL+jSKc8vYKpjwpv/nBTTKEo
tXQRwLvGCuXPL7WH46yX9XM40gYY/tCDdY1ze87rjcd27U9pBK15VWocIQF2b2bW
cTHoK1CiGT2xIEoncf/w5AX/mckRn+udwYd9YVHQvrYpgkLSXvYmqsRCtHOpblyG
fegXuKCPr1hy78uZ2Vo6g4QiiVRczGZ7Mmf3Un1vuuiJsj7Xahg0t4iszaACZNx2
BIV76lQfi8N0IqZ9g5uSCO1BuEY48Xp1SUEWIFg9fMe05KXNfsYkh7RrYIorml4f
xqCPENIoXb2oO1soCIoc2MtjuJFi2edPtUgn2WQweXWUXQ6QczaOGm3rE6ZJeUxL
GvrAnShusdPyg3bOU2T70kHwGif1pUnkBhnDp4Ua5RkoT6ub2lxm9ZRnJ1RYGv09
WelU90wpFeB3f2Hx46pNC924Qio6cPxKIGVGByZxXe9t6ZLGPxKWl58xmSWxsZOY
aUKKXhGE+ChaGvcUFrse4SACCXYxi67OuC5lAGs9RSb6IiIm0GUGz0Px+ooKtlj1
XD3zylVR4z8uxyF57fEsMXu1BpWpFlYCrt2QnZD92McFBF/zYBsPj9x8xbwy1ysb
rwA/FEwMpxiiDjrNyODcaQgQEngKO9aXAYWNNHXVPA6KbSwhNufXRE5E7UcDmZhO
4913GTS1z/x95v1q6ZpMUuAGvzN17KlDvM9A037SM+s6m5xHdH4EiDVGsjZEwiqk
WJf1l0kYbO5/89BleZjvB9gV5yrwG+5k7OhK3IeqUGhCbYJhpsjR5BqV8/edHEqq
2j4IUDiqGN493z8p7bIrklYTarlDOLn+6Y+ED236BlLXAgQdWpPom67ykyd8OFom
e92LGl7Nv4nBbvm3VgA23x6XsPtADSQrEiwcz49fMRp2Zrqf1sZfl+kDhL/ihEa+
dnEgXrD3sK5LLKU3XGwvACXUAHkBRKnKYJUccgoxh5+1YyPWKUFqPMooMO/JKHpt
Qpz5ODW7moN2gUU+pZ4zepynsnijb5WFz2O9m9dHtB51WiJFZP8m/esUGA5EMbFh
DEKPx+uFZe8lx7XRvThhbBxbsIrg4qg95kC+iDNIgDQDYBkozOvvhCzyEPV9Q/w3
XoaHaGd3t9pyom+hMAyehuvTmWd5oaS+6/uo+B0V+QcI2/0tMjsiKDDjSG3f+kDB
YuqPAMmmyld7/TrGRq1NAw317jjlNXfHGATl1X0UcTtYCa29I6rGPOAO3DLPcl+H
VCtcKqui2lerpEmhvKzifHCYNBCbHRSbRzXiDyYf43Tr0j775MxzEZDBgCIbpnQZ
o02b1EiTFaKtXYihLRJD9sKm1uczdpXwJH+Q7kJdrNRm0q+bKdAZH4yz2VTZEhSS
ULUE5UxG9MExv2ejPisXZ3cwWPIq2enbfdgPA5Nxgy9uemoS2dGySkNlgphB9Uqm
dEPWaMCb2uBq9XmP+Qb3YBACgcH8bUxvHAMAMHyQ2og=
`protect END_PROTECTED
