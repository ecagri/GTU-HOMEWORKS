`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4QdH77pQh5rixXk9lsjiujtGCtjtkJdGHNasH5+4F+EHlhP4KLzuSwWr1FiRcThT
tutJdsrSyVrSo/p2bnBnptyoVVe1SOV9PR1A2NUglZlTubSY1jxcSVNDcFXOO/Xo
aDdHOrwVWUXc7+fbN5MXQOUb18i+yFzUEp9DUlSBYiw9o1AR3g+Jg0YOGQlDyPYs
zYA9vKBSCEwfcb+pxXxU0U2anlwfYVdxFJ7euulLYiMXZKUECqu2qhigvcoOdLtc
ToIhUbvj+cB260Mt4dPW81+blIjyddRE2v2+fp4E7G/hXD94HmqPTljBg5xfeEue
iRosXuZeqUJkFSm5KPQaVeF4+NAWc3O9Q5Jd3yGkP0hVKrE+SqbhKjv9O8arGWmi
HtFM87BxasPRI8vzokV24rvgwea3wlKh4ZVPiP35TaxJZXblY4wx5YfoYmVO0heS
UO3Ws4RtMrYnKanV+ruIFB7+DkAfkZFn4zgERzktPApWZybXh9jMhcefQ84SKL6c
j3wbIB0Vv+nn2G8ViW6hzvTq/SJesrbNRWmCDb3oJseBUvbFxhpSsmTCtbrsoUnz
Ed3mw3otWrW55FXM4HBGIQJoSLOqaKHf3cKPfPxOBwuD6Xg4Hyoy2VgTksmwIPoc
6E59eL0X0R1DfyJU9MibFnaJipmdBzttA+ywQZl7nZRIGAZ+yDjlhSR7EAqo7b0z
2tYuDjIpi+2rVKEElNR+baZzuN+h0moLOWDqda7ZJKnPdeRIfIaVs7Cy3Enr1gj6
Lt61CzLTPozUXjH2f0uOwXLgzNDOarzX2sahOMQU+g6gUFwi3DIvZas+cWrds+kR
+GPPWchL84njpn9+9lrVa2FHRRlnjWrR5IbWxS//9r6HMvuasWEpG2Z5ACtGw0sR
BhxAgvqbwG+JXkA5c8u92l7y/v6VWgS/QDCOkTe+DSQG0hdmAR23jKPSZkk+rIx2
AH9Z66RM5yrzEL8mDujok+HlxKr/hSy3ISc3gP8X4UtKvTzjOUH6mtCoR/WVRCg3
97sbW/iN1RW14KEOiauGDOx1szZmjSfhU6xH5Q4yMAL25W6TtfAHU58QYMLaFkne
tYpyIJ2oG482JOZBWwFejGO3DmYYhZqGepZwxgI1OxexImv/ZYiz1oPl74/gS/78
GOeOeB6Xh8fqQFxZHOFCaDAabD6v6pIIKx8ZtuZLOZt7Qi2h6At9c+bHS9Cr/jSO
wL7HL3aGgSrwhijeL2InSIlRW12wutyo/uSBy2ha2tcMhGW8rNeEcmxmay/YZMyE
+4Azh5vnbzvJd4yqgGbCfXOCCsTDkIU8zolCGR+aAhAjVT4uehvaH8QflJUWwFCF
nYzy0L/9Gn9GQ5ljxtB9aKd0A/HPv1rfbvRsGEYoJBcTI9vS3ie5KOOLKDoTMWIL
`protect END_PROTECTED
