`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XzSYWvt1B7ZXGSD5FTL19Sf1m+n4Iv2+u/cUH1NkE8yqSrWXM++OwF9DL67A7vDH
HusOUrTC98YrYfA0ClMKz+GjkLpySrllMA/Qd/g9aMH+y/MdmthODtWBzG+l49LW
lLjsBrWIZOYr2MpIovzrid6NOiV0ge8XmNu7VxxSW5LEmnTEAD7f6zeFrHrxCxpp
H4U43ECW//RnxHimYrIUDJRlNMAe2bjixAMxpq3RDowEpBdwyVe9T4fysCWVlweC
Yo7tuhaUBeI6b4bL2bXUFSeqAVE9B9Sjw093fD7PRUhCJhJazF2aQ4buZLqdREeX
Ccn4VxiqA6stqjued9byNIsMiLMgeVLDFh0Oy9DQZnUNIBSxwgAGMFyFpqDgbJ8A
VNSznZsk5G5xFf5tYjKsZHZoLZ9st1zlfbiqibM2Pi0LMOtTR3zXRoSXtLrjOwZD
9KU0uSXDZqm2y4Ermot59yP3bqf/jIiFzy7JB24lvI/cclhmktPV02+CtPP0ZeXB
Yj+eu4WHpKCPDxssTIvqRfVEU0/UOS698TBSEedymBG7yAF3PXZ1g68QiBb++aAc
fON89MiMMiTcGZmMY2FJIbe+vVkusODXMrfIncy8KYK8aeuXiPvdopYmcMAhnyKQ
UjKV6AYcK/wCF1tGwCCDEGFI8giWCmN+eZ5DPXMLa8agGXI8PsKyRzwHepCugXnG
`protect END_PROTECTED
