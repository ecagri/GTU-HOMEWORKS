`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qzwGsht3Yd0JwmP4eIFrErqndxsqgIcmEP5tJU3fCp2jlFNvv1mUrZaHHwyayv0n
K++4wkH6NxbwZT4jn610DweGqoL1Y4i/Z3HP3HDRIemCNYLBH36/xwU+Nycx0gLa
ATO8AbpI+WZv1ctzeXVyT9RG9tCmtenFndBgkUjIjkOvUxAFUFBI5yILGJx/8fOJ
FsirWKLw5/a3qUQ+kWdQO94j3D2YbP01wOTh3SoyPwRp80RO4I5Tl62wHq9RkHm0
bnX+6NPpHkp+EMt/yLsRRcV5kT0xzgjEURVlGrlJ5YxJomQ6tXp7BOoqryYqrcJs
enOmpX12K3knWuwNb8r/9wtJ8ewc/b/s6wQQCzvUk8+IOdeUSo308IMbjDH2/Lq4
FTOfJ0dDlBPFG3YQeMPhjsDZ1SjJjm7pmfiF/UQcUimt4cZOFMU9Nw3OwUSOURdy
C65+EABECNSVE380+XwjjJFiVTiuk8zNcRlu9xe3DF0QhO/Q2F+chH1qNmSepfO1
8wj08Vziw27k/MtkM0ul5KVFzpTaKvxQcwVMFy+ue96gUgH7ZMlLiMKCOBReedu4
5LWeTi6s/C8V/nh6JCKlCl6QmtpgFQ50UhHyaepAEnhfPWtbjwvC0JVm4/aPd+JW
4dmOkZwYs/E7Tx2B7bp17qyYJ9P3+J/YUZEnCWPNsCEWDEJsfa9L0I0qHMu1lwEK
jMElVJGQB3GC+K/ThiQjinvUrB7h7n1OZAx+6Vdb+bE=
`protect END_PROTECTED
