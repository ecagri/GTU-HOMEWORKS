`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a/EqVsxLKN+Vnn0nMvFGldBzkgZzfkCcui0e3SCRWc8jphHahtHosPuHhjmipNY1
snm2snh9AwRUoWmuRbv9mWUklK8RupwZ4gOnip7lajm763+Ia1gaxAWUc6enpH56
iMTs/SWH3gG4JHyfQUN5C0Ueuh4/MAGGZdNDHxX8LM5SPnBDq5ZQnl0Ya2GD0NZ7
RVamKe/5c/5PVWe63uOeHl4FQPeFBC1dkj25r85FGOBZw+3NM6mpBfmCWXTRxqDl
MBnVp4tFVOHRacN4Gs2suCABABX50tn0YhNm3MThXC10YP21YDIvnacU6OhPuzz+
dThVf4SEPxnvJEzyhXg9pGgQxN7fiUmbDi82fLXo0F6qGFeWV4L6zPqGwIKglatp
DcjV3YbY41kzeRFGuqepQIz68qsMiixPQdPeS+xbdoZFNIWK5QoUkE4E5MXc/lip
901MxD7q3zaJcadVJgS79esLamUEqRpBP4SbhcMwmO3SZE91YUTx7LVGkCkIL0qf
43rxyXZHoDMPlRptao2UIt7zBXhzHOfuZP964Qt6OuPY+VpDLKXwA7H7EBZ52A4L
M108pW51pa10Ouai1VQ9xSW8yPWcS+ibblg0tCurDJO8X0WkjdCSb/D6xxJsN7py
vkxukjrR3H2c34XEq9Uw8ROTa/Qp7CV35SQO7qgDvXObH9QMnBYf49QZaMU2z7iq
Bxw28FApUV9luHslxt4SSwbtP9+lO05IpeDZ0Xi30TAl8bsyvjudER+nW3YiG/B4
fVQ02NrzLaNBQ6JjmIIX00eBB7u/g1evReK+BEcpMkXnfg2OX5VyJ1V+GptLRTsS
J49iJX/EM2b1yunFZ9eGvvg+YGBBiSQqKZUJzVMgA1pUPI7bjebxsrUkrFVc5VWE
EmPQhmNN/V4PJohswm1+dFuWQDThDRy8DlAAfVIu9i3ROiTeWUs4Nr/uIp4DyPMf
s8zD6o6nTVbDZW6QJcsc0tzOvjChkW9sFu3qfx/DSD7WtAGkZ0SUXBZHVscU2JnL
DpFRIT3yR2XqN1E8iW3KsMd0sneCdTtl4PdgsObVs1j7hqyB8lYn1ceXtQoBTgkk
ao1o34GEMWlGs4/A6ZaaHsus6O+nc9dhFlKva0dffddT8Fvzt3bEpf1r+iMev8OV
HwHg5P3POtOa0X0eayuBu/QHJcrmRJAdqv2xwvqmdR/vPWKHw9H38AF/2/0J2n5m
nMVlzh9/NPYonb/lXAAnIABkPVeb27pbq/ex/fjMZrvmj9hIbA7QGlD5ZVyhApcI
/rwiERgLMj1AIqJ6d2oNHvIRqoCua4urDHwavNJhlbLT474na6681WYazxG0x/+q
ewWcaMDxiX1fn4WCqLsvhFxUcFbkoYDljS0l/liv0beziSmTvWDFb729+0aPiONX
PDpM7WwagyePvNRfg/OelcgrA5YJBYPNr70vxpP79LWNGY9+dELm7Vbnoteclt3W
ywVVxhHgSwWH+W0bjkfZ5WkNVuddr7srOlDvvVffLdVqUeZdygYnV5wxDUW6834G
bIOrgsdTGccu+C5xxMecCR72KsAZNizodLxvDfAnqpc1rc07xKt7rsy3XZLPLY5J
MTdq2bo7eNDrv68l5WpqtiG9tCLLvhqOB5DHElQWV7jWgtUmFIkNHef8U1b+WDHB
EX5awKKkjdNrT6X5q2MDa7+DyJCoGX5Or3oFLymntgZVBsxwELkr1nf+j7OE1+l7
GZDadOKKRkRB/GvhI24pqXHfqaRYfh8k4dq0UGQAdngusCE4HoGxOW74G7k3G5pk
cb5TRPvswCumLiRCnbCeseCJLKxEvkYtrZBxyFQPHWuKU2xUBH9FVD4pljW1kBSL
`protect END_PROTECTED
