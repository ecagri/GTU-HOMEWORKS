`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m+UPuDiTVf3bzPqst5HlnZvxQQ1uieJ+Yeuhc+qxZWxrkYYDBwud4UfdCH6Cck3r
Un5ViqOjtRqBPp1cP9CziwHb3WtDRRvcnF1vFPW2ALfRvNGIaaCqKzEMbm3gnijk
Gmw7U0yPgBraa3+siSqdvjhQmg47K/6xal3ggsM5Kn+s0mq0xdfXJx0EVoTQQxS2
8EHA6W3pTjY2CIVP6WALj9ZIcUmq32TX7d2k3MlNeUAG/gAs95BwVnqilb0F+g9l
JY4wJ0ywV/29HO20nRfl3ofLMKYwYyknZKocicy7/qsOzCPGL2GaKLHZ21BTLVNR
tBp0hE420A39Q3XgN+j4IH0MzDlYuJmFTuwGWHTJALkwphnjssUT/NbGSNgK2CIk
mEnDF4lTTdIaoiOUS2UHlzFyim32rexSFszM2VBrSM7iBQrf2KIySTM0ZBNTlwav
0ao8A2mjQcR8HsbTv3UoDjsmaJdgQSToqnM8Akeclo0JDJ27/T0yK8Nr+GG8vkGH
U0ZUw06G7cdjzx2FKEhvk2Clk7rbwHmCcIgjy3rPfgYSgaYpGlMWbDjfu7AzIu24
JUOyFY6UYv6+cYP7Rhv++rH+BhegqiCas0FzDF1EJnw1RIYj0Nc6LjTEr5KWBn7a
zmf6Eveu6g/LMLcAsOMOQzCBVPRLnIVrtsKhasRjirplruvGNPXZ9cbLIhDla7gR
lMFvluK3fqn0SnLNwhCs9ALx2JI4toUp1BA2VpG274ptb96YZSRNA1R/nUTj2aoz
MN8ucDkrL0CEqGPG+R/SVZuA27vHindVIuE1mjdP0J04T41IG9xNuzychPdvdcCz
tZztXzDHjWVIpGMbAYMzHwW8GWcyVADUbyQmBVugRkIJfLh4aNeSc4caH0KTwHex
T773sbV13RnRsOMhb/AV0v4vamtgE3IyQpOv49s8ucPOoVcYkLIA78XJs1No1udv
RDimYP4FRIORE+bhoZU7mwB2oNrugmayQHg4lhAJvo3GMG7tk4t9Jc2gPw5muuzH
DKzgMD6BtDLjf2AeZ1jONqbyShEBcSVgPhVOIN3T+pWA4OIK6Z+ubiJIi1GNnEfK
fnA8oKqxJNELoA2WQsWnJJDHxmB/Pcf0qwsDa59saRm5AzHLbqbXPZd5AlPqanp4
1yZ1mx6Mwn3YkKS3oUIUMY5BEUR645eiDYGN/03fi089PToh9J+2Rip05uiStu+i
yloK+1LfAwK8uA0src5PV0tM5EroJ8vqgPVfHqWE+POvYAU+cDsamZxCNlCQ/F0E
mm/qISIa7GIRU2jdjzpUtlMHwzFW7xcuo/8eQw9Los7/WoLJ4lXFpOY2Rr/tmObf
ynpxWsNKSxWQMOMMR4jfR5V+7zHnnK/kWk+jDkx4U6+ZBZfg+u0bCEx8Io4ZQOq9
3xpViJk8iUshP/meMAmO2I8tutjx5BkzoZfxEPDsc89c+JND2uoNghIBs340nEMv
+JKkgcrkIxEpkYc3Fs+E0tQfHfLTWlz3QNxbGdCVORB9hay5gk7SRoMFpNvgOcwd
JiMeD232/PZ4snBcRH0XnPp8eXDLzqo4xwbet+lZR/G7jTHCR+saFgF1KKq0yOAQ
Vk4UV2JPJOVA5UK/SQW5QgJxUC2kcrOjpALS8eYx6z4YthMLr/TKE5wmK2eo2IjM
csn6NrnbRbYfAVmzvIDDCErpNHDN7+GGRdLR20D7/TPK1n4KsgbyLA87djtU/lBb
MVdZyjC9kYONSPlyqLLnEO8vrFqHIe3bBBVNIqJCJvoS++VHaCrQ7W9vS1vKBZZK
tTtm/RC61M285mas9eTVfaOYrRI2WkaOGkSIhHwUH0EF0r31pwJBBM0NMio1oDs2
TULu9/aOjCYZcwItI0PDsRGIGsgdjZr3SY90p2hV/yCaRRFK6AO9woy6ehzS4Vd2
AfcZ3lgaZY+CrosG4dcY7HhJMuzs1+PoaNRdT8XXYZRad1TgoFOBAPLiKtrovBaJ
Fd3EKB4tEHtPFqyGDVxaYTPlCmMNYk2vLzFGhE+LgI3dqQVSsObuPHyYy+ysaAMt
bXjSQCYLefBRsiQDMhsoJTqPo5/yI3thMnMC+xS+pAEkW0fc1xY8AGlNJlY33soy
o0pBtN7rMnBfB9ZWbCDR63JbMs75DRcS5jG+NZwkW0Fe2VufNnrLQrER7n0KE4CO
sN9j6Qw8nvHC828Hjc6RsHoTVS9U2JVSR4BGCFWrTIPIRFCr8BqO2F5zVIvMHX3v
YA5FUy33VowqanUUh2y6BJO70XvyDPXWExBohb/YgJz5drUh2jWpAHlYVCIIMyxZ
ERIH2ZCGmMc/Zdi5XeMKehYqXOs+rZMXUAPXdB8odqiSvB8St0V2GH3tUbIHJdmZ
OMMJEfb9IjQg9f2TLb2W4K7CtJ6XmjuJ+20pkdaSWWLiFmQ2RC82QORzp+meOjgr
u+LeUduvhccLcu9pUuFg0a1P1nEX/Y96KRRVERzAoIzAXQmm6yQl6WqHjPKYIINr
RezgF+GNomLa8TWJWULAvaJgwgMtQ3y/kqSWlWOdFg86N0vwSQXPlaXACrcg1ovg
+0ALcDT/NzOXd4o+r+QzNTB1b2W2YuS1HjbQiV/h/r26wD9kQmR1lr/1Mx/imyK5
4PYZPbN7qRA/fAeZ5iM7XC1HdgaGzRmdyWLrDneT9XypAzCTKNRw2ilSuq+ZMjhP
9Jxj8X3EzS4Jw+1ij6me10bPZkBSX7atWWPRtzeHFPODklckeW8wSlpMZvXzJ3EY
29zeRQbgUap+kc72UTu2LpXXdJ/juAV9YDL/Nc6DbQUAWfK3167Kl5NW7nfXgytk
s9EXI7gfHub0oRP1KDSn5ytO3deBElQoXTYc+myOAhqszLhStPHKW0IaCGDWalUW
lNlLMdMLeK6U2//RR80CRvsSeERsf1QEEfC5RIRSacxIx5hMKkuB4UsdZjkOeV+F
QlQUO5DJhNp8pgYf7UhpxBB4UUXYkcsm1yQKxgS6xtvtdMHRfTrvsvMDgvcc7rpY
1gaiHORFq0e23LdeRuTPyJFcSRb8/HiHJw8pXf9RBrbEqEQQ0jZ1S9xrsjsoYSwf
R8ANV3/HFbFFSV6YMC68VQb0DFXc5DliYHWWvuvUGK4LFjmTsOkunqgXT7C+XduA
ynSH+A6ksf0Kcx65qgvmiSilLorJnJQhvmOjIDiqg/O9SStbmsmUr296cSdCweRC
05XvcxJiJ+8WdvnAHUGohg==
`protect END_PROTECTED
