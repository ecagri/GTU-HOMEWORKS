`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xOfxjjN2qGywgAekUFhFZGgKx5Q8p3FEgddTbOILC88dnflDmSit4jzufbKM2ZFG
pfikCZsQPxgw21dsW2i5Vm3Sw1qtDoNGNnm6PYQpTEXms6nRGevSOuMUunkjfV3p
X4VW07flmDUUY2OPg8tk2r9rAEetH0mp8gsgFR04kPzKpYQwIJwWAHc5Tby83/jD
7coKj5NUmGmItDFdzzDbaIugHIp9wwesqsFFetn5PX0C5wvbOjZU0tp/Kd2+Th7d
AZrA9psFaqckSHSwhlZbhprFlS+9/yTh9VWK0nx21p1FXFk96hMvBxiFKI9jaxZ9
Re/oBGe5S3GxpSj95tlXYon+passXelt7/KlzAdYwPea3v/GOUfzFh0G8PwTLdn/
4ixOVstNClf8j1dF+uCj92QTKodFgpn5PociUKAIXARf0LAv8iMY+FvgkYob037v
DKwtG9eN9mqPRBHmQh8+WLklMceNqB5kwuG9m39zl8KBX9bDJhXddy2RsbzXF5W9
n+RkryuYIAop0dwZCmjHx7QnagCBBLimuqhOcQKteQrzbFcB4IHi96gT1asfMthq
D7cEo7wYYo6xIRZk/v4BqhEHW0xOTaCCdPS3bXe9UbFbVyHA0QUs5uDkeIW1yIiw
G3xMq/iSbhDD/MFsfg0zrmrAvl+maoUEfVCxRaqeb7jn5dovMUD8HH1UyEacF7V5
IPhqxzbrr6v6s5okvn3+9nqLw07Hmnj/dInyt5qS0a4PbloAjjZI9qjD8ld9cKRL
oPj0aterafBKBTLSN8qUhGt0zsB7CcbF0WkBaxcD3YgRvHxMKuO+xnGVO1lNnPgv
jYeFnBVsgQxh3DkZsz0wbFIgI2j0Im3QYxhrRwA8OAHbg3KAfGhbcmeQAmYY99az
hEQ+kB8TZ3e8NfgTPNfttm+6YfEZIa2Pe+veh1qIjHOrqqERtLjup0SMwAFiXiat
CeRHcUpPTQAO4m1XNVz6H9n6IK5mzbMcZEQ74i5C87u+0Su2EaT69TUOVJXPknQq
Zo++0y3jS0NsW+OWsIyT51XJEqcJVUnEac1pnK+ibYsRsVMorYuvrOa5aXDexqJm
G5goxQSdwc6mMm7Rb9bxNPBofSqEj/bx8MW/eNnpAjhPV3w4PhQWI+sib4T5or/F
FTpkcL+QmRhLlCOlpl5zHgV6gdSzZHsxLVq6hrbwFSSgXotyUovPnu+6fj8H5dtY
A/CpzsSSWZHOGZ4+lZDKcXTfuWjBtRjtURqhpTS81arlvG02EoFCXDJZ61gSG7rm
gBDTXV6eiCOoejdNbSkRHvjOkxqJsPqwG5iX0vGBFN9gp4FSH6CMtmAoJ2WBIw+U
eWXsLgr9sbKZqyUGjgv2xORjamijTUDKsnzTQ37ShmALhznjnXWFMMIdnIrscgeg
6cKUNGNVKihQ9wgb359WsSsMfANxsSl5OznPa0MagkEI/F44mo48RWTbA4pw3Boy
pqqkaGfEVT8IsKIMz7fXGhQZ7wtuPIYqCw039zcbkIbSoKBZFHZZrf/ABwbPxGZB
mJkHHvkwswXU4eM4M+H2B9Ny/Bm2ZzUltvqmVyJU/pdY+1SDdj7BSILIHgfNQ2+5
+ZaRvxXQov44XM0S/rOZgHuupEQnW9lcs/h9Qggg3GEYfDkSR7S0/BCU9/7dSkNu
3+qKXz2EfhfBRoQ/o/fXi01a3WNupyfZvje2GMdpXLeTcqNBUPonPQYnHhiMm3hm
2/G6CC34d/FtZdOa1X5IgsCR8zX5/GbXPIENbFQZnhnINTogwOVcOODX6cuxdutz
rKSM1OBy7YyEEMrZXmYdveT/kM3hB0MRCEkuLY+YuJzvs+pG016VhfF3991Jkz3t
Fv+TQvDmkfIeYKXTaF+gzd4VTU26ri/5XTvtWMIkSt/cNTF+PxvzoXIOsrzTUY/1
xObwu19J+MqyfNdAINS43deMlpXXHlcW58wNOjRX8QMl53nymVkPYd7jeTZx7CxV
dbTrlwh5lz0vgLuAsoOeUs7ixmiFlG/jwOn/Wc15Mc/c522SfgDGP7Xmsu/59f41
JkoUHXSL53Y/5+b+1oK0tg==
`protect END_PROTECTED
