`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pQifV38h5hhoFGQVv58+d6woDzZTmarfxIBqb1XBcwMlVTNpv10i57qDEaQ1Flxl
0wG5TAQ21pDuUFiO2LAhF+gRtCfiOIMUzzwXgIqctipQpkEV3iJwhk6JxUm7Elnu
3crSTIyho96Tm1+jxADzwYx8pmvE82xjB+987lujsickPqX3bL6ZpqHHOmlJoX0c
6L4N86dAd92fe7xbCTI7OUdP8UaGWHZIqw08LYnA7g3q6/XqttysCPCs3odSK5z/
xACybGV34bw+gJuHIs8IAX4JKM9v3XAJ0L7NKCXRu0ti6yM4cpUxhzB13xNHTMJ7
d9F+eN0ZHGMYHrxG1SHSWGD7w9wZOJGPaVt2fXW70EEMlCZV7RsZ9u/bxE1p5IAi
sJ1r0dvU41xxDjjJUOFKhl5LJjPQdf7+Jvzfld853bfK4J9PSpIxvkG9+aV8BlcO
cjZzWxbzEpFnpO8YPB1+xSlaOACubzApYcY6dkl/E1t8AlfcQp7XjWI7DJwPW6IU
zcinwVTSjqlOlExFo2oS5gXYSquO0T5kNEU+CZPFhg6xGI/OUxwr9FW4DHo2v9nL
1A1cZb6oeCDR956snyasMy/rlGvKFMeR8wg1dz5K1mKWmhtDnnCxo1KXrB9dKdIQ
`protect END_PROTECTED
