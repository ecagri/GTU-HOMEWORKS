`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I/opgSYiGEoAvodC7b2XZVjUvoNBlJkqBR1Jm7N67NeK4L1PibpM2NKDIt1XOxL/
jgunrG1pPBBo2KHTT+dU2zQtDkZLdNwU25WX2BQZhVALR6ufXHQ49z9QYfBF2SBS
iQpSQX3OxSnufCm/s87WSzcJRNf8anEdJD4UxlvlKyHfwmqjmXSWu2da4WpmsMbl
6IKMI6zuAR2t861D67/Yp0ndbwsjdzTBMMknDktj/Qy23DTvhM4xpNiSiABsNwvx
Cyly6xUVyREKMwc/cUxfIJlcWSocH66MuqQ7mxkEdirN9XMcOUZinP7D2LCLPXb2
zOwYov6V4SnuHqxA3lMzu9UHXEcO1MpHA3yfO714/sGxsqQRvapMQ3xuUBLP+YXG
WfmDuXW/CZwtrYZ9bACj46/3eDhQ0lBWEZhgcMLn7HtXytAkovy/YpgiGKh7p+eG
T0O/XMT3vyQeFkuI6oEkpp/Ymd06w2djHVJAptEjWPZINSnqYbCt3JUuKq+6Agy0
XHJR6LcjuJLdj2bLmwS2cjCDoxp2sXy7QiEsWftPXon57E76KlOtaZraV74A1R7x
nG4PiFAYGMvIJ+pi93bLu/EAJfKOSc/iEunMpZmMb97f68W1+t0FbkvhpgJ0m5ao
Dc2xfXV6DoT7dneTviHPdDYepLaLqSuo2HuYHAoWdCACYw6BE+mt3lQuXXB4qT3y
mRewjL2PzZGumd4LKgczupBqSGTJCrF28Y9ZPVDwaM1utOtpvQqjETj7pOBkOLTk
9Ft6eG8x6MNmvsa7HIaOFDNP1v5eK1AJfKQ+KVWFF15Rms5Dgn3OcMhdzII1n99v
j0HYbI415O9L8c2/lhm3fi0YzRXf3FpBe0KHtiixZpN+d8WaAgQ53Xq2Swv/wnOE
M2PtjmRz3xhEBcQo9H6UcyQDaZ7Dx7u2Hs32CtV10HlVu7p+/UmHbbERPlCiHq5J
XgYkSz5Dq9VXcs4OPccnNEWOwaTrnLI+QxCYCbREn6y9r2nnqOJcvDYrwph9tqwM
jsaQzX6KIn0DMzcWdB5yvlo+AiH6QoSCw2UZDRrwSx85xask/KiZXMvJEy+eXQdE
6iBfwCa5kBtnbQxD8I4JdvzYxuH2laI5u96hH23qyhVt8nj/BX2/PJAquXJWV7H5
HBuSNRDpboc5hwHH9tOvgAyo4680j84bI3nk+4/YffoplwKj/cb9biVgol0ZtmaR
62lluxOFnZC6Axe9+ZqgngglTXEGqeNVc/vSPOu5VZT53T6L3KHeC2+OovheX7Ox
l6nDi9RIAoK7WnpLFjbA1EpG9kUeDz7TfyWCnTjFyUve7fIoxCbxbILMwimLWy4p
HizrO5J1FsclttqgSWgjbCDXnpjHzbFwk2J4cJEVjZJwbw5FdFSbsJwkMntk6Dxo
0X57MbEv7OVoJYO/jZNPJ/UJqWDxaKGWoFl9g6w7VtJs2EUDmjaia7BRo/Ev0dOD
VeL8lHxks/F3++C1GAc/IJcqbvVQGBqLRxWXFtUxSi5cjy6q8oAZ9qYVOzrUTcGE
h4Vs211D+gfDA08U78lT7argf0b/Ga3p0/Gw2ChPtGUYmzCMU4LfGAAQWrZJ8VT5
yCvcYTCX9V054bb4MuzEA+kQaSwrNat9tpahNZiDV4OkS+sN2cvRnRSXvx/mf6h/
iCeskdaD+QwMsmiDJZeju/I6OZJDTpS4+gE5J1xpKNv8Wph7Z28M9s+i6dUyOxHv
wy4AJ7Klmfy7kTu7F+Orz3CpIc23ueahjLc7PvhwMelrN7tMJlxkADrft2urtv0b
Bv/za0MAcOZ7aFCljUNHD0DNRTp1U3XGTA8EgZ/SrctD3YVYXUkplYVy9VjgyrEa
A2QrAkSoRniSREhg24OGQA==
`protect END_PROTECTED
