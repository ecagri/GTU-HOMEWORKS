`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g9FRFJr7B0HB2JWSUZt9tuLGm5ddFNDzYPVmkcxZpHcBpIlPgd3sA0FE0nlIbADC
AwOdRYVtDDEV8l7IFLwMGbRxi1NEFlRrVRNvu++6ySdR3Vjas85yGinMaoQeLhId
uDVU8S1GTgKjtVoDB7WBqvQNf9Mk0akcgts5YYmmKnFQPQ+6tdUVfXnS+7NlxWzs
GtRtpX67qx83RVf5GmlwJP/A81IjpJfxfWi/wLG4tiAFwpd8V2+R6zwrxiCCW2VZ
DmrIImg+Lzq8N6jBmkNtqrgO+er4OlERu+l2b7n1mlM2pDh609zvQ2NBiqbzgomM
91PVW4H5eXdI9vKXEd7+p7Q/swJ33zhPMHYThsTR7ZGxtNbfv3hyp1a2kWKrA9ms
b6nZ/gfzlw07q2Yic70lW+iASzc/RD1yjW8R6MWlRqJhgrTeLIvUUdgdbTZ78QLD
45Ww12n6CvZu1IdK5NcHUg==
`protect END_PROTECTED
