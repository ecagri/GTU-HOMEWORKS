`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kwACzp31B8L7uF0ckCUwJ4OPG4wtkzX4Yo3+3U62NenFa3wUaTEt2dYhOk0JzpSo
gK7USoBoXPfHEfaOwPdcFklqi3HMSeQXDrZrE1ncsvi8m4H6ChvWT4+wr38dXUw+
TqIEDokMc0bT/9ffsGYZNNJsSYT2R37uYB5E78LVdbnJMrR5cteSFM5OaZZJqLmJ
SwK7qz6efygsP1YxNF0oeM9bd6hw+DUD9+OVMYodNLiqyulYFBtcDwutsxEB5z/C
V8AagfDPCelg8tCsgqLXkXmJpIsr+SfwweBhtYE4tLVCbqFtnuzRYIz9apFsDzyX
y3Np/bS8FCbEYIuWnN1v1tMKozwbaWZdiDb1gVwSHLbUWbnRY6eoaa8Raub8sks8
R24miewsBx3hmXXb2Ah35q6CPnMgrhA1+KVjceWAsTsOLr8kFQaa1be3MyyJoA9e
zbA3qXaa409sQe+dNjI6Bu5pboW/xhXHcXykWnZvtcOxFvBG741e+QNcDWmRI0XD
juPcJvi5lLucoLwTk5WFvZBBfkyz4189ClVPgpkAizynjGFCJihHTEc1L82iuJ+s
G3YwOgnm02XyxaH+ULHZ/P5H70Ef7PrB0s+AIibC8gM=
`protect END_PROTECTED
