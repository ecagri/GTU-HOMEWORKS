`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fHJTCt7YflQTaMxrTEXpNKaG0Ay4173E2K3XXQvacd8jh2XVH01lYe0BOMNmYb25
pEYQflSNn1PqpYJDdS66l3ua9xjjvV7kCGc8FyRMjtzwZstoaZnRd7XQoOKzWnpV
B0JQM7Pc4QdsNT3P9EkHt6+lw5Xpru8x88/4eDEnJf/M/OPtuX40hz6Um0ZqmlVG
T5hyOF+WbXbz0/v576i9mtfJkD/+KGTdHc3SO+OGVLSAk+aRhSWfrNh0dRRkaXiz
zCQM8H3QJJZV+gXbyveXpgh407hsvtXzm/OBdR+AN5z7S6BjIWLHumVeZa5WO/sw
FqGBju7+L9eChaBZfFbwBGpBuK6h4h+mFJrkTWdz0zB428NhxNAgFpKO+zy+/3tb
`protect END_PROTECTED
