`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IZIVJws0GQhTe0r/ViRIA4Zv2OAnwiMVIdi0SoCetMD4//Vf8kgMH7GT3Y3NTevM
CNyd56WjkCaOzNr0QTdxxlOBfaPwtLaVAoP74QauW/Aq2YnjzbNT1nu6O2sBTiK/
Hvd9YOHQiYwrs3EQO3gcVwXWGT15gNYny1A52PaGEZkfYx8tPeHJMnRkpqT8ePCv
6MlOhKWRIzNXu4+vjTN7MU4CRarW/uTxbC6F+RJY/RPxQtc9IndYyLM2cXIXrlYw
Y4NYnhlGgUOH8hf+F0bQJxa3rzStUCSYkrwes0L6b6wczgm8svpvdI/YPgA0uiNF
6nCLKqFY6j5WEPGHIKRiHd/yydu+ElRZBSBVFhuFkZk16cO8T6tcdfUke2XsArtQ
x5GzPNHt6+qhBeh1FnsUzCqomiAkku1w/9AJSaseuouQPAhKVU29oq3Wx7w2Nue3
+JzqS0fcfF2rnpy2QjPGnh5zHOWcz2O7TdtTZ9sbZYHzLc/lEzc54du8SjqdXDBT
+mifST5/WFoeAJnTD1vXDXl+wrP6CQWwPOEGcGNabvOxccPsXdBZPA1wQ2jnqW6n
rV/llPt/v0E4wTdFV3hh57QtuhVlkG5s+Sf/6Yh6mBnb/T469c9CECnwipSLGk2b
yBcIOqMmAhSeWKPDXSo1LCYwcAyVWBo1gzxUc0JdH2Z/2JH1ci2Pb8Hj1MVqsKeY
rQTMvnZGKF0zhqy7ZbUUU8to8ZH+NCfUTM3TMLT6++HbIKSmKr7ji6Laq/Za46jG
ItoOzxx5hD3vem8ph9KhwPoz4UWyp78i8qShlJKouFnaSUwtmeX2PM/QRcS/WDFv
1J2h59rYWPMRryH8v6NrJaTetCBCxE642J7QR6OA5IwCny6dhw3xUEEQqxlyLYr9
JCv2TS7kAj4byYfbTO4PAOiCCiGRctk2qqBzCUMXtOONtiIcptYb3gmtJuS5Pvxt
CX2Zy7/aPx5vjMLfKVsELHxUn/Mi0GvZ+vwSxYJL+MJnpC8AyBtSA4QTE6Otu3D9
KwT1dUJzhX+0k2v66ZERADnV8AI+36iblaUEXji7fxrDN7Gi64bYhzeBdcAuTLuu
dkjdju8Uck0Mdc/1KFYCsi7xfe0n8u2nf5IBl3I2yi6kqbBZ6N3Q77HHxHgjPeio
TZ3V+iLa/C0ZEOEl8wK7/tR4tAnw1cnzk5IdUa1/FMZwL2oYONEkg7xcpGBN+JDC
thADSnrY/5aK3JxsZLWgR5z4PWTe1GytyW71no1+RgS3t/f4edY7bxlHEH2LLNbq
W1jgJPDkI2oWa0IPQ6p8wrKCfNeLQLned4riAO24UEVe6lbwbWpz7gySo2WNrxEQ
Ky1IXzjqu6pcAiGMhuKRrbsGnljTmU/HL5WmynOXi68+JaJyG36F1qIPlVbcYrl6
gRYltfwFMk5Xs/JDTO7aHwkkv3sJeX1heppDWpCCCR6pmQ6mIngXfZ8MBH1447LA
lBklLwjtba/J6qlpkl+KqTfBZU9sEOzyd4qUhVi2P1Paqmrzv8hlOOUc1k+wUN3b
ivu0TDWtAyF8Mk8JkcstF3wzae1o47Y+8JQ1E6Bgixk6dNNgog14vY3BWwUXlxLv
ixGSBzEoGoj1+ua3K6dYQG0oFerXxVmD8xLufsjdGVTkRmo7r1RQuAtSdEEO5b0w
AVlv7QtwpYDxMh8Oim46OgvCvALjwv8UEpIS8gzA8paspqBLMm45mN3fs0Scrym9
XtTuAnJitkF9htLXBRPx6+SR9cPAgswyqNZv3zWkY14+EZeYei/1hEMlWyriIw8/
lOVnVPnvua2XlrOz/6MO0X0VYCngy8vYECQ4uom3w+dshLjORyAFXOpZm1pxlNWv
+ZLmapkDNysTuyjH6b4gNIvASsEkRZGLlfNQ1PCyMtJWtqZgAnG6hLso90cbkQTM
b9oKCeXLedEp2c2vSx7dZTGWGeVPEctvia0yQLqcb2SJLPnAaogULMMvrw9amkC6
/dMyApO1U5/cJeSiqWGFDw2XUQokEDIG7Q3/Gj6W2ljyVORsqJCYyYiYQjFGVlks
CkXQKi+N5CQOsBNuWM190ufTq+CwS4SlasQ0zfqdJ6UoGMiRuNTVxh5PFdPmXWSb
NzqIa7+Ga0qrclcGELfN/wg4ijNNx/plilnZfVtVGJUwW0t+M0uNKXo+VgIVSrXh
wOdqqSFBxcbOn5F2RUWOAbbgw8z3mNbrEut5Zqdm+a2kOvLz1/wF6IDUR2OEz+Kf
nHGPlRa9Vw3oCLBQNL7c6ydJGnyxVaf8FWMZF0Of0MYP0NflFdCmKpx86A32g5p9
XdOi4g6G55n99onAn4pusyC5E/mwiyqedSXn7YDNzpvzXsJFRAzjtZcQ+GJj8COH
R0FzvSo5LoGPI29XXZoknG2rqJccRDO8gdUBhyor512li9d3ySOvj89LQRZbHPA4
MNp4TJxCPFsAjm53B4X6yTE1tWVO+XgYi8BBtmaxgj4sMyVnpOznmGCIGXsZ6FAH
KJ0uav0JMNmoj2hto9NXr+vQwjGTY1WCb+1J3dPiOxoQY3ZOg3tLCVL+xqJsKUq3
2V5UmEM9pxtgPEGUZfWYzsgBzX6PSPINEzH+qD2agPFYyv5l8hVN9OFKUdi6SD9C
x8PMwAeIFXh3xLeMLwqhx1xQyHVrlj4iMrmKfafYxnuURB5iM4SST9ACxoIRT2MQ
p8YtmozGfEebCmsQ0VqnCic12axicnoJ/XIKscNgZwq7WcfLTF0kseOY40MQ8FS6
NDSfIzXden8jprexLd6cko5j999cJFLQfKVR6deftpvsXA/qjxQiyOg3hj6xiwD8
+HJdv42AugYsCKjxjbb1CFSY3zAg5kfQnYU16YDcu06CfBa7sbIKrgU+ViYlLu07
GlKr7UO2kGGg8suYV4tJk9R/NWS+aJ+FGFulSkeQug1kFufO/CEdGTwjuIvC4SUi
NmKOtUp6IrwLG62RY8DlNph2yQ70mvwtQClhnv+hvktuBlSxc0lXYrbWCsayTIQD
yEFTHS2ndJW1HtkObO6HGaQvREmAUrEEIY5rU7F65CvuWWEAIDmM9TeJiBzq89iy
eMWh9bWwzVQwBoPfTGrlKmgZKIvsa1XqtD4hJgfSjULascoMWIW40SpoVNxTwCS2
ItD8aYPwPq/P4u4QYGI5ME1qnm8vvHALgtfmA/x/f/Zz2j58v14+EtiPor1CcFBS
I7x0B5v+wnhSKTXfx49TfeB7N0zaoee3c2XltltUUTzSkJHMDa/cLgBwWU9bOfZS
KIDxPyzbVf+FPaMuPGnx8LF9JxsrOYw86feDY8tSgf2yKJmt1pfzMPSJTDRsaUQw
FaCU0OQVYd9is2hzbx0p7EvX0CpCJYUzz9F+jb6JYji8Ne3eV8IuJtR17ajEbDrL
sQybnOI3vsjuSLHzCrcPn/7WSWvC7B1ZQ9ls7+X4HUCkct4JohA0MM8PSuUIT7GC
4cX+5mqFc2nvB5ngLISd9QpBBXzB3eIyZ4sdfGC+xRQ7vhhs35n66Zd3tGr4nHV0
shf/tt4Z1LVPbI5wMmP3zH61e1S+XtlGSluqhnoF+E1uKzZImoUzHwLfJwpxez98
dW5TPkWvNMJjiQo2z7Vzxn1yAKJIIDea0bOkbdPJOYxbWU6gf4yC6rsrpkQ5d4VD
olJ5OH3fDkklhUNLCdzTbT99+VUeH8yDdIYWhVvkGEnlH6p+un9za6+3KeVx46Ic
GF52W9du9j/Rq8C2QcrwpwUlV1iHg1yCGAOBAqKw8v30Yg1CqaITNsmWy1IZsV0s
8u6LfUcGWIW2XwZwQ3TzDbHWNOigCqlLQRtl7klvUPn3MjmQ9swetUcyFd4iqgNd
9OFLJd9Pd2WP+ib3LNurNL3QUScHOuZk1uDI4tMn2M1bEB+UTWF+VI/0PSmNw8pj
2yBqMt1nCaMFiEKeeHSTty4XS00xGqD1PgU0f6RzKxOxn1gShapmkVrjEZhmcoRY
S++gUN/XbBdT5XKJX/rLjcEFjiqSKooOgQsmwxbocWa3e6koJF0nhXAPUYTO5QqH
FIQ4AeGbLOqA7EQO35zddSLzn+QRkjQI6gp5Q0jv3wJAfwx2BZBbli0pubDjr1Dv
ixl3p7EaSyPLePsyKSFr03aBMp1m1pINVv8j8Y0bYHlbe3EtB7LKySR+os9vPX7a
e4anGbDaLSfSv5r0eN8EqLW8CENb2WhsqYaO5nAMO9V1xDhPhfC0jII9worh4exd
3QJy21siiGL0fpYGeSDkhBnFWokkCILJjKRqJAO5aX8tuSfFM6cISCgwOJ1lkS4p
+3VghW0Q7AYhmPOM19j6bGao5wBToWqmwahrhyMzh6UurHVVeZVPuws0lZOe6rv5
Az9u3ek3IEv0IjhIscDNW27yXUYD9ZN3gL8FvoxvBeXCDf4DmrY6SoEpC+ZWHMYG
2OboemtM73DkTW4Z3MNFPYjSWNMQUk6vpS5bxTsaN/SDJ10zHxaKVyORLKZQIl/B
d3wgQ//0hvLXppgcLQ6jB0XuGS5c1SVRgGLkxMwu8oMILyYFubC/YmPJSAKrH/+X
z3k4eAsfGPEujTyrxC91tqX1afIMhTwKzigo+jrqcERhGDxIAvcbMTIEZ8qtyQ53
FUZFKMPv28hPWu1RacBgwDIhi/Uf8nSdH+lYRfYp768nBL4nsCqw7rWs1RAolRBM
DB1jeR7jAbLPbi0yw3cXNXSe07OGID7VO7IEGasitn9T2djpWyITXG//pZhVpm5h
4OKV4R8+DOuQCm9Wrpj3/bAb19/HL1qMeug9QQ9irO9JUe8f1hk4NLHB9tKeTOK0
BQlU1sxbZVpbhiw9ufameqby+MqjhmRsdd6NYM98c0VfbtclcpfR2h79HOpbrK2Q
aZfVVxO72X5ELnv8nDh9slVzyBhZpCCLMy5cY9+s6b3JCr1c/ttPW0GdXiffqhGv
QyVPyLuADdA4UyEsiOov/pyc8W+u5Ub+vo2OJNtEzJ817uCK/qlbDqFIiJtzrSmJ
lEH2OPPVdCPITk7p34te/cwQzWqGiwwoGht/IRC0TriaYcwCPYheD+b2fDrJetWJ
4DK8ROfQTnwRM3mvxGyYAyxee20EF/umqLXACmnQX3XSOXU8b5I561WiUgCASaUW
yu/lZG0BZ78SsHpDa54w3cHSYVxr2OgDt8EDhUNPNu73SyTQqcLtnKBg13yKIyd4
NqK5HebltUMe1enZqVnqDIV/iANWCfQH9zmw1pV2QOx4vtfzm9Djn0w6A75qPo5b
MdlMb0k+arnIehEhiWjqyKqOK2oKzVftNTY1AWhOd0y03P5c5DK0r62LrjVH6QSY
uQGu0PZZ2BNS2gDKRqId5TZWU6jaokpjUXADprNtnZEAMsHRciXOkgQJRredFWZ1
7txeh7Jd4b+cMikka/yuAAG7Xo6bAIA6Sb8Q7Co4awlePei/jM27ccekssqJ6o6S
zuiR5Yw3NI0wrkf/w8fXRrhl0PM5MAEiiwNSH1ak25aToF24zX8jdukGt1HIA5IO
PWsNX1uZJuHcM4oPr7Jd+fRbA7CwnXMkHK9BeiR/P/susGTYZ9zAfO6uJAhof28s
ZzfJe0TgZ9KxT/3optxCzXQ4AzJO6Wn58e+9z5uCpr1At1wzHc2ayfAwkQWnZdSS
yZMyuJ553R4Ix87iTfLn2Y7I/BFZqwiWphgixmtzF2nFcU9ZxW2usmz1vy+nGV9S
j30ciez9Y/QhB/5Q77rg6cJ5s15i0Yj1/W0SsJRVKVjEZRYKVwOckHYVTyGGkEeG
pE2j7RM8onOAMhY5GPwX+j+BvetOPlbG5+KqoRqJQAI4maUEo5Jw/0yobMCG7g9H
4U3XmxukGtBrDyKxLTE95LL5z9FEM1Ui99RLq2n6+0SyZkW+zb4BeIn+UxRdx7k3
obBV+pCE8Doh015Fc89w25Lo9BTMbJu0QIzfbvWHQeqqbijxsUAlV3fHn3wGiCd6
ltjnGHXCDXszBLVhJCv3wc4YG/BHlymU+B6zu7wU6nzu1CebF1tB2tbo4ZlLtE9Z
1WgxdrsWWLB/7pQYNFZsCUl/aeUNVx/+pt63Vklnc0U/GhO+Y3nTo0iKIlNiCqlG
WJkmNj5GaSXqNLuPxsfKY3XJhber2tnp6SiTaXXFZguBoC9d2zaJF/ItU0df7IHE
T3ukOKZhVzmGJj6DwiSB3HgTR1vWSR4/DHDUu+HxeK4rt4cW/Wo2COVA0dWeBbiG
6lmYzBCVPwgYsDWyGp1xY1sxqUj/tTK03+QZSCjsZQe+KCzFEONUY8zCOqFkY4nq
4RmaYF7PjuF/yyCy7vBBgn0MuSt6pIUNeU/LTbgTNdhpndXnJPNTa4sBESpujTPo
EdsUL4SSByse8/YM96QtoMdEZSrXACTFyyFHQxMyfXz+2/XFuqbsTb3qfy1RASIF
XdDuJk47ETRzuQaRiRMetgq/eGyQyYm+57OmDgcSKXeOhh32nY108rLszVyTtt5J
kecBAs4JedVSvPgY5O9qHjg3B88U38a0ejA9KYl1HpMMcCF5lpW1C/6ZsS3yRtAk
`protect END_PROTECTED
