`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ni2ZlRVL3YPTA4obBe2TD0A6QWMxvwkM//9wGPOGxe1T9DhqlmwRf5QVpZmEjRlX
lhVrVrY/PckJl1HHgFyE49b8gzVHO1YE6zxEqHvO60HJSgyG1I/axqJ0C6FQ2pz4
jdPVc9J1KJL6SMC2nI+zYuiezbRsbeJB8JGzi2bCvQSXHQoqx/riACM2XEBRIFds
iOzPTvkJz6Yk25bItrxMsPkHgf+fSVnSwXoix8M/Cli3TER1+6dwTawySsnaDN5Y
4RR0VfgCyXlQj/h5TwToD1/qORuTZvvNVMtDQY+MtzblyJeuFk/pB7AGc/scpWpm
2MKt3XxelD6cJm2F8d9Rb22EhR56nX6/K2B97tshQiMFq+nlIJGkGq0VpcoAXatP
iP+VwxxsUrTctJsFqfWd11MzM3LsULtiPx5vyHWHBd2OK3KD2L1l9F3mfHhC/Cge
E3vuwOn/gvRyxxGHRGwSnwcheFtr4XLTZiMzQkV3p3aNCjX3xVPpt2mwz+/qoy+B
9OEKieF7K5w/g4voyiOmB/fh+TYkI3ciFuenT9CskTt1tz7TbkWeiK+g+pn94H1t
5nrv1VUEpCHxxsaUOjy5G8IdXWTsTCIQKFC577hVE9S/+DhZGDK29NBJK5Z1HDDo
xT3KVjGi0Rp6o/ZvFS4s0cNgNgUCGRdODhuBXXvYzgjVxgX+jpmLYOwxysddGhqR
RImcRPUfPnpWc4GFtK9fX3hKVwQclJmoKiqWamWpW3noOXja2ktn+BwebSLCpMI6
vA+/zMVRQjsuhwFYVh3q+h4VCz6bUh8Xqomltb9bYJ9xGn0NwA7Qrw4rf3LAzEc3
w6NtCpsAHip/lZV9IXsSuuLe4tgSOInuPDuisTgeHpCwqipBO0UbYXbPWDeF8EKz
8I+jJFVIdjddAJ6k/9ZNQqqMCb5ypuQhy5Tq8XP+AOQBh2RlKZqesQxYnDJeHblk
t8skgcvkcigkJ/8RXVY1MCSRrbKzRrdBwJ3lrwX/sXYwrIJgJ8B87wVGc1cf3M/r
ztMkZP+dfYyA9W1x5FZnfd5nYIM48vayK2C+pNhxkdlc3DWNqGCKoyWbb/1YyJKl
D+6j8jV/pSrsKV8YQBorOJ/4UOMrEGBxu/7vKEuGlKmA2QCjyCN7bWNA8te1x5H6
FJUYtcZvZRksK0JV9o7yKg+bEZkxAecIbpCFRzcMD0YyQb2dynro/Cf1ZUORQhx1
DdAJVQ8ifSDPuG2rdf4uk6TggjkMs8ErFuw/klqCK6v3KC+JN1WDbYopUCL9B1n2
u0b9Am27V4VB9u4APapQ6da1Z3aYlK/bjwdkq6wDX9r8W3u9PwgC6H+7d33bfgnv
zKUwtfxGYGEkZBBcaJOREOFVzse28gAH4wp2203SZedSHbWQ5HVFL4eLOrzvMZDX
9QZ5ZKxLajg7NhWl4Jfl4G8bc1zo/ZoXmPeJn6QDg1C+KqlPQ4i3flYHuXySQwwN
nQTu0Y31VJMwnWStI+oFE9BmsC/cWkCElvAQvc+dRXKVz1eS+ytqZL4odxhkMxH+
jg4152+l9ZwNhS+huOl9y1YJXg9HYy1epxD8Xk8Hbcv7LiQLodcw00Wp6RunLQnk
Ka9Bb4ac2vRFxKrF8D/nz6vx+WskXCxENEM6+X7QMh6wvoRPqqC70zHaKFtPrYhO
jqAScn3v3TjzW/UIs/j0VhtC6i07RTm2M6yXlw3ugMipdOplDOHwqOykzLU91uEY
j8r9+gXj2J6OM/VaC1HEDIx8xGwi2x1vqAsM9nLhmZENzeb5UGkv1Q7Knbus09di
XVFb6F0AIImgsTxGPtESiQAmXAvYuI4a05DgjxWUIv9Ki/UuZukPVX1Sz6zeZjL8
nwSHL1wG8ANKyjIKSnfHo3+aVpIYB3PzjqoIufuUMN4b50DfoXUNdm7ioY0OeunI
s6+LnKZ92/j3AQii9IWUQ31K/oE5GdxDVapD1WzwzjyQTlz8vBfR4+2Fi/EktubR
zpy1Ruhg/pP9KvdMggO0jCHMr/c0WTJ1iyQFNe+Xt85KkLa+1Tib5Awwnn/65H3S
ZMUkxc1CuPMqGYpn/0F6nt0kQuHu0fUjusmD7z6UtkQ2trekYbgRWmzA6YTm8f+O
5pKr6sujgkYkkLXgj1mFFXCNwPuaCIydf3fkVLaKRh4wXXwzuzZ9vPqYKNrvl0Jg
SCmdLCj5SNlOIllp9mhQiAVIXxtcEy7zzLbBQN8f9MTo8mTQpu+kQRBphE5ikHWq
hQFX6OFXWJmvvpmLu2y3sx8V+ZLrMjUcgw564LRiZXegY9f/mYazm6uLJ//HTMgU
TwVBjgrIpyb0Yx/2+1e20B3nc4ZiD7Xu30NDS6BfjkV4VJWA2Dl05JEriSXfaQbQ
RA759kM5ynub6tyAc6NWwT8PAHQredmpZF18IgiesrIDbSvE1j1zdlgU8O2NLwtE
I1i9YsmqAuGfID8z39ZURvHeEyStmNtEwobfrTwbiijmGfgzKzpOhtGzYOeF+0gQ
mHwDqgV0ubC3/k2sfj3BXQ==
`protect END_PROTECTED
