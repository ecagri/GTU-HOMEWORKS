`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0JLLUDnHK8WuRZt3rzAJEaubdN9w2w9A/T7Zrr2wGvF/YVr2KBLqbRhIcFSRzkpk
F9SEbujLRCJMwDiw1w3hqxoml4Ul644rAooZTN9ipADaV+6wa0ETgyZl+B4LAGTC
ml/aCEIX0wUwN7dnYx7MmEApKAXUNIKm9gy7jgzjVSgxJt95XVPP5s52ky6BdWZk
PSNBnrR1PftauklowSCuXRQEvBspRmGETNTBlhEpwyWZmVnX0sQOhSY0qVDPOOUf
l8JfCyrIk4yjfvoLSUHbQzv+Gj4bKdp9/fOJRocztdgohMpPVMeohAifPn58H3+S
TAl9PJHzhW6T5wJIlfNUDZLEbX4OOJ3mnoJkC/jADK9qX2xDuP943JV8vWOrtkqw
sLSSi+c4tb5rfXZ/Xb2y/l6nu7ZzuGrMu6jALSCBqE9hNuaTuDucvnBGYlCWKarV
a7EmDxj9bLBK406avFTXT9pIqgQYmg1Kb3Vxd6IfaDUMEJySONEn/BnCMvYo/A1w
MaXh/o5lCuXEh62m9oYxx0R3MDcUjsW54eZcifPVvRBSPlmwUttJzSVnyhlJXl/N
Gt5zjHxI+kcfwEnDlFTEQBNrJX/nViICVc7TMVlkkp2MzUkrQWL2h2F4VrMG8G7O
UppUlDkRN6qoz9SY+PW56xyTFWNOn5fY0gioJG+rwKIgKQb+4li4U9A9f+OUWw7h
+SLFvhqKdAoLCsAfq+apTtdp7PMjZsPOXvWtbddmIgEIY4Su04V1kWhxZSN/5PGA
3U4Hix9YEA9764E+erixntqh4FTzaNXdv1udIQpQS7eZiSWJiOH5TolJ8a3o9KbZ
aBMB9gXhDLNbMsOPY69xnCJMV6p5gsTBMueHarhNDk8kVOdEXhCqly9hI556VPUK
14ITJSMfy4YZuD240f9nnsNdyw8lY2ll7XwCfN5OQ9R2Us5/j7XkaFZuMhxDCXNy
ahGGdDYoQHObPhJedxw7vbAh9j4huuRKY66q2sIBXY/yQM4LBs6++4W82kaWaTbj
m3L/wY2NBykI2ul8zrXQhiIw62WxUTeOyt1iz+1eY46JLS1NE4/HkHbZK7AbM59/
EM7D/q8fNc+tLbK61nz28OuNYNZKIsHhOn+Q0vBm8ogDe84P+43RN7jSeXKYrF6S
hZmIpTT4Mdyl80caLLEt5MLKYz46sA9amN6l3Py+lqQaDUNWTM4fVMd1dQ41trw8
juwsDl8Ok9VXDUDOBT+hBZw6lrbOCR4v6fZ/zsk4iwnmBInIvzj6CCWtRKAO9xWT
V++bFaOn+N2dNCZAQYRLTzdSVAOQMzHU2gQGg1Bf8NnfoGf3VFSxnfh8s48Qv99Y
G5F6ht+XEZjEp8plDkMg2qzCDaUqwZwc6miPF3TWg37dgqq0LykbobKpnjMULDS2
VtUieRNs81eJiclEyOsR1CwmjhyAvaDgaHfjIWWCAAcTjCrqfiiudsSV2BBfbGTb
gZ6Yl3UJ4b9/RwCWjB+O8t7qe+UPaIY+Q7oqHHmThP2IsB5QTWoi0Qkvpj8ETYoo
9PzC3Jcrfwud1coQ/5xGpvS0IJ2vyUYBQS259+FUQHIZMCCj9IQY7qtCO1xyAj+K
jLCFqwcz2JuYXbA6qK5aawwDMQ+8F1oF51fW4MP4iKuwta1oNzywzAv0H30ffaFn
rJhQB6/sSAcuLhe70LnXI1XwVT3RPtHdKvWab55IbSKBdO5d8reeF8XBXR9li4sT
spioWcXGuc3tuLEewNHBZTPdA0reAzPEUPILYXGnKg1JASXUdbmjq2N4Tv+pIQso
VxC3Uzg2OJCKddB1ggK7cj6CqAem4IN8JRQCwzyurJLus8aC948/WtBgZXQ5he0Q
Fdj3DA9goftNOvBJP2N8EyYOmRDXEX0NJJOQTKdR8Xo0G2MvJMWxwcjPD0omd8d7
JgPiswKF+8+ln1bzrn3Nj5Ps9VGRX75ryIgdrGLCgueAvN/4iWnidT5+PpUFcByr
xLeVtsuLY+XNqpS6kQ/fcv1qSJY8Rg7uCmMDmHJ+oRGbjvVASaYIsG8sGLm23ayC
Mnp3KNKvv70DFq4umFsYYAP7X+dJGm8LdSVUa4s55rIpZxxEHREWATmVf6J+Xx1k
M2XUGHZmiKvoysTFn/gxi1TWwt8UnXfQr1fB00uJXFP2CFs115e0UMhD3Ul3yaDS
3yy7qIHcg6jLWmqKMSZka4AwKj3QASWn9yonbumigNxDEBAmh/F2M2rHTs0PIrVG
epHuPas871A51jorrxUpMn4JyvNkxQxCcTsNeFH0CBtGGVVmXkWS+iykHJ+YLz3M
kFrBBqTY88I5XnJR4npj4W24oZtBumvRnTwg3tjXldo4L74DGwuz8YwEU42Z+RVm
6oPTi9JznSXDg7PFR+4uz7XwAq7HRvMRR5tcuAVPbrQhUMkBUpC69Ym+jxnlfNzG
/gdpz2tynzMoF/rIOu2AfCz8ACwFYe7gTVkS1hDyBOU=
`protect END_PROTECTED
