`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mxg7+ZwU1G561UEldHF+YNtI8C/PER/AWSzeB7WLylvJFIWogsS1LVb590JXwH6X
2rdw6UnkLOCrM4ogzbz9WUfSPkHjAOtXr6MzPDlLSuMW0YNWs23TCza5Vn3wT4bN
70NBN8jO5/xndrCgn4QBJHSx64LU7CCSf7we3TBqWFEXxI6OvWwBx4f+xIc56XRA
x6Ilzyd9C6+iF1zrx2dpxt5SzFNsVzvoJMEzWB7jv9JLYEYbZEVBXARXBpmHUpBf
5yiMFuse1Olq6yrfEYoOEVCmpjsg20100Kc1uLgaGhqQXpPCMlaTUy68vCOdH1bv
lFnK4eAe4oDYx1BuuuI6RrzosLptL/h0y/amdmGf47/MZ+PFoK6UItA+Ky18WwjW
02xkwslBQ/xHtLpwu1rXd5NWlupKxaB3+ckJjVKfY/QDiRq3ryof4yfsyAvW9VWO
cIKBeoDlOn1eiA1uSWCOT8o3zMIhTmhtSFtubgMa23sCTw+/hHJ9EDnTSTK9SPgT
H14/OrrQO9KaNagf1TSlMuhZRESj78OlyFz9IZwxQR/SAd880kLhRERVfcgZd04+
cQ826TSrMVD5dCc7dOXV3lvGAubra+YmZpua3Hr6P5QkhDO2haio/ja7BdrOQoBn
jPEbhLqHWGZywpkf2WY2B2aAKGmH7glUYe9/gUuncbR4yHfzFqor5k1dDvrMu0Rl
hS+imsdtjVNje5jYeDpsk6QdFdkPNbbIbciFxU91n+D/lDQAm1XIYbsS12D/6mE4
S9ai9I5wmNg/vcGDl2YHB71HVS2pt5WE80Lo5QVbh5hMqhlO5peuso8HAwlyDC9h
KdynCLKUZv10LoI8OTXVGV56ucneVE+GRh7KTAfxkMG6iIAq+wmrTcDL4zi+6xzg
AMnl0SYVX0PUSIO4gVRdbL3SqKPfizMFhT6IM5LHh0ThwWRDbNIKlArZG3nMKX4V
GFPuX4fEMKOWf0l+BK653uNKpTTlnr/e2z+fmssPdtAnaWZTEdYJKNa9hFkAc2Rj
/BP4vRgdGNwOqoVKXlU7eQkwvO5CuKsJb9YSHksB8VyDfPJEyycKscV4oqdVr/zk
byqz1o6aynwwbu8r7zhHaxYlYC9KAzH5FTT8Lm+ZquQpEUcSfNbXONzNawpg/vjJ
`protect END_PROTECTED
