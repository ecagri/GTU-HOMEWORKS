`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NEepwZOJ/mOmtxcP1LDtMbFzZl3Pe9jt2dVpK2tVF5V8EWK3JaPHr4a0OUcVbFn1
m4axtrjKGXe6NP1rRFH123Pgjv17zKb7KADF7/wDThrC0/9DKBHrwQEyZkpuFv+F
WK940Kds0k8gQAyL+NXCGTT+D8LkY/ECc/fURWVvHw3W/ohlSn8xFQgny9yAlbqv
AEBtq//JeUN5khVvWNHG456D1xnTWft6/ukvAa4V2RIVYKvQ8e6xAyyxVMeZyQIi
OaXBeKcEb7C0Lf6K3xXubBMYcWVmzxp9Lr7pJOBl3yWX/1H1Jk4saYW93MbPtmBL
1iEq/ufIDqvjLBbK+U8JMWqd7BTP10o1hspPRBZUM091nZsmPNYAjmWpRWX0WcrA
xy9Kxy2gHdI7NRu57mu1k2+6G3tvcp8PpoGGJdNtfOFCdbXMRHAO7JLQpv52n/PN
SMhtWmlSWcrDSUfDU2nqWYkr2hao1IZYfKq2Ka3vs+AFn4CaWpSvDdndG0qy5+RL
AJyUc8pm3Pk1VwtCr1lMdsXQ3U2NbcgUhbuPENErsx3276kuqoVxXpZbGxDe94jI
+rIEvPIo13XbSkVyDeNKS9IpvG1YELCGjdZVRr/uZbHIVEdIKiwfiwWAa7aBdsNI
Ky4qt4O826sl8wSQJ1NE8JIeGGRDAolMABHr1MQdlf6gB9ibODf0pq7u532bKcH/
ebe0qWZDTe4fDbbKdH3cxm87/KoSwKU8qc5x2S2vK1qdst9NPoJfwiTYeCHfDk2q
9Rb3CfzCaXvUynikQlTvqciJPceiRsDe8mXPjBoX5/ILcGTJ3CcV0oqIrDe0FWcH
7OXek1/Qnr4JNloNPi0IqCEq62BG1GEGtgmzBOGBChkX5T9JsR5h1K2KZj23J9B4
Hr/UaA2rD5CE6a+a5Vf0KqR8w8iCuMdCO0/DIPFUEkhOUp1ExhKC+21wUl937WXT
r0i/gAMlyoXNIY32m4P96y/Ow9HKzRvJjQ/kIXGOozu2Ns2K5bs3e3cVGaQUU4Zw
MKN6WGvTNS/IomIubkT6GrELzqf/P8nCBe5ELoSoUlj1WyCWzreCTDwgG5jo1Gea
YpgT36dfmiOfPmJgORoeJVtmbjgVrQdIBRv2zhVspLYYELq6sOXLG13flAUkFzST
UCfxBCOOtcCoLhKa1W5ploHNiEmk7eS9RMzSEsM2e8Z/RS+M36h7MnAvLx7wyoXo
ldUMPg7R8UfQ2jDOqT3okfGDyDM9pSoxRsad4YZDd3AKheuIePJlA4WzeG9YGMC+
rJgiC+P7pvmf2RPKui33G4i+Cg6YVFeT5zRQJ6wCq0IUeAoqnvw3am3Awfz3acFy
BoalLDRvrsaFL5z6ZTDBsMktH0jo8IosgUyfMn1jZz/+5ChkQx72NqjcY947rJEQ
WgMaYUU6vCuED6BiskUvHTHvxGi1bOIVLu/zJec/4r5nTYcU1b2t5zpgDNkgBKCk
`protect END_PROTECTED
