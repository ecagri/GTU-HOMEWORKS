`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AfNX3i0KObolrKRrHXgLBkkLwDTE4ZJ43Dzi/XP2EzByajMCzVHDH50zhbd+5eUr
zKS20In+pzkIY8kmsMqqeDOoYpzQik+Ms42MoMvQA9Y5Fy+4sKLnGAF1zU7jtZZN
iAvcmUU46ZZCUu0NkTtvjupB3h6AaaKvUnmMEi4Ojt12WWW3qA5RlNqul7A0Wvxk
7n9W4zHZc0XkMUE7vPSl/pZ+zYnOFnAyQn8OZmpB+td84E3r55qwa5NakM3Ay9ga
hr/IWmbNbkyGVPTz8WH23RyGLMvYW0rlZTEaw915BnKy2vEWbMSBgQJcR1Xe5Uye
HqY9XtjZlwpoG+EmDJYvNXA7kXVKOHYDwGuUFbdtTWZlfVhurrNiOQgWNDlAJb6f
1AKojxPtfBrTRNZsiELbBo+xJsafyTjKRs2olPfX3EFnx389FJVoo78cWdRBnvt2
UDpXF1LuQjiRMsHIa1geIxjXnLSXLXsGavf+moTR/A1y+mxgjtAIUm1GWO/YhVq2
hyYRxjpO/ply/8ohETdPjLjyuyUCE3w1UP8l1iEfxHRlhjQ1nBoiaA0zXCM2YZCt
/hOuHc9Anb/UmilQICiqT6Jovibh1c35pdEpFqNKUk66aTLZ24z66sjIQt475PZD
+6YgXh642UwOd08cosBo21GpyRr6cb3cWD2tV8M2b4lUv73AgK5N195MvgEvSJ6/
M5hNz+oXVETExgrXSjhr6o9j/AC3egFdn/kJFXp5EZbpeOQwpAq8PwpOP5FRnVdg
XOIH3rruOYxbigwIgVgXu65zDt6Iqf8yIe6Iu/1+FLsDQI52miJ4lcK8pP4Vdz+3
CbyVnE+jQwgixG0Tufvrl9t5mrHhrPU97SoH2ghXn1rXYcqJRzjJdtmIGmLJsvUs
KEfz2Njv8Rbtd2dHJFNBki47LwB9LaP88FsYeqH2gz4aX5zY979BiUKFAP/WCNQc
jM+jRkBot5IojL7vm8r5eJfZdgBYvF6R/OfvCJNY4ApbsYWkSHYNTNn2tMYGOj6f
wy2LhzbBru2wbZ2NFDd3SaOorqDMFPDzt556bpjYCHqjtXC8prh2ktgQQneRbnK7
PxEhPXkBnoEO2/PehQKSBWfyRQym7B4g+3zP4aKqLePbz6MyrvfyEU6TMLdRUspB
cvbeTFRm1lnBIkPUA8yy/yn7A2aJ6Iksnw9o3u31igu87DsipFYQwvczuuZv51m7
dGVfJlzfXHTmXYzu1kXGha4KbRQw8SVpQmztzek978MLIZ8DZ76Idwl9X/veP6Rk
Re6aloLI0SOg2fb8NFa+Iedx6usJlULi5/JCVSeFYm85B+E8FvQ/gb5ZlUL0zq+W
nSxusUi/A1uaPe2fdX+pftUw8TPUpQCs5E7VDV/mbWlbV0E609ZSLKoiW3IotYZL
v+fOfugQCtFBzooVl8z76TV3q3j0/YHE8ECtk0c/mitxbmAUa/wlycig/7ExSsue
kiH3MVgprmczhbeKVzGN8XEJ0dknWumMYFPYeHrwnRKcwF/FKUs+A3Db+paw+wt2
RINzvWhLH5VGdfjgj1H76LqednJewg6Zn23/hgQWApxD+jM4ebni8s8BodXzjDBI
t3ktC+xS5/o3H4XO8AY3VnFAIJdjXdmg+pzzqXaLW2V6sKB1jHbMr9yDWXoKSg/7
TM6XFrxwDuIHnw+j5QXvnhPdlRLL6z4/IAcwbkuCtYtH41pr3EjqWkCjRu4pk4Lb
CeYbsPbPNkrx4qfCcRTWipJosOZPG6lmPxTq/WKqhnYYfJMUwrFGin/jBgclKHxD
2a+vKcxMxtMrb1OoMT3q6JC7PgnqYYAsKm/j4V29q/n9uD4ajCJQtJhpTW2gs3NW
YtXqutVPsdFCnzSUz5i7jnCrm0uxsG0YQavS4w6d34m8YOqWx0YSodH28W6cFxv4
oYj6Wpi4YVT/k/vUTsE4pMSbXXOqr60pgUoQiM2VRJSzOrf8Gtmg6071N9TlLzWl
hh9aiHmfqBJBm1W4a6vX/v5URbjH7MErKAZ53GCPIy0KhDsQzitEOLcdLKMMG15B
Enc+++Xd91NKNqv+lTYvQxMthEUS/Lpz7PGFvEnjMpDERfwJAAlu7lh1HRRzqBET
KnFOtF72cXEG9n9ZM8SIotf5WH34S2PrCJfVSzTvgqsQi/ec3EG1rC0wcEoYKlPT
HIAY1lzda+Po21B1PWyuYoE+J+c5JdFjR+2ivKPcZgd+WtojNSypTgMcuI5shLJ3
kfl+FktRye3m9hxA6usNPEzp+fhRrai2BzhfRSkJJo+5PB6pFIIvfy6S3oAVkujK
JgXZimoptRocHUC6Uj4XRgRcnhiElKP5wyjbeP4+jpsITmaQdXRrSTMfOUmZy9Gq
UVBry5VNGBsoLnGLom0BzogWtGNta1O7mFaGDya9e6vlpQ5IEvSXDQOCdzF2nHbC
rkCNOmMe//Uzn/IHP3VkAg35N2ajDdvWnOnWMoOGTxwEPYjn/9RYumMAi1PQymqK
E3Jn+teahJp1Fqku3FiU8eP0hHv+/WzHc3bisqFRsEC3iJNiPHVZl9YggRJH1pFA
4xL1F6zmSZnt2ht4xI2cPNVjUJsIn/xWGe8fek/3l9ydkXIdUWVwn4h87QBaprdd
X0sW7eo/J5RjJZiqoQuQ0djPl9FbMn+A3O7mcLipDKR2gvsMFkzNpGBNNZhvthhI
zIOs74VHCJS09Rm/zNPHcfCD/LQorTmMTkoXJwIxNXoAyrePvpqqx+sFSZ3ujVLH
SRCxlhbDhJdoYGWWE586QqaHnfy2yWhBEeXZU0X37ZEpCgmJLSq52E2Hrp2A1ubi
nhAFKVe5XEBwUmR9unEpmaPw4QuXhNuCNB1q08yNY2pdCWd8WOhE0udaibdKExIh
UdGg7eS49+MWd4PDeF3IednqMjFAtMQzsibBJtIX2f0k+PAOpbT+faITyyjroOEu
+wofEJiDs2V8+FeNAFucv8FDlWwZeT3WPrtpca+U1t7/UqTcghvvkYmCdzZx8sM+
rUfZyhVhAF1xw+5c6vmXtBhIlQNqnhR3DLQaaDK6vi4K2IkWfTgsexlSOJLbV4H0
QTrdDxVUUyjQhuhqjAhjVZ9VlYkh6n9MWCNXDCYyJHYlPjm8A3aQAYtrYbFSGi7T
j1xMM/+ayd/tE5vJxDNzNkofoAWcfNiZM6NFeYOKOXDnCkMFiOwwbO0WS0MJgHUA
ePGz+TE99Gp/l1n8SenOB07gT0nLjVjbZtL6/b9ZnJoG7IvTRlRMueDYNNRX0KGE
vnRbSeo61ee4U1tFxxj5ST2cYE7RsYNr0TCfiIh1AercYhnvoSL0QcTqFy5fXLte
w2DFp/EnkSKQNn+8a/FhLTPIPvgxH/G0/ULMTMg4G4qdHFz4MywvQcZiaHNo1OGi
0g1Dke14cY+lFUq2LZdIVbu2D21wZ3nVvORpHuNbPSMSyh4X7MjjEW98BsZcYqC3
yhC0D7WnWAtR3UmIPF+YKy1KpVRf9nttgYcJIdFQHEmDhP7dlUbeOhJWrupW4ACo
`protect END_PROTECTED
