`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kjjER3Zy+SiHPDw/YPkm0XveGy+BifsAAsTDKk2fHH9Mw1rmk784vpdhn0k7EE28
+Ppn4trEqTHbjX2A52OP6k9ci1aH3Bh+QuWsSMuLLIdCx+fD/L5kk9QiJ/utSy6C
sdPL4jTek4PHirheoO71FcDPX2/18u89rqk4f+pxRGEib+ZVmT0fc4ntPHm1wuTY
O3Rk4v12xM6qTrOakW5timI+3HAYJAOz+UcPppP+x5dAmwuXnzPtVbbSi2yi7c21
QOTpV7fdru8gdDqo6IQ5wEXiLOLOgsZ+0LDXV8kAWkfykFtQ+cobXXn3z2ZbIvaH
0VWhLQz0kVr3yio+a1HSdncIcJFbTcc52ZFveD1uhMntGGYIU8YtTUOlpZmzn2Fo
ACayKVsJ1R/gpOKYJi/nCGG7GN44tGlKHhJThrIXQEGTkLuKwHt9Xm8lAYenTXhP
a56WbEKkdZ2WIoS/E9gymi0Xvd0tNvBh1ek4piGuEkWVxo/GmxqtWqYUWCUT6q9N
CC4ddWKw55kvVzIeV5I6qAzfD6ikSIBEb6mj2vhHfjbblOWUE38oE13+CIattVIx
BHUaiPFZuRJa6rd3XsBrZ6KU05VKPZGQtsva+YCqaFBrUwyXaamGfuTanRx3Qtsx
Q4jpnpATEZRN81NtdIQUyW34GV6ij5c/oFrxI/pP29pqblGeXY4nckwQOOJW+gjS
gpDuI0NZcQjjgGaWLaOMWT6NqfVggHn5DYuG+zuKo6ghIsRK4o4VcmPSB0PwE5qI
e3emYrM39R+3xtfPA/SAmLfjYyfsKA0+VrMgwkExhA+90UCE1U6CfiT7TOf74cEj
+IPS/7/OWYH4TEK6fvoHGoLidhlDkL/9A53Rgkvwd/1C/ylxQVNXaEY7AZUGjZoj
9hpAkVCxwv23NTrVCK+aBOptK6frlRG+jWbG4Xnftd8qGMNZ1FwPdQ5TaMvzjNzA
ARdopzwLDZGNKfy7LjdNeQXmFJpH+xGltf9kxi7py5fCPr5Co27k1+nggRGX+MOj
zf7pmIg3RVg/v8ZdJnLk6C+aHBByfu0GoD7d/5D5uULIHIkKGR6NBlTSCatloQlE
QE/pJr32pLcE60ZNB+Lvuhp+rIvEeWtBvj8N3NQDccET2FptbWKybmRtgpQBnMCy
mTA2NOetiK0lCM6VPYhOjoirLXwcSaDvB0FWoZ4UAQur6eavn96e5AWMG8A/wVm2
ttMwM3KpajeTPAqY/KRaL85P7xFT1KXFZlijBcfeCkMnW9M0mhefJWROSlh+wkJh
WkH3la1vjBvbOSSPphuPsvA2w3pnTpb5+5ud1lchAVVGX+NA8aFEjPr+LhDdN8Pw
XcCthQUOynDa742hcp7zjc2PrO+xrSKjMXTVtTwol6tMUHWPz1aUl8oLCkU1WsjH
NZqhkmGr7NSsec7iWzfrMg1pxZgik066QMJun6eM+zdEq8WZ4KVPCjBtpWANGvnY
vISGlOL6HPYJsLtkel7x2OEnI4V+PGwvK8CPj8kuraHOzDjA3TjZuGpWD7jBzwLW
sKook1QKbTQbURFXqWHreR95TYe99PKxzRHD5AJ3ZDXNsQVpTW22qNDI+D1xyqGI
4++C0kAV6mbd/ORPW+0xcVcreDbRs/R8wlIRyzksNGkw6TYVJP5eQPhWMsiY/VkU
4+M7yZ/ROtsZsO1rn6FwBJm3aGhN6InGbgxk9ckqFhLDcqOF3fmAbX0ZYmkppC9M
kVSluNzSZEhWniXRskicW9Kl2U7errYzSxFkcnn5l40EgsCKO4rP8qXsJqbJ85nq
+DTyfugHx5q2cmKoFkzrxmk7MfcPJgLy/VodF2YHjjwL1Xhyo8H0fMjoEC9hQB6Q
RySjTAXiWv4MF70En2YeM5BswGri2u3icaYYocUPBs1dL+0O1rb/1udgvNgqcT/M
5cxmOodilCmkX4g+QotLE5FPebqpjoHfJ42kEFy2EIEXvTaG0DcITj2b8jOactGh
CW1PwPg+r+DjM1uO//n5lRGk1xxYUU9HAgQaPrryQttP422uH86JDd+VxqfiVBBI
lhAZ+u41nRaaNk2TH7nXzEZN9e0Y7G5F+AWZUeQjO1PuzjbR07S/1Sa2QlautGxm
t4A3slVPx/LUa7qlzUhCfKVZaz4QoGFel62ubULAF/hyGfcBhcLLEa+A0fehdvJw
Wbu6h3sO4zQ4IgYErwcYE/iGs/bPxSqx+DkbS+gCJ5If1PypDN13VaaHhoVoXL48
kZzHGmOzHIvpqemfX8FMwWLySeMhvKgBBKJHPG6ds8rEGgsGTjQgg7zF8djlhihx
/2fIKiHvNDnl2+dVKCAOavxCI6fMQdyXYXl7MgRrbLBxL5knX7ipdWq65ueYcp1o
xaYrUZdd3wrPi/cPvsSBBni16fA04FzslDuh9gdHmGj7FOifgNXQtGfKEGFdnj5e
yUEtzG+MjFKqRc4b8w6O3OVPsOr+hLoNPEjCBDtnZoWA27a+yeRqyR4BnUv+oUKl
QXHWRhcttWBW2j1V3Rn4zvnZDJV8e8xRWNxRip771KiZtn7MUHKcIH7KCfWrTFHZ
PJmQ0K+IV6F1sOUhznad0s1gxNvidU7CMa1ni3aLLLAuD03+ns8ALPExYRmNedNa
FKxIfnQfXHZFyAviDAJrjTUFOVVWSk+VFeGixuVS9O9tvH3vLS6S8E+5KAcUBzJu
BBWCZ5A2Vu8cwJ5zjmI52h6Jgc9uM2CuGMt2bKez3zB+EIdqOfbr8PXi4jR7oWZ9
LMefJDE015SYuACoMfTG1tRrSmk8VKJmfBgiL46eQfmNnO//lBLevLFvjV9kaDIY
47giQJgaMwP/58alMxF14v0LYkFeRmu5KZg0dqLXYSHZ+xNaeOyQ1xqaZaSjPRFn
qtUWEYgTj32Scr9zUXZfNSApciXAvYYuJ4rHZUnq3EaX9RhBKdT+3XqJhyp6BfCw
AcTFPZiLZ2Vk7508lcdnoxKeuvVT5/cczia4cXbe1eeFkYyStCGsiBsjMXNwBgu0
BclduuELLreC8+36DbJBlIopVJIOOpO5sNuJBHmgXEUivWvLnRg+9EPUoVFt799n
k/UysOG+MgrTyRgNRnttsCRHaUdyUJsIQERr0K1xlLc3mAnOJ10792VFjQpMMFu7
W1/iNP5wdvhaT7nyN7JpQnncSP57zsTnH/hRWGcg4NwdhbmWu0vV50rrXtoi8Slm
dqsgKSt5AS/s11xBzKgKov43KrRMTkv6pIjxP5kwRnOiPouSL+UqRVQRg1FBHn5I
0XrYLMVeLO/donxUhGQJsEpqAHq7q0MBV9xtQfmmjq6VgYhAR+C0WYRu5Ffl5Koo
pqTaUmHYpR3VpuupbLAqqdm9k6ChjLbw4ZiePrSH1Qs8k5koQaDcSQmkxLxais5H
ikcNaZHpgZJNx2bZK8aVNkracO87Q5/LMR2iL5tCZtZrGQAWvrfu4MYtu6G//Pn4
/Oo/J2G/ac41EnEW7ddI32Z2VS8PfSdN4ITAja5w6h2nHTbf1b7eIERwYWbpPl5N
i7cZgnDmrrTL6eboDysU21bP+dOWUl12Dr3ZLNvj+h6ywN7AHaeuhuoOqWjxonTR
pfPFPvVGk9ptQnnwMNpzXdMaOj5dNeP/TZ8K9Y0TR3Y1VJt+/iLOX6k1qmqhcTFo
FqgQ4RzOo6LvvryQmp/lsAhXQecG7uuu1j7BGKOsLifyxIUvOXHlUp/JfO3wc9jE
3xIBWzWRLOXUqioJDNEzFkceV5ARENjgrMAVd+9LlgyOjl+YfJtZtTHJv+F/gImb
8VXPU32s+IJ6I1YRRU4n924KsCge3VlVn8CCgCE46pFu+5DaM7KFBIKvL2aNxIrQ
MFKsH0Vqbdx6Rts2Ac9e3B0oPTEdZD7I6OfXFCqh5raNG6uq8hcdFqdhAIcaCK9S
/gPRfmKSJ3wqC2q0oGFjGxWulYTsDPv0TJaAZ9XUPWtTMT1Z21UN9OxW4H5Qd/FD
CP8ToLukrYQbgZhQ4hbthfnMRMa+Y1xD70tMPiKQ8FGq2JWkSzjD0xFJTrJ3b38O
DFma23MbIWOG3ElKk+1tq0Q+tVf0v4//Zkg8HYOIl3bxckNz9Icc6V8xVOJh1CjR
v0N/Ivae8TWC5/vHdsWPHGUeTJQlpr6AV4mdqnlDlaWm3EtZuq8AVl0d0gWNIfve
Fr053Hg1Yq/ag+Gr05/5f+RTzRVS8ghAcrQFKGYzT0l6uVa6Xfgv0To0QDmEPvKO
39VV23yLc1HlQvzLqmXRvxFoE3h65pdO8/ujddukkpDKopVANJAmeufVP1JRGn80
Qx22DCjDf4+7iKtmoY+0XemAjlXX0FIAkpfNdInFVNY5equmwGve0T9gK8/dO6Wr
gj5FaRzt1sHCaK7P2HY6MIc8nYXbvtbnRSXwSsC1JDNHEQ1c5Xd7NlJBdG5LKVqK
E8OA2Sx9oHXuvpHeNDv8poiQlcWLh8TKnNOdUewIfJeV+Ypt6quf/Y5RXTl/HvEd
og+LUU/wtmhMIl+t1OGhGvqQOVN+d80/1TyZDyB/0nUVDmrbZaNEj/HdQLms8+Ys
yJYwZp2J3l/7dRj2QU+4oshJ3e0zVxr38Dp01aPO7X0LuYx3qQdXv6k4NUK70XPm
6a/WTsDW/7fdPh6M1yJfM7O1rR9T+P/aC7Lva0dFn6/zNR3sni+w7l5N0twCbGGK
LA6kDKrDSEfvGit3Ofnvl1q1rO9t9P6u97PdloB30T3r7c5d0sQVqwXP9fCOG1IL
kuuRquhIVWmOmjInJu136GvzAb2JNCaUGl5Q9dXiePcQOSa4o/vZU477nNC2UX9T
Aw6cmWPN3/jlFMSfBbGJagpOYN6XSrSFB7aKKv5GKqBJ5qlqh64zm775FL82llwJ
AGOLnLbiGVSWydKY1wQvWJBlwhuTH6IGNH2p6Fzo9RXm1kTVMCEZEeyxT5ONC4l8
Sj+HJeU4ysHLTuWl+x/mB9JTI1rgXUQOFSL+V9CY46u8BWjZkHYv2Bk+57N3ZvSD
eMsQM0wnEcSCiNeWUPRRPqq9mW9GjAtwpB46Cuk8HBq+5TZVsRhx/AuS3uaV30ff
djfih1T7foSgUYdYNorkesklMGKG69TQYsgwTgHNAT52NYb/V6Hn1YiWno6kIB5t
Zoq4g7GCja0D1XV/MO7EBVpJ2L/5mio1lUIKiStF/QVb9nZkkm6PkaH6vfIgrZwE
gZ2EcQsYjU84CRMrxcADj2BqDeUVJqC5xaStG4zI67IdrWbEAh3Smk6rhVWiT95k
D4nujnwpNWnDPIVAA9MroB7mx8PBIS4mclND89Q78CyPNUTeTKgGV5GxmqKXuBwE
S3BPuUwF2BT584+ShSLxcgpoWoY+CLeJn77EFjleY2Ztkx+G0e7XM2IOd2bBgcqA
ZLruneFS93EnSifKp2z6WNK/XME6Xn+SFFNrkEXoDobnwxZ9Vl9yUcIs4jN20ciG
HNAWpusCjxKKnjg1bWYYdEkioXY4dBYDeZwImhhhXkvW1O6Vn45akoDqphJ37GjJ
Jd86R78XFwqVKCdSxiy+GW/YJj9JVV8rGMhVgUxnknlS6Q2QtAZAMfkPwaGDw6vZ
oZfnQjFA3ESO6GgbrwH+rcyL5GFm4xF+0qpUM+l5heFzsiASc+OWxTscxycXOVUF
+601e+7Nw+MAroBeuN/hJgmwfWn0pOaklO4fABFQsDCQdTfuAD6v5uMIeNn5wbK0
6L+lG1tQTbSm0ixkzFn89d7XRukqUbq+CUmdOqr9DUGH0creD+Y49QMXpWiJJj5N
v5HLY+ppaaj81xcG2xzOlnSbEI6uW8X/L6rOLEW6uyfVIK4YKYIACnI/qOiqr6jS
00SLp0b90yssqmgV6+L1XVztEfbOWLzR2snGhEoY93KrPUG3Jbt7vBZqe7zRIP6R
20ZX8QTIjNz/R7DiLJjIh7N/78D3YOxqVPlp/Nol0EpEArJ8LFMh1j7Or/YMgNDV
m30o/V8QzkrfFDEB2hYt9SrDiS4wsT6nBp67RaqOaUb88tqfolpP54YbZXf++y0r
Bt97GzS1lokBp3sokktPpsXW2dJ2qZa6hNWQLXl4Iic21lP8eHndBRuUJKmTg5To
keht/Ayss+zW9ZnPTZWUgtfC0YmCL4Y2zAu/35gb+NSulr745QlRn8Y2FjmM0/Ij
B4zKDfBkpT7c97P3PYCGMrR1oiUHxygrtnCMG9YQUzrphAaQYbwi7BnhTXRjtIFH
nw+nkk5mH5BWiKG8UfmovotIxSV1NzRZhDztoaBnyi5BIY84VA2NuIZkEnw1u1dr
Pgs4tGLLArYRYFTbFbtuVWGOfuL8vmyi0Dkm2k1c4+r8T+eXUfw5rjpvInOkAZT7
28zMj6DYCCz0msHl+nq+PgwqmLqkGINPGj734ZwbSf8tfbBEw9wYDOxj4zkHfogN
FYMlVddDH1TPxioj9XaaE2/gFcXKw7YiP1lBPrhfvWOEs61QmQnRoNFB/WUe8YuA
+GWxUk04htdyBdD7WmxDmNhiq0x6nH0sjnStgW+TpsM241thakjrA8EpxhxLRBUp
PykJ6FGVkZpu/HCIsu8+2NaAfguuXuVjufRJZO+OUDBm7ZBxPenTcn41nvKJ8qSu
6knDHf3+R+sqR+/DUTN4xx5kIIkzzSPh34OrIoy0fOTXwRRzBntwY3Dx2As06Eor
O/K0qgc3/C0cL0kZTuwktVLb8rW9wmevMOcJhw2SSKoGCCjx9H9qGOZ59bDeHrMw
8o8YJoGQFPN5lSjc5apLMJQYvPXAsDq+rfWBzE+nIKK27kNA6Oqd7oF7khhKY/MK
2N/kpCnbhHxspSAjqnJOE+uv6DgbmUfzeaFQm42WLTkKl+1MN7pe39ZAQ6RtgG3S
CQQnL2N15zs0398NiKs3W/PUuDO7WcR54bOeGW7Tx92EP62hsYlgMzvPB6Bihvte
xny41PjZ0zDDAI2m5lQojjrr7Zrbl3dn4KcSeXULjdz68w32LRwCV+wtboWcD4N/
DfdtJxP2Kgyhw9JKg3NZNavqJahA+89OA3zwHxzsIkI55KRPRjRPNUzslnGc3ITn
ql232ozZEK9D2YfWV0kVyAIe6h3iUu5HiTEdmYu0VuiFMkB1qct6mqTzeyZ1cYG+
gm1kscY4gqNWubs6bCp/HkPpokOdrROi209Iev/Kz78PpsBwZeqyfF5iUtw/29RJ
0va0k+am2T22K94CY6sGMf8D0dnP8SxEX8NWopV+X4DCxgemTBdAaC8EejpsnuIt
lCJr98mVzPM0cfdT5O39s2WvUcy1e/XhuXET6HkyMXqeWujLtcqFpBbzLDOX97rq
NGakUVnot0IPZhSqQhp3gnqrNgluZwiSERj4J3cTMVm/TOK7e9hQCeu8cJMaClPc
vJzzCreQfCxOfLpXOjSVMKHoXI4+2skv0ZHC/eY+fALSi5N7VngXC0f4zFyT9Vs6
jErWDQOfAm9yWxLKZS72VoWwpXnyJXFibQANayJD2+pNCMdQNKc3iq9AWjxKEwfv
NLThRYCXWvn7dqUqJaCWDPShBV2NMjtPj73dSP7QsroZA0IBaCj4hY/GU44EAW3D
HBfzFDEh2nP6LhOeI17le028jx8qJhxJlNzTwkKsycJTsPb1Jf29GXyXjF/eaUyZ
17XoQmH0CgvTJF+qHEcveuQUtT9TvKef0pl03NBBzufRRci02DTdSg5JutnA81PO
cZp1QVY95wTU1TOqKh3gOKY/ZkCAufF+66n85YOEwi3dLzXDquhKXg24gc6WmJyu
0XZ9WG0UdqWkeKJnf8KWHDtCDenM3xjAsM5pBEg96XKYmE0HybyLSwO8fdLHd8dE
cDocxJrmOUudcMfCL7VvTpX3yI31y7zBS/kn4mBp7HrvXe3bCIsDQJRlP45R9llP
ZT0hz2aABVMJwEMLCYnlbknwW+KzfRwITidhsUgi9rS/8EFqAb2+IC3pvDM3bjaz
ZhqyUYWkjSYQUnHNjH0rkSqTXKBw8dp9C58UM2TphoMeCDVOPHxi0ohIy91b4h+T
IbMYjBQI3yx/U1NRhImBGp0YQK703h6wPX8YS/x6vvfYMpwpU3LyEaMtotSA6cSy
c8/5Dx9hEJi5eKlVCKDyCfCr1RmE/N7m3pJ43IuQDy2zAEiDD/aimDrETiOESUNR
Uf62x6yErl3sV8DmCXme7MxX9Ugkm0oNPKUbNiL1KqPhpVeU1kcNRG3DqeJiMudV
EcxizROgBevBL7LCtn+dVnomCWvJ/BXTKm1o2SLFaNjFC9XpXVgnL+ug+BMzvuq3
+ETkXEnD6AkvKCuciJZbe1Nwv/TnjC9AjU4pNvB1xFQR/7Yb2r0AbWcZqlv8pv3f
lCUXylIat4kIHFdFk94TCj6+Ufdqfe5evwKOsHKPqoBUI5NYNTSQoLNmaPFbWQY0
pbzSL8lI8CzBKLVY1G3u/qcObm8P9c12hva/f/eveDuP6Nj/P9K9hVcRMTiWq02g
QEd5TaBe60MbdMQN7/yTCTsbKwLE1iLfnlBrVRMEwTo3N3Vr6Kj+QSGm0gCdRGAE
sCWdlTkZ3psgsFE0WbZWG77+oY5Yi1NuJ2Ts2R3wiQJjeInRF34CFG4lDXGSoUX5
3TPz+2VG8Ygv+hvWd4Q1USwq/KIqtDnKgO/milKER+e6PqQxDh6r4yyvEE7KY6Ci
HC8V1eDTAxi5hZaRnM1spn+TuGHaAprCPwLK/82XF1y3Ww23PfwDRaFGYCp5VfU9
j17EjKOmURoLoF8cPhHkDBon0UfgYgS5A+fYacQ4KzXhH5+XW/ABkrP6adc3JRAI
n9QEQ5R21U93KlZ30kyFdwnIZI/8l/ED2nYsuhrZCfuLruPdPhHvPwQoi6UcBN2a
DpA+SKx8M5YGe7GnLUP1q/H9qBN6xmMuvhpne4trFf/DJaE8eedtZblqqnVzdjFI
64i2+BGxlbnBQU+bCFCQBz2XLBrNTlfFd6+TnKFIO9yhkyyhQTuER27ezPFiacMi
0yAXre2hQjwYsB5WYa0+UPEKOLDb8EF0OcGyYKyScrXlp2YIeuKYFKeLH2vgpAS3
nHH7lj2OeaaDGlg7OIW/XTwPrzshILwZqTX2KoU6a+7vom4JaEOAfxbArNxaD5AG
rm26IixxqI2BE+zu5BImC4xtCLk/Y+nMURyGVmqghSrBlRxBj/6YGe15eiHaBk5n
6/+rMFIvHOWmbwk51oHzmRZ8dJRKFrEdjFEHO44vrU1mjJh3bFCsEz5/qGLIHera
XHNWUXwxvtk4aVYeifMQCRi/8u7Bi1V7dqe4VHMUE2UIG/a/kg/4+zsEa9fv8JsU
pJ9xZ1rQkqhWYc+N7Mq6ZqQtGa0lu1KfjKf43VkNxzcYWjglkMV0v+gWSDOW3t29
gmoPckW/ZbJfztiAx/hE4abYTzctGwGR0Ibn+rGsKNVsGZpM2yIe72roXvF20tJV
hf2LvtGZmDyO8TqyNQ4AF0a5FykdWB3NLrTJlnxifVO3Fbba5H/8BCIKyOM16Ww9
2qg9WW47WFZYij3UYY6IucNu2V+OuicAzQrn/CydbmcnicNo9he7a3nXk+mhdcr0
HCfZx9nNOJe3zo0VpeHfroDuAvO6oFuvtGU3zfQKk7z93IQ1rU7BMTToPxR8OsTe
bhPWhLLo9UmDUvAsdXPjDZykSB2+No6bs62m4oeYv6Bv29KsYHp4dNZDGxsBH3Oz
NDGdDZxSlNpYXaJ9IanGXNphkbVUDcHVYeRP4B7CucveBesh0/YsSucAbA1riOec
XPEY3LyQ2rNKmXy+Ns2iXn7vYBBmWftDo8hzlu2NQXRCFw3zCsgx+lcXpezlw3O0
1uyKhbRCUTXg8yQ8z7Yedlh/jUcigODe9u/s+gC/XWHIqNIrmV5i6nizi9pK7SFs
/Vo1IAFO71QPrYMpsf0+GWWqDQx7iyfnZ7fHSX94O4IzE3crRCCHk0KpEbbb2ml5
u1V603v0kSyw5GdLCC6ulgwPN4VfWVhe8lR9BJE8RpNt0JYZ1eQD/zc47oaixnpJ
UYkL9ziVP1Sde13BAgvk3gjFm1o9MaFAS5ST9lM+Aet9Pi7J8AmR6aHFIx7zW9hC
MP5PiSIuIx4I9K7VSiM6OvlZ91TzPZarGnofYHgQlgDYSPLtfh2iQGBzVV88xBFR
n9YGhpQXII3kMTlp/qnGpvi/ce2eUqRooempK/momm8pIpD+riJfbfcsyH2kXacx
ptlpXcyVJPXGI5reR85jEGHCDdc6TTPu0uqARjuJ+yOoBVdnAROkTm6vPWtKDXI+
ydQlB+Gxc46h7+wTUCKFzMxFXin2CXg0qWb968Sli2fwQw24RMPylxxcltzX6kxT
pVayLn4Gc8VwWPmqKALy7HOQQSu2KLXMG1NF0O9eJMAFzFbTjWrkYC7Rz9XYLrmX
IFjI2vHyuAD4FMTHguv0oUlzzueKqPJ4IEvQe0XG4J06p7dZq2A8k+/h52FSiSAt
nqS2GLj1/uHUL3yqWNU0JS9a7SCckN1b6L4vOVyNd/+1tuuorjHUiUNKTvNylzqy
IeFz+TSPAK+tWHxNob9OlQ==
`protect END_PROTECTED
