`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BBNrJE0N/umBY6QAKdHoawcyr3TVhRtHDVwPke6saZW4G6ua989Y8z8OGuL7xe46
ppJ5BuhWa51s2M7EbpTCu+rf8RhjE7+LrQIRLso/t0V0z84eMyVjNqDkMxnUOCPy
lgviDls3M67fRUZudkKG/sqcr1k2ozehW8T+DUM+8eGhvgXTfkQFkCUhuOFFTjai
WXU+3Eb0xJ9uogWXw165w2KagxOyChAFBkWVL4dZ8EwVOaAmttcy3z+G5Ebht0qr
ly8Vs+6/RkTZPiYa5EN9Mv5AEsUR7VuNAdOtmWx3x4WsoKZnMR/s8DPPtNbCNybc
LjeLLKI4jwXe6w6uQli16m1pnME7sP2FB5Pv7/qhFPFqRFfLNUtAvs9RBQbIJya2
w+hin5uphjc6D5DbbrPPuJFa/dwcJ/WuxZzLKbuOLIk0iQ/KhGjvZ0HVGgyoFn38
bLSAN6Hn3ZYXe44qe48xlPNNBn/i85Gp5WK361zjO3EvCukxZxgmNG2lN/zlvFbQ
deKgDx10PyKxD7Ba5/YQIsMpvoCFIW24zsBKNp+i0kaGl4Mj3nExB0GP1n6HfkS9
KuqcQ2C3gE/Q9n+X8nZBZXKB7EC2TQPZE4iXoom/deNt5Jlj+afP6zLF1QRdyeZl
6atIGJGm53IH4GlEuOzV0SzHERtWjbeNZIz2+A/QvIrXfX2AW2Hvi9wde5aAtKvX
t/ZzmvUwNPGV+KklhoOmeQ3j9u1FwNLp2sPaW+aNomQKfqVsWdh0t+cRFMvESLH9
kcgxZf7dl3sY3WIw4aZabhZhjIdDe1GlCudXOj91uy+FOUwZfv/0+iWkxU6MOk09
C1uDlJX9H1KTQgERjofeKogJyvww0HfcR+NeZSjdMHHJOOaJjqkVVZinEbNB6uCJ
9p2YpR6ptuP6zAMT9S2VAz8r+aVKophun3T1TE5dTGX0zKxtYKR3u034ECwDnKnF
EdtGgPM0qTiOEwpebjM2BPUdxxqByj8TA+2g5FzHTQ1nsXmTOknYQD0q0tkMc/OZ
ngnS8KQMTMudmFUgKuvFlbIHIAf4UazP4VL/olYRYDof3bgvtAPhw8TthtpNRJBy
SvDwrmsnpzKLOPnAPo05VrELsLtLbPXDgs1H8zQNJqlM/xWCBCSI/4+hl4zCyrAJ
NkG3vLGq7AyxKmgNhYfhG/zupyKRaFEzu6TU1J74ee6aUHARrtaNtuXSA4q1uda8
/dy7CCX5X5Ip7IdqF0JTUhpkaM/ScqQ8PAzyttkl21VeWCkOYqOTlre6nSva80tb
QWdUZ5h7FMj5eIqtokaukLwb12E3Tlk+9q4l04UjWoytzcfIQIgrOtzLZokNX9h9
6CZkEztieT8+jtfMN+DnZ6bjRKDoAsNJ0W6Tdr9p4nUymqt1bfhYbr4zKJMQU8Lq
2PevGllkNpuTV+aL/leX/ult10h6+h8m/55PgAEvtScZeBxSHFEJX3ZvO9j3vYd5
6u2HwPmrvxl3Jg9byx34nLja6jCgexz3CLyv6RxihbdQNIK+K5lT0e7ZvtNjU+wy
wsS2GIJTgg+wOBBghv87xQT4l8jDsv9NZlwqCTXvx1g96sKlSCPGUWaVUkDcaWzA
OVPYSXfu8whys7fxS6mCPx5CG8dz5SGdmGchflcH8VjxDCySgeaDgNo8hd1ZBx//
RrdQH9vy2AWyH05Ia99KQoWR51maq2yMpNiA8MSePVmvBDeMYct8i9YxTv22gzrX
Ve+rSZrn3CLLH1vZYqHIzXqcqUeRXOsT/RbBsccM5Awxlw1SVOm6N3tBJhXgLNRd
DtO3S0Cj3NYgUhpHUH4/Rs9BoVsbwCNlbtzg0ezfxZ1D4/FCN2o3QFjy5/hwlQec
sVbCXyoKOxtK+wyKfF//jO9+81ToqN6Mwhfp77nz0bw+xhgUocLYQ8afM3iUwTuI
nobTkbSntLGtSyUUMCXPpTJcCULulEuGs2Jh9/12yc8vxEDo2CMJM9vuL6U9zoQD
fivjHslCXnfzjBJxfKd+NGFQE0FdwyyqqBo/2f1yrDiJeq4kKqIlbEBWn9qtk3E0
6X4jawQPwPWDYOg0dqsTPgknZtgr1Nlrt8l/+Yc5m+IxVvRnyH6DyV3+KPbyLBEJ
3aNFnAr9qo8T1Nkg2fRHrNxk8jq8D0FscW9WEAuwBMeSsC9zF4qvdYx4OkPTJs5x
NegyG2A4xTyga/ABvrDa65mSlvag3AmZaXfY3kMszTFx+cnz/oNx/VFLIMr+TlMa
oJHgoYPwqfKt5z5B2M4MvWAtnvnoCcUfHfNtei40HVe0lZi+MdS1Y46hLCbtgB99
Z6+jMShkYNv7V1RTMuVDTIU7WdrBI/4a4TEZi/WwFXbF71dng4AMIcS6xEks2J4B
90zEqsZtVeoFm4Nuh2vUb/0zqY/Iqv5XEz2vUBq9on9xa3lxLdSz8z1ioBzAKw9u
CRL7VhxRiehqruDw0lgn210kx1K9qLVayF9MQUfWpD1xhKHCQnGUK+/H1ktIyPN2
Qi1/YQe7KY5cRyQjCSer0p9QTh/RJj7l1xuiI0c85w7wcN/t+OW7N3gBu8Z1BkyD
i+wWH6QYtBolFyf/ntvpW6F5mZ3NVzD4GXB8oGV8Vex7UJlD1DmHAFoJ+p6dkiO3
P8TzPRMusONvlK/VcQiUftMCBaBrHDypoOItYJxLTwwGF4CxstEqWCmRZRQPZWkU
N9oKWE9C6ZmQ1F0B1HIANIQG5b8QaiMolRJvK2StOrBy8m4trQ8CIh1bNxkGh+h3
RtlOUpdaJanL5V5uQj3qddgILAuODE7EkYlDRZxMiGJXGgjLwRD1Y6Q43HSqSDfB
b7ZdVbuLsurV2mo2Dn2uGWvThYbMs93kfzte3vsWza/UP04yqEJWz5qAZf399m6v
rXmG/B2/Db+tm91DZ1PdvBtPcukJJRz8toquRZuUdgVE4V9PNvvWiYT4Gd80myK+
2lE5ip2bQp1MkifXHVrpl9PKNLotkk9DRhN5ta/+goG71bqE4dHoFFzjWUXk9A0d
lSdIsKFrllz9LdQsXBwD2rRurA4vowTrqaVpmYumdVPp19AQGtyI+zQp/ShkEdqX
pjzYznQyfYO+LjClxasJmXkhagLt1lPzwKqyhFpgaI54PtQdsI/7A9I5KbwAj1mI
RPtRguaPXd70Sf9TrC7mP6skHWBmR4QgORDS1TF3Hf+6mZJPCOSPjqpEUwTy0LI1
JD8OXigHD2A/jJA3gfuzvZ4jnMfFGdQchEaBouFirsYd6W3tBR7UiMkCjIi33Ex0
CtbKb9AuCOk+o7fqN6YP19JJpAjPLo6rD3GDkKItMzzJFYYHh0wIBNdmhgO3spXy
yByeqC65K3+bebO3X4T6smukgonbu3SP4/hLFfcINYciP2lOYk3vR7bDsZOhv0WH
q2z3KMfBfC9RMtxeo+zzOr4p9Wu0L0BvToyFAcKAlCDYULYWtUfBenwFyCBib6lE
1Az0Z8f4yGggBtMFSqV1ZiZ7zFo6oNa8NuCcHE2D1rcUuY8OTC3Alhbisfg9TXfw
k17jPk7R95KtEZle2aCrjg6jxb7j3rKA2C1hq/lYbRqpcpZP/trta0fiM+Vy0o0K
JfKYp3saoITUgNM+KaeCstsLZSA3ihc8lV7OWXoHCxx+ErZwKoB7zsyjrGNd17vy
FS64XfqXNpKh47hDTpkeq7MEeFJyeOsvq0fB1lG0nl2RxTwTDkZQymxfeAkO1pJF
gn1wX8DJsWoIr5PsPPAh0PmQo8YOJ+ZKSZJJdhw+02T4iJfJLtfQqWHyK/pzIs1y
qPnJ92a36BJxfuLprEDJ/z7xKwZhhzYkPc83qU7f+Q0d70Zl4iSSzIF0EYVBmKyd
Jw+aS4hrfcJulo8Ogyk3qPVhpSbykbQLtsq3WOIeqBS0cp/Obkg+EvhAL6vFs/wo
8Rdq8tsOPPQzr9MXGTN7Q+hbH3pZS8kav/OH37IIo+1HSNR7NK3vyAIkqwQUabgs
Djauzq+KNw4Hqlnk3TYxjH6YJ8UzkmGXy+D2hFASv4FE/pcE8jzq9VGtNbRyjMuq
/eVYF6aII2vRGv9Z6wYRRdt4Bk7j2fIMTxpdOfTeWJSfaic0qz1b4cJyvfuQxZqH
x5QvKP0N/KusuA1vLjcBEXLY/l7q+VT/x69u6YxHI/T0bLbqNlv1dhjn6Oz7ZdZx
w0LJvq5KcVR7oofQdv07aEpQ/Qku8AiTbw9vUiMJFMdv09vc72UCsOCMJVAddiz+
vLiV5A+88alyPtG/9SDqqjlaUGbLNW87LkrMLchMEA+7nKxYNJPxE0w4SxbfaODZ
Ek0uTBCsyC7PxfpNWQur3URdN/Fe5J5J+qfScABiYkabPQZ+5gf0imqO8vyHP3G7
BJ6K37QBKsNocycmT5rbR7hRgqtjEu0GG1vxyFbp5WH1GD16DTiPOvtf8kL9GeNV
kT1+zyNxTXx95iPf1unwL5z0oiUkfp/hGe9YTgxFdOLrdKc8Buutm8y26ILfr/5v
1rP9rK5pmcDywb6D7VcB5gwXD2qEZzPBxf5K5ZVGDaJJDmAhq66oaGvVZNGlLG3V
n3pGXxpVMJHDgElvOR4goi0cRwpwZS45PhaqhFhuQKFQowGJJBbunhbwYOCD2FH3
J+zCvbYxy3FF8giNal4tpZeA2CZYI4gYxHW2g+c/N03hxhAsI+Eiw27SLxOApdaO
Bwm/F7JU6B5LhfMMWn2iFneC9mqHtzKtA7Tm1cBp/K1O+gBMJ8Axx7a1e6Gv0fzb
RSQehdB9GrO4NAdD5jW4OYsNpAyvrOVU3QKrivTpU2qaQQ7FGQGyR8Y0ASxD+77f
3iRJ8P8VTku8I3psBic7AKjz8drBPJjeOVF2NLDrj8K1KXcFhZtBs8BuLyLokade
UOSJnWwEF0Y+cvQXzJ3w1RwlfoZmT82+B99vYCtrE5YO4L5b7xqPShgnU6zr1DB5
6uIqAyUlUDm+2ES1PE0MpTPtw3oKOek8VXaHIhR6hkCMoz1FZO2TLxsuZ+NzYIzf
jT4wvqaARUPz+Y7oCwimJ+0x9GaY7O6ei73otvh2mY/nnFEEaPZjx8peZRQGATIv
PC0BwSQx1Wo7Md0c4Urt615YzpaLalSzvkiNo6XfTNJXN6u9rLIIyp9oYq3U1NcR
uv9Ks2G7/qEdxjNaWBtjOf1R8hL64gCIh8hkRR8Wpqz7kLZiDqHJzcY43SDLZdDj
t8znAmcUTDu+A9tvd7k+x8g3WyA8ojzaY4afFCC79dubmLcy34Icfc0r6CskyMua
0uvSKr2YQP77Huc+RxHQgQ5Bhx+OxL5gIfbu4GrxgGC1+NGQquQxXCYl9j9S2SVF
PhbRF0a1QmufJjeDz6S55HidEtzcv4dqTOWp+pMFExRMg6IcepJ18LRZR8/G2cpr
YrUtgPaylPMq4Ry+h6TL03xQQUsE6K7eXYBK9CcxAcRM8XSAgBkzgAo4RCgApeCl
HpOhkx11MxNVJGMdXXQN6PeJ8HVdtM2D8k0EBvuMCVwmHJ82KDtA/T0S3eEZFbdT
Iw3+0pBbyxkFmoozE8f+Tk1Ca+CU/SuS4rJVtrDCxIP/4bKmzreZcKdV+0UO5UzA
8p5vCBJBYS8HiLdyDOXUTRwDC/0wO0ZpsFPrKN+pCHMfVNq00XddYf0LHCVEjq+i
kcvlObMG5yAoTdrhVJRzZFQe0JVKA1Og4N2rqkObFcqS40SkkrJ96lOOiMLbA7qZ
xNKYanVKCMgm4VJuDwbcCVdc/XdgEOHpAG8vPmlmE1uUGBZWs8KyghoY8tDJfepy
rm3OYt8MCNFAGkGq1HJQntIbqsdFARGxSWLIEdy/drn3jRtLkCUd3I1iYCHybWmv
K+P/mZoZY1CczlSykL3noufe7GaCSWSQDzrOYbbVeb3pkA5GEvhPH75aMy3/apSq
rnXpHibrktrlUC9OQtXdVdhbKiYzi0uhdbqH/zx7TMmVYy3GqpzCG8qwpqZ1kP5T
21DiRkQnyqE6MxKvaNeC6qJsdl+ZhlL7l2WhJAqLMFArlxnmnnj0NYEfgn/CAqE0
p51ptCkdVZJy7T0vIwFOD0djM0gyWeq/zNcHVGXZFlTsKqzPRhgVynzd94QxNIF8
rpqLIt3B7zAQqrf6YP5kBEPDaAIcz0hr8OjOjLf0wpxDkSwb1ZKgJeX+RKMhQ7DO
GWWMmOnZQpyACH7KcqWjFHqMx8JxTvsctkh1yYZfxkgiO8gmW622s+vg6MnDz4aP
fkn+mS9G/g669WB1dZwPKORjepU73XOHiN6f01mLdx6jlRCH98N0YaLCNIF1h5O1
IgBlJFWQbO6njPgyMpFD0Rvn8V/9zz29DdmsNpoju7bwk4+q3eq33pJVaHGwTORF
FC9pCegdcohrUYWNkULaXNEhDvRccbtjyA2geoHx48Dh15q8Vkom8uvipTZAPhrP
/NwGGajV8Jrs5OqjEHr8iMWVCzbQHjtou70Gc3KBDjjBt+9LNvA21RLFl6F+Iw68
GARRkdekqkJof4U772uWp4igRz/2fT8jP3OIZ5sS3i9K+R4Kej7OAyrFlYbRks4G
T6gCxXvdclnJkXUNyr+SHxVUfiktkycCrnwL4EY1quFCPgEg1OpOOWZm3s+wfIvl
wbp+ifN4KDrc05ccBPXUUSE06WE8nuKOLGe6d2uQPETGR6lHrt5ybGC9CSo6WP7G
jMZN4xQGcqei/yBhRkzs3w0G4fTDm7h7SwLFLWfY/pWJzwtteKZYTfVheGpdtAh8
H3ZstVeESmG/QHqS7sn2SF8TafKKQdno6vTnz6wIQiDL571xd/3o8MMw6YI5Pe+H
CYLY4PsMl82wzaNVp1k20L5YHgHdU4KtSwjb3wIftD+iune3IOGrR6d5zUumD/vw
gTWmGsQHRZTPBTsSZeFbZ0JUum4TYZt4RmQ6IGFUDjCVOCHT/Yk5Vxll1rS0nr+N
dlK7C0eNiyl/XV7SsF1mXF5zZrnEma6F9eMQSjW2IHJHyRCPKaafv9vJVlfcmfcq
v+XNanfyFXPgQBvUPASOJVTbbo51614Nv/64XBpP4hu0CnlMfcZ+pL9s2a/Gjvlc
3GRAlobTWJgnDPXIE4aRWwibPRAbkCEElR+vT9h0MxyS96EZUrpfx1AnQ1RJiM/B
rg/fbFk56k7qX/jPG077HSR6rpGy921b+FpOleeRDxZfQe37bpBS7bVheZl1ssMX
wt7x0ZoRvr27Vxg6fY1/cdpvjVPO1ZEsHGvRHXQb8Kz87hEo62V+EGtqfZvP3xnH
15BJ7d7dxyU+Fl0YlV7V9ygkL3dREIDtTm3T5Ma2qitAysn54wtngS9RQoE+2JUi
bDOIBuf9D7wT0AuGwncq6Z+I45SQhXyB6fpSW1kKSaXFbakW0wUbWKtC6FyCk2/J
eEe9cdaALNLbc9kr7D6NevzJXjO9udvHUuIbw/+bkW56obSlnZk7AERd6Kx3cOEJ
/89fdwrKYRtIsUGWAvyNkcDXI2y03L/FPM2eOqi4xjfEXEU10HbVQ0m+J5QZwvNB
mpqPiLfymYdu6Z4ps63D9Alk5/MXgCb6sW92qR6izjJe1s2e9urOBhFT75pfcVmB
aIrofKM4C+zKOri+BA2nE+dohPqc8GnIXu2kRgDOwmw4WxDa646OeUdVtsE4eHlj
0uAOshjmpTAflvBYb8G4YbwR1HSi/+Q98HdpJeeyHhngaIt3di80BOeYydc23/fF
5VcMbMjBz37sCBYqzLzBXjA3x3FklpbihgfxX3fPcZF6ztTTeHwrRe5bq8Jf8kyV
7xSoga6RbmsteUHL6Jz9tb7O2VO6/MYpsJzGzG+uLEtHdHDxuYOrJF0nEmo928L/
XuHDfN3J0NI5XZbLoKe3N4kk3aDkZEUrMc52GZCc6QJvuU4P6LF2tOMd7QABGBwk
d7u2Jp/M99Od1fvWkG4rQLRH01QcmFud7YlmwempPZtAppMOlknStWaRuV/axl3P
ehMPKwgotVgkiDR4s0GrstRTvF9cqvxc4CHpG0eE2GM57dIPiC1PrfAf/Or/A7CO
GlLDJGvE389tpNUfowkkaqB2KZFiwm6elyJuFUHs7078aYbQktnKp30/Ame6CDyL
T73L0QF+2NXWxsPpZrrYG7yeQMRlDxblISlUZY85aJdpEEpRhQuMzIk5SDY9Iq0L
JJGq/xqgLPvD1SFs3spDeHrVRMGPocZq1qhPEaQ+8xRSlIf3ZRC3MUyo+uIYXwSg
rHMHpiFqI+AO91MHe7JEP3hwFdXdvEY7WsY27QLUZCP8s9FEQMx2dIq43aISzIkD
BuQXbdp97ZnkmfakHLIbXUX57VbkcWJxx+ciKn3a5IMeZA/RqAlZ8aHANhif9e9q
qOdJ0jLhQgKNtFmn1gNK6s1mftTQolEhE+87I6Yp+WOn08CPkx2sTUOXgblOh/eC
MwIThMJV2qDhEjiXKXl9cE1oiPdHF3t6gtW7pIjDNiUF+7Ll+EQL+TxpmjYZT9dE
WXi/G10FEIN4hvJ/S5hzvqhMKEdbGL5a336gI20XlBgYDAjvfp1snfQpYRF3Wcb5
FTQINCkv2++cL7PSXZaQVWg5z5gwBMNAr6foWdVFbTxaaYJMZizomUn9dWaJfT1G
sv+Yy6WVTB7hdjVOEHJhyU67yxxoGTmRtIgWXSqw/sZDmGFai/vx7WCKmkNc94Un
KAbZhU9Zq3ginrmaVyX+/3dNDcy9sMHU3pXveVj793qjBmiT0iQZmzoNghVHgHch
gQmIcE+AXsctFzOW44WvMXI5rGP9L4q47SfyiBlH3NdPPye9KJTc/kEBMNP/uuWK
s3r1qnGMmJOL6HJzrrxRXSWHHo2h9kOe5RwgD8GSnZAq8TcFiZVemJ0dAjQzopw1
5cHXLRXS7c0L3A+yCS33IAoyYpB3HL5mECiahzMQ61+4spQsyEorRjGHeNd+daN7
RNu1XXdtOrvp3psaV9fL3RZpDtr4aA3G0Zf1K+oJqc01/CWcILc5xEFWyUu5H7JE
SuvaqzLEEPoiwW9gX9NYQaM/JLo6Pp8EW1dqReXQhCUQx2T8V4wdamhlf9XJrl1o
pEGjaF3lIK3wNmznr5d1jHXkhVv+luHqymQQF5lw0vmSdfZ/ShSuKAhnJ6BVVt+H
FHakv5c6A/+IuLY7E4vl9T3uCmwgu2/Dj2ghkmKCgC6n99r6Psv8pw/evogY2aTe
8dmEW2q3UpNJAo90BRaENrkhYPVa3JI5ulBKWD9RDCpqsPPRUFVKZiCNrPCLQwf/
qtFo/1riZmhQ48i3ujKJZIrS75itOvbgUYZmDMCeJMK+/9bOHsftAHu868GuDxJJ
gnCGekMzwuaNumZ6Mf52eIbuM2qZnnGGw1n7BTZSn+W5UAKksB9b0fOp37nFmO0S
ZUbhqCBkwd2iPnAPz4Fqc6pS9bdUa9HEpI5/E29ZgNEuhqJTvCs5cNss10UBtf9i
A5eKiwgwz0FagWaf9B5SCiAfWLgS7eWsJQnGSHn+Oow1nFXxveQgUEjI4qD2/MrD
C61SRBA7tWV+SG5zYqUarh2l1cCYJlmykNgOjkeWUXfZ5zDST+RJ84JL7NDuMAWf
6tn/vvlmgxiY0cLZzrOtZzX873kcuErco1AtNP+oTCPM7INfS/fLmc2wkjh0OUm3
7/qy8nbtOwtrxLa5sa+lGQig/MdabIFx6KRh5LRvXwPlWE71tRpjBdDTP3kp1HvB
WzVe632g65L9hF1p33JGEDw83h9ycEk6EljcBlDhGNPTddlGXqPIa5cHGW76Byhf
Yj1SdE5V2+pupIpDS+0+5T2bAqkapjpsLu1snBcny8bQ9vioLtZm1sfi2gJnLXKA
a2Hba7YxLXwG3oI6LuVFMvXnuSCWf76Rthy6tuK/lOLfJXlCN0/jEw406qorqDht
oBQyvh8W2KC7tqoIaOpkIgYFPWmdLQpS72Pq1ck4Mz3l61OoNvEw+R8UoYgLqoju
YvbVdAcDTqrd8eVBL1LpuosKQ5TuRloZeVVcNKeoodla3H7XYFieFBBOBWznO/pJ
zgbVJAopEjhrapH6cCfpJe5EiJ3zvlSoj9N2kPkP6NqVK0mmEJE6rZAov1XrDOfA
MrWsOUhQVj3KgcV1ImviweohH+4Oa+8uX0VAoGRcU4sw45v4xnD87o9iA9wZi372
gioLD9XqUGLaELSZqBHvMLCqqCX+8fPVzDlnujtt5e1x4z/x7yTC9xP1GPXaDgWn
A4a9w4I/yyQfoaS+omOTBPpduCM8UcU6er4jRBuUsvQyGVfO4ME1Wh405sRDgsBa
exGjqnGDEGvQ4a5PN2tDs+exqYcv4+q9Dg0YZtdA2IN3XVqcOvKyIrp7FTwNiZx5
zGaW0A54gnXjXLycjr96EyxQXFOFGJjgCVVierrjagOXHeqZsTQOMBZiK6BsWIMZ
LLuCrYaSdEPMxPboCbPiKT5TH4iJ5wgnnUyCyfin9TQvy9RVUq4OE/7Cp8hN8m3N
z4a5CCaxYsPM+mH8NCdzZ8UCVpodYl3SM2icNv92vdFQfP98eheTZLJVa7a0Qd8H
K7uzeNszi05Yfb2kd9TRcngcQ+Bn/OwjuzwKZMMFYZ5fBHpKSrP5uvFVQ0XLgkV+
jvHPONwqFHmNFtw/VRXMC0tyDNtXMM26cPGto8IPw6Z0Rt3sHsUiwuflHm0azMIp
BrAb/JTSjyTeCdMyouAfxhzAPTKQPCb+b+WvUz6becWUr05+OJ9q5+x2sFXvouqC
iM1q53MxkB8R5F3Jo6W3z88bI0NhtBHeKCxnRuUMXniS9f+6M8rF8EC71z6bgcgn
HtSA8G8D4gEDp8K4XIGqmvX4Dk+vLnkIYQwbS/EfvG1/d91hHwRiktbdwrMB6bbH
WsGUpluWxD/jL+8YMnpkMe7hqyag8NfBLzC/4vAS7Bi45Jracbp6IKQrV8LLuKg9
i/6fODiKYKwH5HZHhvKas4p5MOVcCdDNp3+BqPiXt2uZfSPR5byYOG1eLgPO7nX5
InMGIuVkvrIIBbp6ZHSQEhrtvv3xzUo9kK74sUv8dDIq6dK2+QH3XO9s893tqe+O
AmTk0qQPA84tKnzMM7E+czVC0qFynkPC+9sGP2f+vvyILF4vgqcVjEKcjPMCyIIP
f+fqwZ1kxyT/vrCSATdP5o1TQZ7tY++sR5uoiGHW997pQZJNk10MmJyvR1BkRh+G
SGoxrruG5cVo8j8wW1KSUlXU3n6lERN5O0KbGbeJSIwaIwaYHjmXfB8yIfjL78MD
HZQdVQc0z3VfuPaPbUfcR8B5CsBGvTVuloitb55cLDhrEhJ5JYYJvLgU8YUmiXzv
lsSJn5YNtbD+AWhO9NjzbmYlr1KMBbmpiXKdVD28U2Hsda8jFI88IE6Vv5vY4gyd
N/qj+UfpwdrmaOmrCW2GO7jYg3pvdWsX76YMWIdD18eI4juQxofW44fM+0Pqo/mu
lSai3iA6jox7ej/47RzgRj/pBuUWkyHNNv734a5M2H021MenpopBrMbXhe31fyKL
p0y/FqFuOcYIMEkE4ybrfhRtvBEhGXKjis3HTjVbwR9MN5YhNJSy2uZjKyNZUMD0
6wVa6lFuAgeT5ipJ2YHFBPu1f68Uv6wdpw3FtCehh7Sbt+xdVNQjJe1txZYFDDVt
rQsoatl2PRyVwg61mJkecvigiRBx5rw2SMprrIFTr64DTlAHXVDTop+nGowuOtkB
mMmf7WI6tKqUs6jlVaWplMX/ax+6BAtVoX5+G+24xix4AVjUfWq9i2ghvlN/L10C
8BBcwC75MhZz3RhNHIclTFLNd70GxYEiHUeetDYX0vAASc+LB9Wa0brb615akwPz
g0ACurmFI6DcuBMhvXQpHdglKmum0dvTdcc+DLnF8V8qdiol3Uv0HceWKe4+j69j
wcsJKmJ8Uo/ad55hEC5fdz8c1t6ZaNGRRVfWBuajtiwbQz1gPj9oK0j4sUHwUapt
a8a1od96orCNpjlMI9XOJ2B3ZXqpo4nZXBDWNsQUfnSxVUbQqLldcs//NP46ICYP
3LPOYAZRRg7R/kH2iy50OmMW1nvCeBSS6LPSuJCxGNHre3F9ZGxQ12HLUiLMxKZh
n23THG2e2rwPKVJPe6w7JZV1BxIzS6xmsjVKO31Ft40jUivbJXlFJ68LLcF3WEa9
154CqV/8RLWGJXmtwrUdxWDYjX4a2xFxaKdu30EE3pfnYlhH/1Li6Ym0iXhzZLuH
g3GzYJwOS+HUsbQGqIbyWrXN/DkUNsYlVSfWqg3SgMJIDMI9pDrgDErfEByGW1Y7
C5GL9GF+LtjGlYP4aC3nUrOQyZNwfVuQMTRkTbJSXnSh7jBCH6sc0ybg0KlpsAUH
Yg8Z1nhmJ9gpltQM5Ty2fdvfytMEqSPBqkmbxYwoj+RYLi67FdC3T+pxinvXuS25
TAzx7DpB4Ve0lmb8KyDwo09VqO8hC2PYbyYEWPNgvpDPX6+zu1V3dQoAgouACEEi
YxjYUlCHHrO6P2WxxoMPsf9jdyLDT6yn5v5SoG6h4MAvu/uO2iZIiA9hm03mUx9Y
8v8fIzY5dkb6evWaBseDasf8xKSMUviG3BASg+SKTvb/mniLc7n90CbDGC1FW2bp
dhBDDvqkBA1VdhVW/PfE2Xb4S/v3y7DksO6ySUM1JcjCR+AJ/z4AXYEvS0vCIM/0
IwYPaj4Fkn3qwSzmJyD92A1fU189cI+oDKjb5jOyAg2h+AyYCWQaSxDZ1bfcHN5P
IEubWkpmwRKHljtvab9S0XCerHGKvyUcuOPZ9zSbSgL8A37+NdHupacUIl7tmUsE
xU7y2wIZRucRjiYbjZ/6P47K5/zo9km7bLJJX4ob04SfU9APX/zVl4JQYoxvJKt4
bQK9i92OuUSeNkXrUbHx4WZvmjGLGUKG/39LFfseeXa3Csbm+3xSZabGF09Fv8R8
Y0N8c7khrghMNsYxWyy2bdaiO6MVSJPNCk7PN+nG2cvD+9cXYpo1E1mZprJ7M27e
Y+Uobla8FILTtGR5FTVM/kYeVV4P8yruID/SeqF8QaPEYwt9aFvpifVux3X3yqGo
yc/9+DsumMThdph4i330kBa5iq7KuebjF36m4X2I+4R9ns1Hjr/aGSQOWPLRpdUL
qGKmHO0dSlCLgTC4FSGheaXDgJVE4BB0YN5xBhj5Qla5UBjh/GY3OvxS7gx5mVS4
938Bi0/f80CMB63tlT+daWHeazlZmNgFjBwmpNIwkP0SZMchvyy+WkEkgHT4G3Yb
ogXD51TWf/LAS7nWXEh5k7xvHFWms1XP+pEmmyqL7ghnmMh2qgy7ttjUC5LR8kzL
EzgoM7M11Eh4OaxWjhRsgJDnJHX4XYMcmjsjzrbUUE3zZK181fbBnLIAOed48hzR
opX6UIAymHmkYNRz/SzISTuBQ8sgtAvo58DHUYEO2t+EpNIMIWTZ5p7QNY5+p8Yz
bMdc05O7Ng0DH1SsZe88Wya1W48dLeBTDzNzB+TI7jsu+E7IiNmLy4Mii0haTzbI
d0Qy0bigyko9uvYejkN4ZU7BpZwvFDaPIND8RlKsIPS7F7DBzN1Hkl4BNO4hjjX1
M+vSTZHbgujf7y4kEyGN9IbCbypV4Xty4RlVU4pVmqS0jXtDArqq4mCdu9WBKelF
GRuIjsy+l+B5UYO8M2EVz+lz8tIQ86xoGZmwqATm7Alg10aldsD24CF4TJmpq7aM
OTC4iv7nHjr45XscN5Gt2JO4Swct69ga2Ff5wHTngy+7G65AtVQ1/zpsdYoYsXqt
M6EpBWubQCbxjAADKbUZANOGb+l5n7pwfGrgh2cqx0B7+lSDX6exS5rJnxeehYDQ
ld1JIACJXJmbCf9pQ6EkfhFJJCJFl117Y/OpEPzs8ktGJLW7cpvQyarqIa0RssU7
+SdCrFrXxtmJBp3YQYMuDCxuZo5rKj2btRQLIJP0fGmncSzxCicl4lv3WoKAc8t2
7lf3NB/ovFl3m2xVpVmP/99WuNULmQE2g3k2zcs7d3C47QN2q4ko3gWE/oyPwFop
pUa3k9Z37f5aeTqfO8gWY65+5NuuY0nUlNmHOXqR0UHg+S8QwDsSBQS84xW9vNc6
4kYA2JFxipmkH0FniV1HRpeIhL+dq4LxmvgSa1VgiAz3SFayRFMG3QBQxm7s52TG
CgsQ8273heCInoLs62/2gZxo6h06R+gBkiVNp7k478awBYDijZ1MEjtan+ZSRAGY
f8N5I8It/72Km3lbvPzMl069DDMD7QG9docDUiMi9fFz+juO6HqDq9u2of8JTxda
79irclfqvWRBMB0wzPKkGmNV48dmHrilMaUzx6cMwIjzAuLGqrIS3Ei+St0/kelH
Ljs+yJXkmCxKKot0sibdEvWhv/JewfDFlHmv86Tk/ETQm17TdwHtBno95J7A7Oes
LJMA/JXNvkZLhX7lLmgXBe2CF2i1AKnlhR6OJSHXi564NszRGjBlwclZoSKsVZVk
naBObwQoQL+a4QtFwvSdY9Tx21b/u4BrvhYtxpBGNFgYTwCatbrC6111MJXE/CfC
uWQLKAYMd/ozGzeQJW8EhNP7bI5TUwWEvm4LiZ1Mx8vdUNVH/EI4d9RXV7g1Amuf
PLoEg74Nck7C4wNiSpS/kCMESoqNRl93x1Vd41mFqULsEx10aIP2LcooBIdOZu8W
Q3yN6nqSVR2Ys6c/SNBJR9sYm/Bdi+UxgGT/RI86BZMSLLnW/Y0PWBRdYW31sqKo
wkyyJfwUG519ga0GK9v50ud/PAyc8OIRFU4CMokeicUSDnVtGqU4C9zh0sdl7nbK
xTg4Jtke75MceWQMILgrpy0oU58ZnVogQFxt6VMWnK2EpEE+58ajl1lpasU5D0rJ
ITpuezWoqSDj5wPHslIG3V5OQE4+9TlBKytL6+u7zuVqaMiJs4TsXVYte2CvO3iE
FJu5AftwgE2u9Fbfm/sUcQ2AULWA1flwQ6lAQ+b7M10UI2d/u78rkdCCkjKoedgC
bkEIzQwpO/AHQLRqqsr3u6+RGUiRqmEllRXID2wQmV3C0rk/ThSh3ar3iovThPC9
dxLSua4JGjtjuKqxUAGcHKDe78pAYprK2Xy1KYaFsNqK3IxZj6RO0rlY5YIDf4sf
kemrm25srfV01Mx95IHUsp/M5EREOM0Hzoddpck8WaS6hwv2D8t8M8gTxUs8VREz
l+Hp41YBaQmumYH3+7W47D9O2jo5/HZAP+FysuxokliGdriUjvFu2y0UB2FJpWXG
pPPc3NU+BLYVAyRVBjDMJgw1TuhkCGHw6DB2xD3kR+9lm5Q+84ZHDgiaUc1W0pkw
EC+OC1/F1qkWPC0QT8RuDKOggKvnQFlzdz0XwzvMk5Ls26jpSKM7gM6on6kcmtfo
/um4okI0uB6xKtPeTIiSB1nlJr6enK6QkCK+WEHD3ONt1/4tiwea2P3rLPUGK0Yr
RvR9c53IpAO8uvUkxZwUJfjdMH/Nd0sSEr6MrRCFk+XZ68jmnwcZOENAHHMi2QxB
pZg2gcJCf4XqPdh3KFdPHvGwH1Bi6x6qAI9jPkZnHCEt1Rn6R/OfDvCzKIxpw1pA
pDRtPaBVa7SkRLVZC7f1VKQgdUx5RRHktCtJA2akuEowU5QYPlSn+X0+b35o74gI
Op50PbllS2RBkOwtTt2oLdZpNyoEfLUin6plBCfHxdsZatJas2583nNrkxlpne/U
iaVKdcC2AZiYZ2CjpUZOCAEgPA1tXKOJXgO22FIadYHrY8lEXBtvt9bEDlQYDJAz
3zuHachuL5xAnzeUP6y30JCJfQK7KKOtxSuJP1n80bmHqaLi7t7EAy7ddDCuIKMS
zwv2dXudEgJVWs+1eIQ/NH299ggQ0MbOCjv5AbdbMJLYdWHMsVhFZquIquzjv+T9
xlsUJT6Q8x7hHtwW/JfJ1ulI/aRkA3j1zmcPqMlM9sCTcWH1zNBePRw6JyraktrC
iCYJELKzjN/DBuyDioXNcx7wdkxdQFdN530Rjrq/77/pRyMcwJTW1cU9+u9Wkyuk
xe3DmdIVjrWyjAg/+LmlyzWfHDguSCqZpVeirh/sIQpbRb+4lWWCtc431oGlU1jj
1TLakOl9o4scgRWLHLKd6j0Rwcx38tF7GIbToTiJPd9ENa4CQ6+MYBhf8y4lach2
9vogFU4jZuU38HBbmmZysqnkWQZAeWn7iVemD4ofc9A+lsp5pxqDK0FVf7i8KDKr
9Qd/DQTI+AOGAMnrEhaTCccXiMXDO4TstBUynceUxtVmOP9/hFHyzV2XrZpMsrw3
z0DqL5iU0IVCciCHU6Umsk8vpts4ykZVPUc1S7CJvd7EE0jYWbTVI7R9T1aw5SQJ
bmEYHa+Yv3qqxvC+SYUZRKC8Oi6P/hlN/U5Zbdf0Qc89f1dUrrlWkPDsQKZRpfYJ
1iGhOnPs+B/rbdAj63HgEFDDZPRaxlNjLp5LEUE0oABpJPZ7Rm80zvCOiebBelCh
ZBxk0KGrigf0uDbEUPpUhLFxt4Q7Nf5EEWSWSPq2dPKXyoFT24N/4xJdCvBwr96r
9iR24YYYJtWkfOQr5GGXa+vPL4n1E6RB7uShAOOOYYXbX7dakve2+DTvjPkJMtOa
lDsKD02omp8hIKj/YHvgSgeH0lqYm+JDgmmdyALbYTLHhi522e9qTF5qAVQdnNAT
hcUhHmX6xB/dcpg5dQ7+9/UR8ETi/ExNHN0jhHYUXBw9HC78XlTr4AlRJuBw/+pY
54kdhKbyoOip50sEY9dbS8CP+4iyZb9N+6npePiJjE2KV11Vxyo8G4RX/E7Nk62Z
1mX5Q6RvNYWRXmP45LHQs6uY86w2xuvXnR3P3w+q+tzOVjfPDt+k5YU3wxfRQLsv
1Sb8IaoCaaL2HfrzRHgSlh8naNPIxw71t9GZcZe9EZc5QYHEy0GQBwXogXYDfn1C
BgaOlLk9RXIZDicBl9dHrjPu0PbIcLdxvJlA7IJsid/1rktv+xMALYePq/56nwBJ
fFGpZYv3pZvFKDHaMx6JQHkMK0J+dK7uXK+i7Zs0dZhOjC3cwaldAgc4rxO5pT1O
T7sSuO2qTOc/SRu5WsW+3whUPS5dBS51GGxwZZAOVkm4k2WRDivDx2e3Pg7GuPzh
HIeeY+J0b1zqffqikTgrqqrIDTMjSH30QHNw2Fat0GkGuog6ERcnEy4uS10su236
eCMEVp8FtqjPuOmpPi8ixKvRSUkCtS72fy5/ujLixqEGuCqoa8IKa1NIyzMTMvsW
dE8WKsn7Ze7BHFTP1/WbSVnvdAODt0CGRUZjfqz9YPgVmQb25zZlVorUE38UqJoO
8IFMJ62JkPdtkxx327CuD9rE/0FA+mSp03H5dAD5IgZe/fv8CXxrkypMYu5XF/43
RJLkjDzVI5IF/pOSFVdbPOT0GkRlGA6r+CJnEx6nf7RfoE1h05mOlQ9YCQdZnWj9
zFZaI59lkPAH0Vef1SPUfLe5HexSOPnKpYcDRk9b0pxmokPAwZvLOw5sxNwNjBRC
dNE+1wIDpHNb7OxuyVLuEFb7F/6zS6WGH8IPzHa7IHQ9BxHMxgjDm82zU2cxHQLb
EKWzbypggIj1wucO5muo/W17XmGkZW+6T66RAx+KI7W61y4nAg+XmuJQumSwruSU
2OdGzecklWRRw7OfHMPyxz60QFHqvoMTP9wmcytzZle3wGN2s8UNGsFvqjBEmPyg
vyDDCtR4tTB5q6Eg/0svrezJEbJCdFACQWHk6Wa/MAanS0SSx4vBxLeRs+PZ9/G4
Q/gDpanUM5vh5h1D3JdyAUEkDRkAVW7KxUWdIwaQwJBWKjp6aQnSMdceMc/Qgc8w
jvZh5jdYJdO64V/ZXTQhqo2YokjdQWWjy+gxEdiTjwkF3J9uSmLuFx7cBLRWGHPE
nXFv+aMLkYepXU4TJsCHw+OmfZL0VuVfwXukyOamZGI1zdy/aOPaAqUgvvviRABQ
kXGAMPVPoPXlWIsj/aKY13gHb8rgq2MLTLy31rQ5qJYb/rLj5EXz8rSTOfEZ4B8B
J3HVOa8G5oGjVKOkHfz9qUt0qZ3DIgL6avAxo1U/MzKiFuPRisE5zUWEPiVsHUMS
z+5rCpTE5hhEdX7Oc2xqSPuAfb5FWmMQa8924diHhMh7ITwVuO6jNl/hfDta+XgB
l7kboCp/n5FoD2fVsYarrWUV+DGnsrhQL6BHxCagZXy9l5a1lCDxPEDh9Pbjf+7n
Y4lJsNF5Ci2xshYgLpbqtojPh4hY96AsO6FTyVIIcvXSrRSTXSYLfley3gRovfii
h+BlXkEfcVrSo0+25vRBUcFxqenTF4omky/JZOwO5lMJI4WeVzWTpmQBtbd+aIxm
1g6JW2tCR7LKjm6vLQE6LX9mkTvKQEzt+VFumjvcX6kv4EcvSm3ykHkbNI6+hBvT
qNDpiX/XyHPrdqnls8ewj9yhvEi4kUsXFtU0bYefe7KSZBlOYHV0sm73PllI2Jtr
JpwFVaqGM+f0CgPEG44jXbgZDBlnWBIbh51QOoCtjJSvmo/kgRFQNHAF00qu9vAF
+3aRkv1mpxzYtcDCGNlFhyGFzXMe/CaHD6pKzPgUXVnf7F8dUrZ6iQhwyABFKRrK
3Ij56cXLIM1gZy8GWMOa+82kbWGEsm1NFZ1zupvHqXfAkgPPHDeYVNSuN6Oixihc
wSaaxUD+hO86CMdl8cpPJMpmpONPEhjKekIXFK6RRJ48UnhRkbdDX4LrefhXmshk
xAW8dNCrXguGjuHsUd/ACodAAX2fWN1f369ohk+c5VIcJGNVXjtMHjjTtWbPpw6Y
kuUr2VMeZ+3xp9WGro4Izc7tjTPH83/Ujhmq1u+XRqC0ctfK9xPtwoLUh0uqX/EG
xTGrg1GPdYn8l7LG5ya64k46gMVtZojhHS6xQusBLdcStrQh4yYMc69K+flzO3uk
s/bxjbXQL/Z3lPQt0Nk9KlvO1W3BAtdoW+bHz3oxUr8UAM/Uyn9tcrZAdQM3F1WJ
9oFmfqofcDdaSO5IcVNczaqxI76g9U/FONL6o6kp2djbJjIzk1aGVLFeoYpQ3I2V
XVKnGb7QL8CI6a3OkaqPr+VBof8kiV+alb0IrmKW3vVVoIYRRzK9MeAhEFMvrFQg
+R4azkjTglXqFOa7eBFagUyMlCGLAXDGuINv/VkWrC2EH7Wa8KyGqweHcHnVnJMe
JqoDiwiWAMsQzWfS5/tzC7wtleB5/5qugViLweqp92VOZg4tvWBSO4iDPfQtAfJA
mbC3CjEqYnZGqecixnXKGBQwlNOpYF0smPjAXCsTqdLFkAumTqFOOTXQ5fWNjvjO
PyxXoG7FEm57XDxhvsZzDgqanZkqaKELIZDF3lI+eiRMLhsDutfoy1OB5RTnLfyk
yuBgXjDLEMHbUv85BHSx3Rr7aZa3OHTdV01UM0HRV7s7eh2P4rHv4RMUhz8AGLkK
s/hfeejHUgiU876qIPICW43Ocz6eeBPGXASVa8cgR4invYUNETZpA2PQHRcj80v9
s1pwdWR8sZ6JyXU7wjmGBk9/ngUle+31Qyf5iVZ64b2R2YsRke6t70xBtlgxFYrm
M7dJtd0HfPyQwFKd1g6nFKZx0yqMbOr3RpH3HSvKMl7oRes4DKt295JIxiXkxqAK
jyVn12UeDe3hI9SsUeqo1kplu6FA9WaB+RMn0u77GclXCaC5kWt6GJlaMHPtqBm3
O6oltmDSz7j9MTJA4LsfQtaiHCp76qvcXGVu9Y9FlMLM867YZHGhfjP/DMP02po1
xdjr8clXBINijn5Fxp9hYGSn5IKuOk3O5Ix0GTlEMnwMkJc7y58eEoms8CInF0MV
1hktWYYUdxNgrrhjDxGiU3XXaRWhLWVycECd0tooKCGrrdNKOLHP1mVvIgQMlIjC
fkO5hyfvb5EA4Lk32HPbF1dyuv1S4VL901lFaV3nQ/C2pBNVNaUhx9NNMga5jqB3
a+hlGdHXMhRtoatoUfJJXx7QGIVzm7iNUgPlJm8PXqcQuZDYLowjqd1IVVEZLlHO
rbQ3nfF61xWwbvEv9uJjpiNW8XWrQF41iQqvRwqLpivtmEZ+ju1x1FEWi/SL7MB0
agWLsRigwIpJalN5gSoB/RMbEv2Qycfg5dTgGgm1xSQLzwNYwV3IPCaKOSz5IrjI
8dMo1qXr3o8Ji6oJyo1leKDb889No5dRq+h0d4CKLlYT2H1su4zIzUzXpb/uOIkB
RHlnx7eWtmc1nNgJhpXjHaamtxtpZ+q73QtqEJbYk+rO2GhbgBZKGPqmfxwe6gM5
0yqjEbtx4o+psY1cHxhV6+XZlLDYcr9327i3P4+PzePFRqQKyrDECRvz6h0tj0kx
FHknZrnIpCvaxkSt8PANpA6zRUxLKSrVvBeHvMMAgr+pHxYAcvS7mszF/5UOBRl6
+fh+XQCaKy8C6Mm4Ly5WQkGZIQSXMQL1cwan/5zBBodQF1Y9C8WxMtzMxaxI2sHm
OMFScVZNL3fAybxKOwBW5O1bzN0h7ApEP+zmL/EJ/u+kwKwCM0lsi7SVDsg1n8wQ
S2eu4SY36WGHm7nUH258uRY5Ht2Cb7jSxIp+66IQQcD3FbB7JnvgMRJXXChigZed
6Co7M8piJ8wdOhuEbJJY06XP0qgzoopBaID/u16EQkHUQFx8TpEZUYh2xsxxXdPy
bkS+a1DWTSHbgXPrBTM/h8Hi+drATYveRffwVvS4rgLYIowz77TCfHaBxMx57vJU
Gmm3Tq+qB5TI2+tguG/JkLhdBy+YNSRp06ip7d6S/0SjkIXdeM0NBtlobAhFAhh8
0GBeLM1BE0A+f0acuIM/uWfKR+rVKPItD+RWLKR/lXjOVfPyYW0DyGsdanE45M0Q
MLHW9nqapvAMIyjgrrUhQLgqIwglP7Djn1SLzHX1O7LFRsNKgBKTYF0lKGeB0h/U
i3MzzkZ+8R/PrmxDkAOqUjfODXTC6sj2OmyyAV3toxK9/RdRBMKNK645VlQPH1v2
GOsmConkDxmvnLOElPSQefsMKVVDTjVtD/BLNMHZSxD0FFTdY/dP8vM248d5bFhG
2BTcbSHSPdpqPgqhRSG2nBgLyQo3oeSJF8B2HJwDB+Rzsbai+UI0PdmxR2K3SQ8v
coP+bFc0nReWICC+GOoNcCxK/Ojis5s6TQ4UNrh2gZFdI0vgr7C375eylN0yMcQK
nRMXx8Ur7KjILPlVD795mxTTimn5odLsLyTiSykPoDJsM6S87BOzOzJ7QV8ddgZY
aa2syRpvsTiPmsG2sCa+nUmyP+FYPOiOK/iEFb3lahAThqX4qEvhDsxI4AYVY1Cr
Mi4cV7RFovvqcedYOIF6vjxSiGdMlTz5vQQykSFYnnNhqvXbGbsrjhDf6JUkULWt
QPon6zK1wE5B/jtFwEze3BwIRHS96pwxIY6WqCTe/raLszAih2qPf1sQ15gdafCv
9SEyHId49M7ryvDgsHPcSnMv5LdINSOv2vwfTFop43veW6yockL39iNB9o+zvkre
iwZbKSY3zhgAMggq4Oafim7BKisrN/TnVMo89fvNxVwJKnvzbeAD9rF03yMPtFBh
EeEQ3G+C6tAgYP8Y1YnQwB+CcGkVKZ9fTb0j3NoERCA9OC55MSd3KN/kTsO2SVGQ
anymFMR+De31eMyKgOOg1FtpCjkZ+LV+YXAB7sqTnhGB+75TtM5xTlI7KryFPpeF
RA2KD10F5TYENx7bWLO6+fLBaAkTclldFYYNhLfs5/wQ5uk5sFnvLyM/FAOO7+Vj
WHot2+cXrQ74MZ8ve6fs0NbRlMtExF7AEJqueb4fGUVT8ydHIvexcUp1471vRAeQ
G/xI8MOvw1lI3yAL48/mo59fqFPL+CCfXPGOSQXjQ+X8ueQQ08DdXr88Sz8HBWJZ
7QteTEOa1hqCG6UaKAwzxR9q3Kws/HvAE1dC09zIYAHQN3C5EKtWWarzYAeCQcJu
FoxWGRgn6q1Q2eT+2PgiMDgXEoMPfrjVoFYpH5sE6fiiarOcZM6kVeHyMBu7HYMf
4JIN7bXVt0BdnCpTVLqE9crFG0F90h+u2t3wkYZMWSsXxJgdtOzY8DPObJU1wLWy
gakvkdGFaXDhVoTuqYGIy82rU1khFQ1KVNL8DRHvl9q9eu6zFa9P6GigIFRKFNn6
MZN/qZUl0+JUOuTKFS2oL4QR28YTWMuDu3yzR28BBVIRgcxRhJsFtnpbufoHgBVg
umPhr1UpJknoiazRegb+xpIB71+nRUqv1Gkc8emkvB5hj8bRxq2GbKo9Tpmm5bJ9
i8P+Kgsa8Vs8a7ExdJi7yyLTYxnEJ+5vpXwYTWM/OUafqJravj9CJlhfqwXPjINn
wzO66XhyjcrLnVY+qCIWIzQ1uN/qjinfEdE0evkgEK6sIRjk+tS9E75mkjK9AxHe
RfSe9cu8wGduKxwLsdWBo8amv4u6V7zyKkPCvF2AV4H73tRx2oHa2qB1ASMq+fdc
ZF28a9blHdtChkgnaO1HL/oA3XIcOMaeMfeA37Hw/BStf1+3oOjw+jUY/2/vysQn
u7/zekVizVDTVC9QPbPr93UpCBtlXmVwCgY02j0X9CL/vHS2EIHyqtMXAA6HWn1P
GD7HeDPvsreaPg4rUH/DIBSw34zxaebbjzYQ7fPnTl23zZTd3/Gba+VqwVNgMhDS
Ms+R1ugmcEreara8mjm2jLlKirZTkC2bm/YWRQexOf4hC56o0Bsiq24oVEslmOYM
kzwP9zDdo+B6/KfoRxdNjrhWSCEMQruCx4GFlRAIMdx6b81trWY0A25mHf6j8QxT
LKZ1m7uk5U/rFZR9T6fy9R9uxwCm/S3R4p7reZU5iToa9CPSZHOYBs5KalaIFlQr
ID03VQ4J3AJEhOGuF3HMfcxk0VyncRT0oKPqRbUv1E4e+XaS6lArHP3QWd31cfnw
C4lpAFYsPNMeU2xBIkn4tCi+TQU9RN04cTvN9DgytuIoOH7H2JD6BjLnFXbcvR8n
9+yMDCQKz87HCUq+BIvpGh9ykRB9GNumO0/KKvSaf2ckd5x4Ixt49pQ4TPphlmmG
Rt/c/WiQrT75wlQSeEb4eIlbB1OMsBHlIhqnYfansQldEywbZxO5SFVtMsDTEiqR
lQ4Ugd33w7uKJkQrjXJJwIZvi4gb8uK69UQzQ63KPfbCrj2sJowgy8GuL0rnD8tG
TY+ogooIeNyuYlL444Fxc8NeaceHFRjZzAKXZQaf+liSohnNin3CZ+Hm4eIzQKXT
0I+jgL3xW4DoHTXq8ouu6+UCxx0CKSY0csttNNdq5TwU8R2mnpWpWaWPFxtig2op
evSuuq+vacDehyiuUf30DHxhdPRoN49cBp5O9czVCeX6BzfoBG3uk0EilfLhPi5R
7XjPnoNLJbcwwOYtX3OddFRUWZxUPWHvhQNRUuJNnodImxIXkMjnR4FCx4XgVbjW
oXc4IkWuBf+NLZ4F/5zcJq4+qHh67kLYPiH0oGOXsxm1o+qvMj/HhEM0sioPQa4r
HMZuXiYV5x41J+443JTLuWXALgQU1KRvMrmkJb0OIlLDrDrJhzgl48ROR2wTDGli
ORJy1yi55stAGT1tWDO7WF8OKQcUm3yZLCrTsX6ciY3rI9ttwgddJh7/pPZF5sjm
Ip17beF/29JB4qlMGw/NqXnURZzvrfXQZgUHJ5p1a/RNdR/hy4IdwL6lgjh793VP
0GW/VUJXE+Q0Z5dYczmbdrfEUFenVTsUqP/fP6VFBrsOghbA3PIGnhYRReguNokt
11eTNVSvyh/OKsCrY1LR5Akuc7pXtWlQGdfb4ooKcis+T8UFJltZ7m2TfyDV0tOI
AD0l9q8wkR0XziOAU/d6VPKmiKPikUbBQ7bjhJn+79Ahwd/6jYmnI2BLOPJCvNvt
X0s/5SirIKJGIaAXglNJAQDj4RGN1g1wnKeeS/un1puK3alQIZ5J9ySmhu/8UKMy
dJzCwYjgqIWLAXp7uEaKqYt6PkI8BV+Qm3K8Fh/0dFtLt2XTcUuw2HXQXafgZsYe
eDrCpMnJrrEV/+ZCvT+EHBiorpQvrZv85b3D/LO/77Te7n2lFpgMJaCa/Qf3xzwf
Skh6qVaL5NH6vTvwSSMhxDcyPZylH84xyLPP+lYqiDztAp9AKSuQ/D/ecZhR6Gkn
rAuAQu3TaUxBzsYHLMobrdgzhXTx8rta/c6aHVbfw2Vny6uQHPZR7/uhJCL4JzKh
KUOGHKnYWJPzOmIExOODoK3Y+byhanhzrPn5FPoFe8Rfgx41ESozivx2nSwNPByj
tyQAXKyO4dpuerx68KAiDP1ENYrPvfxPYbanok2g8O5otwJsBaxEZEmIa5jqsL2r
okKt61lsoSobHrIw3PcF75HyN9cDW49ebvF4+t3dlaH06Vf4P8ZamBewQrT8Vz2G
FT12CmutsI/K2OLPaDnvf07+GaRDAhWbPOXL+epbp/1Tls9LvjVsGVM8e2G5oTQP
19wRcCEppxlHpEE6vjz6QwRkIiqI8A03aGg/ZKel1cKPnc0UPMMnd+fD8TJsWg8l
8/GtibLsR9Y9sCbEy4NBMv3+Sy8jmf3o3K0kh4sbhajYYEhKNTlj6X6J/JgkdUF0
Z3EekD0w0KI5gFPYHO/3ujVkg7woYZD+GszL7OYYj+2QFS52wvfcBF6GafOiiXJx
OOPPtSWnVMCPEGCqpszGArNsbi4VmjK5a2bf42tKOiJZOP/5Y5pQjDSrqyNTgszj
xkjkDhHCCKDDlUV2+53oZ+dEyhiggs4DHBff1QCxyUnG7pTXsb2AJwNI7ClIWzxR
8dBT3l5D2v96P0LxC/2Z//E/v6boMPfseETamJKE8lDUWcJ7rCPHD12l1WJlaq/3
vPJYQ/uqDSOaE3TfwlQJ0joGqcTGTkfAW1yOrpQkNZLFBZh3UV+otcmQNd461MFU
PwXPzuN4wOxtbGFQ41B0/eE2HQeUf+vGSuzqKMcmCmTgCTXNNw+cGXFsTc8zt2cR
yBFHIjhQKZeuN9Tw3UGNvGiYpc+ryj5tO3cv+mgK6myDxtiaRKymt48zE+9KXXUt
bp++s/m63n4mVtMV+ZlibAMkjFWycFseW08aXDAbASdwDv5asZgA6AWdKaiWJ9ig
dYEvNj7x7W6MgATxLXT7QOOr1U98BKlNtxR0dZfMUInuU8MwOERydLRQvFtlKgkM
gcLayyuxB8WO8kXrbWcTcpVywZ507pNUZIZkwRzk7Kx+U4IgPdCkxfWyTxtchDQL
Nf0BQYt/2QVEOyoR9TzvdDLsm+3QhqCskzwjE9geSrkLJDwY/Wd2Bh32UrAWg6Zg
g+XHaYIL79Z8XwOBOZyzO/wdZbmYEA36klSHZa9comjjnja/pAk+/AwEVBWj0UVi
6mL+y86ixBYCIrSIuyL27Cb3l8p9zsNAG6SbJmGexZhU6lKs2/4k2E7q9pku6cmZ
qDrjcoBdOwGUFpyM6RBWSBuLMalzeV+HQSBcmDbTY4xO/xNxBgRZv7Gj+P5z+11k
U6tDFGk9eLQmPaEZlt4+g/BFbhjf39BX+gll/cECGZEEzk9F/vEOL2Bt2VHIh7Jj
feWVASVjQqectqOxsGClSSoJSAQFt98q3Oi1PO2gaityXWL2yRXwG1Ty1VSiI4ZJ
OzRNB1EbOZuadASkPSZXMVOO5jr7HACGr+0/oLRjs0o5n/r7h9drl9UtOOF7WgOa
+wy2prBubUNtcjfwvzezb/BKOEF2PZbrAqxMewLtBEiB1Yiq0oQz9LgOySpA0Hjk
kgz843Jl0DWzbC4GS2DgE28mjgDKNa15lRXHHDOF+l4UCc4O4Tbi10inBE6F5B5g
DLryyXQDyGQLUv96NMtV/ePVM9OJI64O6IuyoczX4H5mfLJC8hYCJ3x0zv9ubSYL
vlqpcWLp7WDrUjrwtU7TWHRcZTfsgh85R4lKlGjwk2Tkm8ynW+Uu9XvtCDHhorfK
t97lQ6+uOPujboKaSMEaVwoRVelXV3/HL6Ut5smHuavcbLW1MgMKHZtSvLl/XrcG
vRlkxQ5t0A8bzEL05FGgvut8pkV+U8l/f5MWtQzqVUXvXz0fmWV5rKrFwtayQ2Q4
EmGgnSf73cu/Bas/bUg8lPbng/tTWoQBLaln77RzSSE8A8NiUsING0URNI7ndN/e
CaNsNWEdZnnfCYaMFpK5bQ4H8FtICg8WMYwM8VgMrMqY/tA6KXKQnvGxqlZP5gRA
meuVwI80KkvO/JeGfQdq2xCX5+FFli9GvXVtcsgA8m48v+9FOrJJ+OM/40OqRrSO
69KUgMtSMrW9+xgttpaojk4V8Iv3knZS7AHEIDWyrORKa3xNPitOr4GZSe8a8oR2
OcmaaLs9A1zdjbC2fkoiQ5r6km5+q+UfPYmqBh2czXv1/1zRak1cdx+cFRIvYAkK
98CWnkO76Z5K06KfEuOivoTtGhDsHdz4vFq0oDMj+Ow9z17juwmUdT0cDflL6GQa
i1DsDX85YkipUKiY4mcn12o71mwpd8Vsyp6Md3SsL3nzDK9KCr18Prb/Xkhv3mbM
ah0Tz2IvY1lWoFbKNaXGRVBuswstUv96ViZ4cc/imfAgn9GT3yb1UIoG16cyXG6V
3NF/P1VywaMqGT9GFVk53voy0YbWOKVZkrSU/5g7oTCamwlKSfkvEuDf4NFEqKiG
Myx7gAOKJI65feObz0V2ywF0TeH2dO+3JPQM9Dtl6mhT3K6cIaUmQ6l33yfBzsb2
LCjbOEoUYlqdTGC73R0qGt/GZ0WVmK1V+XExjbQJnCitS9S8rebUetTa+kgJ0zt0
bykMzbAGr+UxtrFNvE6pSwgIZEPHIeDtLQEg0Oyqv9l2Jpsr/FkwpCb3kWPNf2i5
LaEseZqNUrJ6M9zDGwfuCKvq33LkwSQNOcPRC6TcZYiLp2jimkyKszG3888VWBb5
ZYR3PsbeqnkZ36ndgCfr+BFhhY7RnxnulRyrGTNWLzy6Z9YW/EmZlFm6MQV5qKVu
h/VsVbbSnmR/8K18efSQGsQ+Lh8zuTtCHQL539L6OkZ7Bj+9H6C6CGrzlsGHNMA5
5Q+Wn3A0l2lNIKwQtlRXsjaMl7ucNtOiJrff/wH1VO/dr0YWQE09Ywprr6nb/dZ5
ddReps+6vVo//kX70IKyduhsyJR37ZWmla50yrmwH7e2BuPPkUlSyolhu21ebK9k
o7OflHV56f8ipN9MncGFI/UhAG6gTFBLssLmpejItHHfArioEUpwyTV5+sdIk5lW
4w3LHw+HBAO0xExQaex8oR9y3mXao8uV2gmpuSPeGov8LHfxe1M5D9TefV7TIght
bbmT0jQ5p/amwqRMHKIlO+CmmZWATBa5QIBwDr5i58fpmirBpAzeeLfAmk3IdsOq
GHZ9BrAD03/kNx7ympFEJm08t4vBGOALxvnwfV9yjI7NoFw2yrOPj4TpukhOWRxW
0RJpsw7LCNLMk9uR0HgYCoeJKxI66/NWy1mUQ1MxGJ6vDOrKrmON7EGFX2k0nH6I
gTu9ddA9+phCwS8soLP7Ya54bn0Cs3joNHFoGuYmxaBUSEtGGwVzYyIRkFJyDe+1
iADVbYJBv2kclmh3GmxpFqS/HkfJOCmE71RevP5yvFZAnjaIBBRH4MzWMlYmOdW3
wvvPGmgKWkIKDYPk2NzPW3Vf9DPfTCD2mqmfGGES2m1Mxl1dbtnDSrm29gtDCFhl
ji0eruQ6wlJFB0AFMsx02kVqjFjpVq1Lleciv2IwPeoYRqSydT6pN0kfRTwP7OSc
ZKBi6/9rsVJgp3LNxN2RdaDKnb8jud1KqGyH+MCLNQtx+pro5UyRZqHURW8ZPIRb
znUO4UIWSd+fh+Ig/4L7lZsWuDxeZN/wrj1BIJKZsxu1yG3G+DAKDiqd4kKRo36R
iTE4NwRXqEGT0XvYUq3qAv22YSznBkpwuHCaVvr1lHqsC5TmPol6hr5NQa+J8ozF
q+Mattq+nS/MOgm+VKWK4ShW532R2ZlPghEgWhP8Fh4b3/US5nnMOLxmMiMJssRD
h2Hw3eabC3HtgnQ0Yh0Z0VmC6m8mmRzTcncHoUGSMi7v3yS3/fTq6I3Sj2YdECM3
xOYJyN46vT8sgkwju+odr5lEOSQOfb5HSOq/0YJa17cnGBtDTW3s9r/5b5z0RBC2
wODfTdOEF0afIPrlbfkrFWtryCHugVdASuyt/PoRzyj5SAAFQt5bufpSpBswmL8L
lK4O1JiMR3/70jQab3m3EzvpJXBZPhuWRMlqsNiWXddMRpjlw5zBvSRzY+2gllW6
zr3ZlKm4vLRGTZDcIq1IZ4Q+ncjyz7eXNzn2q4iSFJ+03Bz/2VqkXXVW79s8MvM2
ui46l3WzwkLSoMPxXmFf+XjusXwEvuMb6kKVw+8j54xiL1bF7q7kUbHrU6/QTieX
cV4kU0apF5Mt7N1NxRtddJ79FThgkbsszvvZBaOLGKDCCvnYfVWBWF+HRroh6a5f
iYQnUVlXE3GdT/ZCqh7r52gnLGR51ECByvJNCn/L1Xg+JJNZ+QHmnW/IvjUSRNs1
lIiMplF+cjB+uSlkZFLIvSidFe8XWao1m3dSPcPvs0tLFKUDnI1y4oraO/oLtoKu
eD/QaVUL8KNqTQ4NiXxgzXZ4unYG5Ha8FD1lsKhm+aqx1Ef0HTsXKohAaROUt7jz
tHWDc+hdwulCJt593P7dZXHculeaIF9yH3zCtEd/+j7NvTlUjIMgttnVYSFxfrul
GDfYkStdCLirfl13LstfLQGtU0JpFLV8iYDu/EKRUcq5TQe3HLWZeZToT6gXETqr
NIRcd/MoHaJ3SSJRZCIpQT8/IcB7ZbiQLOkzCNz3LFdvz6lVNLfVSwg7oXKLLBTd
UCuX38NAtGFSkOSlM3HsIU5IAvC+tieFFlDEBMNzxQdstcIFEZEQ+T17pVocWR3I
BNoyQXKZIxB7gx+HASJ2x6uiYkxpDq6Mdd7hIdpgMoxopDuH3xoiSzk4vlp1nqU3
0USChX6DKRI+IHfOnN3KdNO2rnyMkO56CAkddOv3U//fpuhqaB8KdmrgaFxLZXm8
zpoqpPXKn0GzaICewZQH+7KjEG0wnuzh1AhDlKdQOu3lGCCNh1G19nR0zg8Q+eiS
Xv1sKB7/1Ojcpoe/dx4zd1iq4kAukZIAG/ozIW2EWMiNWVXnq0F+EKxv2u1Ife2I
RRuABBXPgVlBWAPgBaApRZlyR5upiTF3IJu2Zywm/OTGoTR0/Xa1jJga88KHLwrR
TWIGBy44mkP8SNZeBxxIxNPU/SQm31Bh7yiR8F7XryPBqs2aLodpolRYn9cNrabp
SethwhL1Btr9bPsmeqzBlTzuhGcw4UcTbWBhZxwPB1LwMhEMwmm+Uj77e7DzE0i7
aJv13mXmyUGr65NZ12e/VtEQ0L8rlJd38No33n8CdGmgMyvZ/F0GgAYObK1zlrUq
kQIWt9uU+g42B1j83ymvtUBwOZwhbMIVEwo3jKz5SMhp3101VA7G0dFxHcsc/jOk
gGV+axACzXKIKPUNlT6+uj0sDG0gtpp3zI/x0tSbsyCyxV9e39EFD0umnyIZK92f
Fbv1xKSfOCYFzxxXlyfi916BcwPeXEmSqhIQg9h6S0ie1Cz1EXV/2lvN+B9TQs4l
KHxLjJqs9tX4Tvprvmhder2D2cOpSi6dDmxp3cx7/0qh2dIOd5l9U2txgpWpYqsy
2NDMMG9SF+Bt97dNfwOiybRrg+kkPUuyHL1e+HPhIczR04uRzB28N2EMwOqkfbY+
e69wyy89AExErrlpWpi4antBR4A0SKJH0OX8+FB3VweqMECnn5PODctZYYm7ovr8
EHHuujb8oZ+LWbmVo+VAWzGHxdW6vUB9WtCaMvMovZVLUJ7VFt8ILdLoiVQ/Tk3V
G/aeILnNBAcyC7a+xNzv8jqfPqcsrU/KtXvj+cCRkAmgPbS1/kZXITxvVeonSRyJ
BgO82H0HYZ9mJIeN6froYj4L3IOXmRFceWKypSkwwCklwzRKTmMnKeKuWEyCIEnR
FAT52lTA1wnBllE8TXsKFrJO4fSKAHl94jRxf5hEv3qIo+SqgLJ1a8e3cvN45YMP
xGuaS43YGbFeeXDfZeIX7/Y0UmqGRzgeoT5y+lWNXcU5ziTHGZXcNN6kI7x7GwX9
cPpSK2qwcedtObxJ44jEWFOzwjGLbzxMt1PacZhUZoHHQOGwIAV1MdAJwmQKMZZN
gXSWcXCyClMStVz4NUUds5IHxUbP4Hray1975dUCug+xyE1OOR3wxzVjqB/NimlY
qZALscjPs8PugSKsUnS0EQI+reo4gp0/RFzF4nOE9ngvxh7LCeSUReVyz1WAYR7r
cLQAsVfkM2AAe1rQJ+iT7PCqaeo0KzRZrNTETjAoG0l401kYlSewdeM5nq8c9DWp
zuLXlcKWcERjBKu/Aebq1JCVWRLMvyCx+8zgk+zujh2ogS81Wnm2YdNiQdNiwrq6
MHq8DD3LZae+Jh/JPBr9fccCl03o3RhTTt2TwCtsbn/j0dQDMS8gX5//vdQOPBUG
Nmt0N0rNz2h5hDfiGY3ySofpQNxzYntyLYnH2l40e4B+K20D1+zZ6ot2Vvu4NiP7
NJw83rLrxu/yScA0jCjo1k6mYqBHvSvpK6AahjT8KvanvtBqKlWU/lfOAQN7paVc
YsXau7A1DDVW7yFbGDZfQU0F56g3nhosnepeAgf0TDBKBYxOVOST92gODJmxK/r4
ucJ9vhzDabsApW5MOfTPLPjbhJYx19diOX3WlJFbengmSnavNIgYbCAzJP2o+ywi
uUeRTSTYOTOnvhcStc+NznfjJi2t823UnJk7skkACXNxamPGkHmB6HOHI2gvuhF3
YV+Z7l+GJ9FBN+/C3wNTu9HimsIs5X5NE0uW2/eMb4EYPIIx68hK21zwyLXj83si
VAtwbkL2AzK5LLA5DN0o77UJAql6tIkSTaxogLRTkaJDfo5EEIueC4mmTm94TnrL
zaE13zTWqs/afFXrgpOzunnh1PivA59ZA9mfD97zSY++TBR/Tw4v732Zo7yMrOdR
nP6qW/HcibHBKBgNG9OzNAu1G+EOE7NGig5PH6Gn81MQPpIoUyGmrTnW6/byBUNQ
7e4qHu0SxPY1mESpwC1cVSHVwjUSQIBKC6Hdh/GUOHx+xfLD6sKJBa5Z8w6aHGpH
ZvqlWuvyNUAD3pFnKo2vrMLvpDYGoiZzYr1y7Kng8EgYtLIybQbtnncsU7flWetj
K/1SO28xnqgqs+8dpzSp0XmdYhhejRAlB5GJG2XNYQvivehsbNsdMf/kwBl7v8Vu
O6e56BuDeQ+zcDYLT4KqtqBwmLOQYoYl3ehh0a4zcyQIVtrQgUMxdNqzjOSqLwbZ
ABcGhSq4bJmJ5URKIiDC/aNht68IKkMOqXoXO+yfCKARSCkogHqZMz2lcGx3oFmn
s/Wenz88tZY8Vq1Tt3gMW7MzmOqzvxYxkbOHHzvOj2ULL2vnSRHboDaK25NcS6KU
he8Qg7FJ6mkXpuVpH78j7C2WY/gRFiucEwVDvtpiYNqjDXhfb/0R+NbHbdcn3L+O
mrleICwPWxeaomhHEMVwRvvEyRaa6oFeX+QqSv4oroR7ZreJOCkupsu6Apc0o8ZJ
/jf3+qkq9jHilEJgaz5ONJLWe/TmRwtybWfRAOk1ubLxd8etKl/Q9YpJwTv3a0BZ
ed5H3WC4CbgVs3HtMp9zK2Uw7AvkQqqkTzh22AtSwAgVc0nduAOxmcwg2MhaI+A+
iWXIEy7IdzWf3dSs6Y+7xCARodeq236yKM00QVAlygPGjx7EJtJE4W3jkjBU0PGi
w4mg1SZvgU3SqmgoB67Y1ViExeUV1XXwKocV8iZ5SYwXPT+Ha8EuLuL/5YNG4OqB
xjGP2honbXkozeE3feo1VhPEHXnA8WUQ3Q+KfPo6XkqcA1zLlogV/DTu6WXHZFPY
CfzWWAmgZ+xhX6qujpOp+7kBD/2wkLuU8OHe7WtfwN32u7f07tC3fK8FabLS2PI2
4Ep9b8F1DExw5D4GCrwxQlcPX/QBnJU7uTHWtwRwqegxLsJToX3vNDnW3XZExPIa
SKwrj77+0BOdG4iEddMJZgjqz+QapVloJo0pX7t220tCH/Farwl2Yj+LewAuqcZu
0Ys5Wvtmspo2wUCwVlcO5tRmAiw2e01+bb9oB9jwJ1cSfk0mPSAplU2+ygo0/g68
PEVogHlCap0CAs01ErHVnKLckCj29jTSEpBzajFQr2HZWhUy0OMqZFZqgVH5iodv
Q2MVRr6RLfVXaHQS/56VSUQ0jUMQXVCEwJYv5m0Nw2c2EBYGmMdOLpTZs0U7rV6B
mkZ3boQAoiw+atjwMFtASXDPydRFCszQ+Y8IZMwK1tUAc+N/q7mhiiL8tXKolmPI
VqA5d5mWWUSfmxOjewdGh4oHw/kor6fVxUviOhiGWA2t0PKp++A5tz/eae/xsAub
2V2lebRYgHWVkLqveW56gPdzxyaPcsSSra1PVb8fT/aho4kPfrHQEoOEq5qK+oEf
6DeuSLSmEm4wuLTEPzpLiVbNUXKBo6Cjy65yPNQA9TFQgmgnIZPSVW9gxfbyjqic
gTFpr0XeeZmECGM2YJ/DDneekffQ94gl6WAt/ak7ZgngfirOP71FvsG1rQk7t3zM
wXHkgM3Gv7DrVWnkqF1TPZk1L/VeuQbaHybzUJasSHoqPs/+Y312C/Edu2CP1i1W
sbIRaxQ34AVxsPy7+SZoHdLmL8PFZqVYJejrfUZQkbXbsZiQ6uP2yMcPjNt1QxAN
HFQKZey58RyG3razXwjh5/htxmE9ty9u08VXbHq/SNNJeHBNU+X0OEX2AFhzQcQx
/Is8ewOwbZtDhwhhr3XFjhAciFMCDCcJ3pt7SGFtpBNGNT/v+W2FIX1T56Hgcemm
iarHF9/8FZie9N7qZCoSf2FXhD15apnybNDZDZVrvPmCkK4dDgsI977Z1M/O+0cD
u+QyrpeUPu+I46vo8A7sS4Yl96RsS3JUURnO5IDFtmMvrHEkv7AWP4bxhghm4rtn
b06YpORmDiGMpChwY53YjdJ0ooRUoKoX0wD1Pt3w/PMBifCMpujANc5DCZuyCQa5
nEt12xHYFRbok1Aa+TO5C9EBuyjbBjV9lWbdMd2uJt5QP2wNBXQNpDJ55R12oFik
ZxFLWrJ1vyx2s/Kt9L8KfNtFjk0jEuZArNjqEpigKSMmael80QG1/cq4XAT84y0n
lTFzuKhIq3L0c0kcnVsug8lJpjdnkqUDvkgM40pGWyAR+5BVQ8sTz7qQ7tS1lTFM
BhG7d9HCZ+rLVlvaog0NcFTAmLiLFuZrdn5wgEhsvztfsqHxIAlsRXZkgnWUChH1
auxqpfskDPx3UfVY1H7hw9nzYTF3gcmTqW5fg0HuOlUhZ4KeUQUoNtENnKvTkSPy
qjSSp3cv9L4jS2nxEouXt2S4Lg0GAD1lAZnweHfL/TD8RTBSZOdi7B6eMz6IYJPb
ToasApWNuEETT4KQbdTcUSk77mQTbmHi7RqMeMRhRpQ+IdH1WQmwcW6QEyn2NyTU
fx5mg4xL1SGz04N21Pf/hzTI0qBdYkykZEblLr5U6DXgG2iYWrYpmV7qNiJyy8We
xlP1ZzKnrHneW9JKjaTW3i9j5cCFgkDjwIdk1lrMJ/ISPPTIc4rw2k1OIrQM0mxj
iqQp5Yww/S1V6fNu6z4OyaZExhPvctoYAW0YDZPwHPikHYW5PGIhLbwI4RVRu7DT
YzEg5pzsoELKmnYMOBpbD114dCjR1s+9s57uNr5w24C5Y0KjqAQwjzomFTTMHwvH
0olckVCcDTlUKvLphvxKYSSDznAwyoLswSD5vsSNEj9GKAQyGWDa4ArpGWSF4eRA
vb0QgVpgW2dOT7/Our0G9BUjT0k1WFZp0vnLEZ0MT5ZyjzZbEbZmlsWou1tfgbDs
7IrUr37JAbImtnhumIy1tppvJgwYCayC1LO/aJ2vTs5TH/C3rO06UHpLs2wo7BCj
FcEN8rmqY8WRQrsopv3SoZ7GlUEZl1PS8UpJ71culbGTxpJeu/6h3rpfHIDbPo/E
eH/Uv7rQWc4t5wK+zV9GA/FO17Q4yRFiwsorwKpK/g0cWLyzzqZol17rOLkZALjf
kyBot44lx5RV/tHyOSmr6J26YmO0aitnKkNggVCiyJbIE6u+y104r1nmHRM13MqF
cVBHTUOH77WkcDHpUGb/zNtQq6TkgsGKZwwwfCGNYmDd3zH9fYHTOnq0vzkgd0mi
mwlDyDrUVliKUpMit50LbY89pTR7wbid3g3vC41LdCom/a4/s8/R094sv0BoGhVr
twwcljrffLGKhe8qzib2Ug+mTXJvANMe7UhpxGRek4tR1b9CQL2v2AYSsycxDPnM
cjlwV8izF+8nwrhkYWFtbEShvjeAcgsx9RiYZJ8ZVex+4VOifkR3IwrZTwws37Tn
PhN05CM+xYO7FvXmFR4utS47ntPnXaI04SkrV1D1GbUQg5wOjZFcKYCACDerzgBz
hANyOZmhOp4q74/aT2FkX6+yg5+27pVB92aElbcmHYD9e6gqZ7DZE1qzST/iW1RC
hpMrDoUaTnGcYYxGn5ziQN4v3OdeJixjG2OtEcaOLvozKGhFewRuIpoHucmIL2gx
uQpHZKIGq8LwyMaKo96glbk+PC7PoGU4K4gx9Ej426LRsEdw9MbsjW6I5ZtlUXwk
RT0cdgtygVVZAgfleZgXpdLIKLoPKW11PjQ3+R72xNGKkJ/fWzb4T+QeKQMq8+3C
SnhTZV75hOBMm0n1s9Fwh6hRbkmMZbzXGzQSDua/44X7UnbmhSPAL1px8Hpe8Xnx
0F/reA5BqUl6JuA+uSlI0Kf3F4mwg/UCVf6PVpxGPzr13TYskK/BUYa9fbdFZTIy
adNFcOz4drdwT33Mgcm2DPk7AMGGjmR24XOZXIRXuh9zHhHBuNfcuXmt7qaXvG1Y
FJ6VeSkvM2F/V2K1+fzAuMkGbY9Hphhle1UlHx6BTjrVXNCP2kYOUvHfhiNAfXyO
xF5I76asklIRqUMkZ6jgdJFtE4tHIFObnqty0TAL95HS95O3AwRC0ezIf+D5fEmH
HIyCzOZZn2pW3gLwkGgGi3h5ybhMK8wWeQlNPhNF8smOs6W+I6jm/o0LiyWONQaA
EeSOYBeX+Ac0/u7IAbFA2HKKuWr5nQpMnGUnBUSvFjMD5HLPDRACkLaZCoQWsuER
Et8jfuc/4oCvVtCvJbbEJAEtDTI1/p2SYdwFBbuh5VRTmzEWkB+t7Eaxm3rZ63aF
KDtsTBk9J+dFfj/45DqKoLFnXTjgRXxxraLCsHjF/WJAR0/GlPUepRWVhjl5xbfM
oSlDE6k5XyZm7YPx3TPEu5jDWh2UQgOLzngxL2V5rFh4gKdZtX0KyHauqfqGv+uA
lXayYcAn0d+R0dC0lo6BA1o7uVT4F3qqVs466z1MUdhn1pmIOJa8FFsyT/evvxth
nIW4aSLtiHqtNE05k6P7W2MsIyzzIjvKoGhfiDROTrCucVCGN/Sr2kwa67j5NFuC
CR3pV+BiQdvgDDPw62BfJTALfxtM4CL+ACyiuGaHBUAjb346Xode+I3gGCxo0sVm
oZwFtPzNncjKHJnCc0x06fSIksTDYTudlFtAECgKpKeRQUCLxvYi+9Zxos/jWLP0
9dX3QJ/o9YkMS9DxsoL5BCvSdgcSvcgcQPlmYEM3LoUozseczOYTtNR1s8SVzQOa
QGYKqKsbjHKjV3c4DcrgME4ce9KnqiU48JR+9ngQW9nEV/BfMdWNcl5YHQiIdGcu
Rb/mHDlNZQ+kHbflicHLL7qMx8RFCzCGyAfVzbOyo2xVXVoJdpkWvLUcg5e7wvtr
rYUvEtiQTTD7dlL/169VpGYasOsPPBVG635sVHYx6fOtCSjWJUC7jx0+70z1X+dB
EtPWj4f93MYTUSODiVHs9acdUTli9O2yeScd9hNiVK5AT+mDapuGBH6+eGq0V8G8
bjGwlxodPM+2pAeV9a7CfRIprlQY1EmB2AmJuygwAU1vxh349Pv1KY5IxEGQpXd4
mO+1fCD9NbMnY5G1JsudliHu/efHjrUSGlCtnU+sxVVkk9FoSSYl3kycmHiRL0lY
qG+Bb1CxU8lSubSL/vTWYvYMa/0glXEqfgII0WL4lwKoJJ9Q0dV+zNvegC55nhuh
Ldd1YXQFWzg1+YtYFdE4uGywTkukpMQYcgRyrc8LKNYDqfdx9Z6bWtQ0ZS11BYDk
KdMbBKTKqL1A0FAm/O66PVa1kQTxOtjTjA0oAu+yb431MkKiEJ3ltBEiSiEa/QO4
1y4BE/QEuV6JXWCxGUUjIZZHSssI9XhhvCatDIsZT0WcjgcDlEdzeqKMLr8uEuo/
B5jN81AAMlfal0fu0w//bgSxfqfoZD5y3pyPxjCHaqwKN6enCTSGeKoX535Foqsg
j5Gw2THOr6hWrbRDMfFmMgu2EcCwwj4ssTg8HHAilhxsg2JrWXHmdGCGQQiNdTVi
SFqArKirqd2yQwz7YRIQ4jN3VB0GhLGw4/doN7IUlSGOlYdeazs3uNDwpIzsr34z
XYxRg49N0QYLrPv1S/dFT0jqnrSO6cKhGn+ENT0hAgO+cKQyssSlhsDpG4JJtFBk
HC7xlQ8DL00RWiC+kydZTYBwNQ3+mtJBgqyJLBchYoawNe1rOfBxHuI3p8RvWhO3
9QCgGYau1lP4k0K2Rn3DgAroa5+tBJYP969GN5i1GfCwcy5LRViWSCXcdF+DYWyM
7zFKeRXzRmRRUHXUzoZCGmwGO9fzlUDZHkERm5n1s3i6+FLk6nLGQyIGi5HlqlmM
6xxLJAhhk46YyI2my7mKJqtGo7PYX/1/AukXDsWrH+HUsFuZP6pGVQeQVq+GOiLq
S9IqQmEkwzmqDPEORVaqfDJHlzUKA+Zu76nrfuDXzE4RVbk3tmx1qE3l+zJ+HKhz
AVL2TrHht4YcGsVCOot7YlF49HSOKseLoA9ZRp/2BZOjTxKIJcPuWw/wpXMO94rq
75pTwTJOEoYp/w4Y5VIsoC0jmPHRBKXbJaSnzA/ED3AWL/UufH4ZWiHz55wlL9pB
hQXI5zx1He7EKOmsDPzUJekTZ8S8j+agVWshlVUKqHgv8EGDPY03GKf3MAolL6Rq
tVpMkNl4HR/NSmDVg9Y3KWY6X56clXipTuE4JP8DfGwOSmWfGh3QWPt9izlo+/sg
9ZjGSt8ZHzql7i2llL6AmteDJHue9DDO1rxRmvNhZaGARuP3Cw5kYn96ovvHus30
EVeG2RXykYl2u6x/1zBN9iQnd69dmEI+8V/I357Ct8d/zg3Ke9/PDrYu9Chcf8Fg
xWIuRc+CTWM9yWMqJSqjJktslYMHp2VEhqg+PagjU6L8Bg0vKRS313FaXOK0VzI5
UrJJvO8sUgrZI0a0T5iAPH39mUv7Z5aqV/UERpA41c06lYZhHe0pMWwp2jogxMof
sGLpWdqJQ5txD7VNSF73K6JZFgU7mG8H+7wMmBC0Z9gsQwvvwWpPSh7kot07Egc1
5RaJCNgsENYTF+wdr1TaxDv1RTmxvG3hTE8e9vYi+GdGyG82Jhlv9adohzLx3Lf/
soMnTjvlYVT83fMASBU4RyR/m80u5Hhn8Ahuvlzv++n894IDVB8mO9qaiXOhf64m
O/1AtTNm2m5HFvVdB5i0K9y1+RlX5t0GffGy7EDy1663IFS8utak5tXI60Cbp3Xf
QVcyMq/I45D0d5fKMJR8TlaeNJdWlnKRmxU/5FMewOObfe0qfFrH1drkSWvI3kSY
4L8zj2nASvb15qCCbDa4jNADzsgBr0ChIQdc6Ex6lkRwMnE/FkvMWOQOOBhzfmjJ
NSJbK3bY+JRG7FJgGOPFxOjr9Li7hivZYdkvG6x1/HYcUiYdP9jwqoQIWxMZTKws
sdWlnqM/1AZ3D3Vf7p6lIq0InlOR7SG3qH6AomGR7nYH7msAGuAPD3agN65MunPw
of6H2sAPyd3l7PaSxaWL4QHhn9Pzya/MFIIUdkb9uqLg++CXg1q7cKP1sZW6XGdk
Ovy8zbcGcX7GwV1JCOj/z+fC7mg7noNmJQoKnt1/WdYCMI12yTfI4QyN+Mo3c2ZQ
UWK/384an8C+JA3H+avtyC0xf24l0WO8iE0OcZ908kC4kI8FKBlFOGezEJ5DDpHF
f2iNY1CoiUtUSjfCATJhc2lwaBLtcqFqziLksV5sfGRHxAnutP8UymLXSNJW6WEx
vdsvtSXQG9vjy7CoDkjO7bIXH0PXnfbC+yZZ2dZTc5Aq2akNRih4lD94iVdbK2dO
7kueA965M5aMOMOhu4C7uTEZv8qqdc4JS3WEZHBRI+G8Cy5vxxoztohL0njyBEbv
JoDuP1WR3poEk/cxd9Ck0Q9IqHszdkswDNgfDLOgE1WgPKs17WT0lFqvpFiGTPuJ
jZ4E2tqem8hN6uJ2uC32rKdeillRpZjqn8cXdYVhD1yvpHoAZpZ3rp9JDqamdBxT
gbozk0gpK/+frPZmzH0/R8DZnw/wlvsbZam47//UtBHdlNUY/97jQcEXB+LBTzyW
Jm/uHGAtqy/jeO0tv6GBWdh3DcTDY5EeoE5C8cLtfI5IT0iIEPs4gVHnoWcY/7GY
etyKhodmOmogZ6fd3OhR+yNFk6Ytt5i/tSqeOv5FFrT/JzIisLG130qu7kV2Tbn2
Mo1tAiXMQBmldWZAbZuL28+7aFKzPtlhTdV09duXBhSDUNd4brwDysDAjdTaLBoI
0fvSC8HgmtpZi5FcKd+OaCU5imIT3HGizw0wZmC2qjvCPB5qHN3bIEdrY6eUBcnz
gGJWD1G4kSID549YgYsR6LqfKByD8OGpNKwy0uo5T/ExPJL8qD6ykbiy/7vheOc+
65vJMO8DHDFyB3XVCSJQSGXwmyFm5Jw9HHBvQyi9zxqdmKgtUYC8sXDUCrcK2VzM
AzFcJqSFxDjtCbbECMaZFU5swN3rhDOS7y8E+kUsMfaHgZ+VCNxe8viPiqH5P34q
jYMSphhffsV6qYwSaw2tz5zemwnPOiWgs5+y2WvKH52IukVQ5l/0YeA3S1PbVoXk
3F0BpYjQDoR60vBh8o9v5t4mNG+9Ar8l8hZF765LoSNcxE/R1fzfoxHsFTTm7I4n
rL2s0CcigBeEcHJ02uFcbAgJXafKSWc7o2ZfsWdcR4A08zwH4enmT/mbss/jrQgf
LaOSrg6GAamOYi3O8ksOuR0rAauIwBL5DRJyzT/mSqdnP5YZm4ab5VY7MAUPirKy
KC/EmqcTYc7SmsUhmmU+7/052/PZDM7X3Bfe2pufGazV7iNtj7+fWHVI7zw79fv4
xeVcK+DomFU49h6rD6JdJ7g+MZbyVOk4Q6mStfb4OfagokeDHGz2lwr4Cd5zY7OG
4bpWZjPeSveFJkzlbmxw0cAYW5cvq/UHuoaGiAa63DXdvtlgh2gkUL0F3AJLI+rS
m2jXNNgf7Y7glmmYXObxcMgNS2JjE8VE9fQkMzUWv/j+q7R10PYXmmYwLN46Vv9n
sUbvsgrF5s6WAPprpyQfob+Wi5d0zArF4q55TTfWPb+/DD1XWndkpGUxKUR39sO0
v1IOEf4mwP6hRzVLPTAQdR8mXq9fD6gZ3G7zUBUi1QyLWUyqbFFbmxP/ymAC6xfN
gvPm2Lk15ha6vMmo9ZF88gDSlwsk+GxzjX8bab0PfMf+3u0GJuOiNsabu+EN8Lav
sqhqUZSbcuKvGfKCx5uPSsdPhEaunqGs3SoKSrRVqEr7BQdmzrSu8/s7CTaMwhYI
Kh6seXs3J8i77hgprDDXK1avKXpM1rqJirb58SAplv9E1FBTng1+KZ2hQJrnQszx
dayUA+xbQ6SGHTGRf6+8xslM8otlMDTBb37Sx4RH/tQQUHB2+g/HTLskMLFocvdo
e9nvRARnuTFH244pLC/ME3TVN6r949wxCWte/XtOIeWPrkyPb+b6XzBC/4qiaB9p
mBH3nk3+zm3cSDU4totPdIOCPyxq0NTlc15+uPSy8Xfccd8unTZXmZHVuZW8Dkus
v82Z5kloQUefb+60YuHqJCkUvVgtNQfdMUyG5dlcpGq7VQ3pONphVbj4vnNq+0uY
sdRs7Moxt4vr/mHmxN5w9FTF8t18yd9nW6TttaAJ5lptUdf2CZgvaeeHSdyM8NlG
Rz8Eje53Uu8fZXB3MNekZOjSH1jpECI6REXVMDOpGniVdpZ2qkdR251LTpbk6qfw
ibxaCVoOl5m4uzLHh2ln/a8UhDVWdSoY6Ov0qe9/wONdwU0fyl7+dXHeTxfF6EB7
S73hjjuFa9yc2e5UygJjOKO6g5KPp27/Xuht+9zV/P9L5cMDwajTi2UwSiIQUQu5
RLdCFT36jqaieIEEWPgu1spERXFJpHj/5fQF7kD9PO0McQ+0XTVC/s74DEsC7oz4
BF0K7dbe1DVcg6obj8he+ILGi/MtLzpwcbWSU6UHNEmo8shix2rPXdoO/dnTZJUX
nMsZBOWtl1WLeGsaTo6HwfkSA+z4eDfjYwT6S9CTBE6oC/xhSqMF3FvOsHrkHVrp
9HSTz8lQkfpB+KXkgJNIZ7muHRTd6UeewYaIweS5nUq7qKNUwS6685Zxiu8B8a/7
c0xofIsjXOmhqw4pZQezhh9g/+tcQs/7MLOSYdzE8dRWQOvTFEldN2w4JwMfGMjL
WsMw6lCEq7PPLTSGXHbSM9C0sMbLAMvf+jPAeswvaxAICM4ApYR3ZkSb3JIqcNVx
CF41iSoaoXXlzCx1FIPVkhLcWTvC1O4Fn7QAd9OUh1aIuFdb5tpklZQMjVP4s2sS
K4Hr2sVX+btglDnBueEA8qK3l5EJKzGJ5/oEOKjIKrpZMC1DBhqRvjzigkqAve32
Yde/QlAoaQXTepf17nzvxEFFtNDYC7BrUIuZxig3pa91QqGJjOEHLzcoBKNjOlT4
ZcO/F52+F+TOCoyAbctDJLRhq9YG/+usFC/E4sHUFSThtryDbE4CI2+Z5n/vvkgU
CKjstga7Dz5IRV6rqbfA/c9AyJzoPnN2Dr9FICieNFJId0artcHycE+lcJKMtroH
Wbsrrn5XlVbJUa8PC+IJfy1W60XfhLuUKcQq7wVmclgYsQmJSAgqjSuKAFmKVbBU
3x98vEp2wYmoWPrd0Hq4xiitCoRO7KyefqnPKb/6YUMdV389Jm53IlPedrvZzxm9
4M+4Pcr6Na5VK0+3L1AW/dKWSe19gw3c2O11PoqcLtthSCC21OUgo4pEtZywvPQU
Up2uGs4UMBzkXHAIzM+mt/QknMeLC/Sw4eMBTvkYO5qpa/wa1EyREGlb6zXuU6XA
IZ77AzdvNc3PLRh3SpyN9TgqtkRYdSIvGUihqel0iBZ0WBMg577XS9wiJJn6AufD
IusYSGtRB5kjf33g8r/p50Lo4/ez0ejB7GgqfRx+Krx/pN1zr+tg3zR1IHxR2uS3
xVK/Qtij6r1wvGlJOBtw9cQW8HaLjY+M0GDJW3N9kKmrSNZaQ20cQre0CX+SHRGM
G7am4zE3+6bw5EfmTv6kFuUspORBPgSMWHwlXxUZiKKuza3CpzAe4viJiKLlMWXT
tgfP14+dsgMtYMb0vBpmTPUPOeozaKLGsoB481lythnqa4eK2W13C1uUY+Q/a/tt
voBpeTdWX3ZSlr06LmNXBa2Y0yai/GaNXOseTR0QY9NKiOMaYip1j78QW6WPHXvd
jkLlSWM58oy5W2O7yLLfCDOQCgvBTbf+iEoc5WeXzAAOIMBmxwdNmji2qyD/sGhH
jUQ/ZLDfNJopvp9KRL+RTt8SvB/WCttWsZOYpNm6/7nb8JkXMdrCDE873O7Bvl4G
Cvk2Z3HusD2hxtSLQGk32AJxzEIJffQ64Ip2mN9QMNEem5TipEZttuNUVqiVMURm
6QO4j7NKhckYUOYfukU9cGtBooWCZ/J2ij26vCd56w6JT0YJ8qYPClxXCdiMY1cf
E1O5mmRJ8yxKhv6dtFgqYXi3bAWwf2WdZvDUtH83n64lOYdnGdrcmdSpkoz1XfI5
TGJ02fnk8/yp1lmZMx9W8sJcqCS3kd1XhwZMuJRp2EYiyVjS03/VqxLdjVuor1Sw
sRsTr4zh6me3pNOQqv+lrnwPhG83xtguBbJAe3rhqgMSV1TvaTQNM5+WwA45nqPH
5Q9E1UZQOFapyfKIasFx6SBflA3+vDn5gyYAnwAFZ9bFG/og6nrbLD7QGOHIS74w
fzWcHhOYztSMfZx1G1VKVLFTwEOoZNY9CMuXA5aMyFeiV1S+q8GnalqCLaBXQs9u
9QFlDyDiPZcLlryh9dQQcZChT1vGvE/R8aUaYnGeteFThog8+58W/4SOfxUokJSW
ov6GqgSmyq2LKNzNoerlNgvRGzmsHVd86lvBaBor0K1PXDWVv7HEdg31YMAPOAIo
o9MCbHHkdKUMVaMchypjax+UVnSCx2og1usRfclgbCTUvzkv54xEjAJJPbLYW+pF
rqd2kbv18JpDDsGnvXsE6lyHCk88nx1kX7lXb0uyz8drNeiFSzaUjaxEFDkgl+p9
ie23+s+pHH4NcaaLTGGeZpA1khrqNxnsq5zrf3lp12tlhNmD0ZxuCNnxxPA2FDNS
MvObntrvEkZgLqQRieWdHQ6PJ1PsNvy4smiClAkr6hkzBxhsaPPqwoAJB7lsbf5k
pluWIzJdSCEjhxg522dG5jNjaT1tEcxob5ExebXodb13rjTznQyf4K0oiSZUI67b
7kMdQtW+smIurEgM8xHIpwpoWVQxMV74Llg5OOFy++eJrdijJDZJ55MNZY0UQLo3
WJ6nCxH5oWiiXDzW58LKiuqd5riwPLnbKwj/4zu/BKWZIaGku2Q9+o5hXo4ff9cc
eCWg7zFRJzIcpqPUtmivnTxDX6h0N8rSI5I4gR9zkWQ3M30tLwlnYY1tr8/lmMcb
aCY1enjA0l5zI3OrIfGbg+Jxz4kvw95TxlS2tYpf1NjX2pjgBo8zob5fRTesrKq0
dVCoO0+wHeKvXTTE+RN+L90yAZbhjA3dFFmlxueEhYBtPTgVNLfPdXeD3vLxhJxm
rmIo2gPjTNeSvjSGgV/gDMIG7al/CSwB9j4MNsYbj/wdyu6q+up96o1pg2wKrxY4
S/UqGj6gvygx4HQT2yPDGAnioSKnVbmufjh3dkqExTu7h7dvK3PKk9t/9e30Z/lg
Ks6Y7o9uXS5HXBzodgHbY8ujvQxXy4Rn4Uy6DzlVO1YaUFwOW1sUcTMeqic3UyZA
BWPcgOsuRjGkKQL4/+UcsdJvo/r3Tn1I2bpJKJx42PK+Jqgp0sLgicBt5op0CfAa
szB2RaO+caOEDk9hN7oYF1O5zL1AkoR8b7Ivd9j60wmuVOqGYT+6crdTgt4QAtcf
pVCdZJlyLAHGthUqHEArLfUyo7EySOaKI8BVm8Jb5hh0ZA0QuMOM936Ja4ZEA60D
dqFhlz6XV6k/aRDv6j00+JSVFVez3a5VCXj2lxNGiFnyqbqgIgYQKi6GCuAv5073
ei9xvsdRiaKtmtmFa2Y6DWFy9jR/59IW424geBoLhpJ8wrXkIZBpjho0A7ofxA9H
lqwt0RR6o68UD3k0C82ivIf+QwDMtSltycyh3FaYIKn4vm8wrMZGbYPIULD4wm9B
ANbIr64uXa85yoAMljkUhNuoO4g8OflVoPiCweYqQ2J4PoJOwh0h+Zvi8oK1Yftq
mgUe4su48OClSfX08CJuY2mXvENkVP2q07vyD3qgOhbPKtoZWh4ARkAvV/kNOahB
K9cvH/IZ+cefKa10q5lLQkpl9OO67dcyR4Ur8z6/Gw/y9ciiR4zHAG1GzVoMhpfx
pQJpNrkehjFt8VvK5uQUOq7RluKas2WrHz/LA8d3N/jCQny/gqA13LuE6gN3Bx3O
QlsCQVRBGB1qsZqt4zWTlbpg60eFvekDyVMKODhaV08SIw5sxafQV4SYp+w+Upky
fjtVHpRN6UIOVUa+WmtZ1kLSf0ALDFa8a/6Riq79LBb6kpfmo41A09oRmGZOuzJ9
1jNhFtWE/zACmme2CRjoOfbefv+xH04SkfGzqxs8YnQ+fa4JGxuGM6UnvW7ZPSd/
5pHkW7akfd4VQWOfNGNPf4kLehhdMHk1b5PrDaATHQMGPAII0KlxjInzqnGlpNwu
Hrn3sX9OlD0qGZ8Sox2x0yQ+mzFSKZPg79FjlLcnqe96KI/fmz9owDTEnnNZw5EL
hFdzmIKl2BBuW12vJXoWn7KE3V2pjA7tm3IWQivyxjBnD7ysoUfTRZFfyrc2sk/q
FL3VQPFYgmjnsdTPrJOH4Mbwn2qbO8eFxbi/l87dYQ1IZ2V4CQbk932DfIbgIp2n
PpUJZQqRvPdwTENBkYSoR88FXpkBvMUzjSFbaUhDVG4+B70z2RRKbr5Wy4fhqwe2
0AVd5wF5CGMxUbDPc3rWR9YpOmXY6KEA17llbe4FY3SJXvWkd/S2bVxLPhatWAWG
cykAEj6dekjs8rAffD1wL/fMNSgdAkCA7+zqFiOTVw5vPCNlibo6xPeKHHhjyKFO
BYWQt+bhGT4hNWdXGv3oMMhgwGjcTi9CQ3eL1aHHdmDpDnIUUnix3GKggTVLQJKa
Z6n87qMXUgX8Xkuhg8JWJAjHOtoSow6IWhgkJS5oQF8NyP6ockbiTcBo70+yUlwk
ulVQm0R1Q5aaoyqhnsrSn4Fz9PwDO0zfRyZPle7OiJJaZvATg11iqEMLLIYT9qtu
VrJUGsAnqpvchyx6cwZ2xAmAPLkH6lwJU9yr34Dgx4UtSOgQR4mn8DfHVyCwHPiJ
AhFfEgM4KvLqRn0X9KnZ39YbENZBbAJOoRfv/D1+DIu3CgvNlDRo/L3qxBNJmP5C
AWbDQVszCWfsLeN/SpBiV9uCJRBdCerA5rl2zjaCuuYyOXMGHZ2qLbgmQ/u5H01Q
CKK8RoH8VC9jKj1c1EuRYhx0pya3oQxz4Fo3faC7YTB1uA5oJZ4S+zAO1pN2xt27
bZy026+tMrvxz5J0/seD//rXTTB5nJiiMKFgb+TUBipaljxOfZGQJHEIjFCuGkvZ
2ZdHG8zAinM8t0VRJapDdrmCDDhDnwKUzIM28AVen0HJsMKAJ0tS98HspX52vFVV
RaaINJUP40BcghZooj7NANClq1RYXpPKdiC/O+5qoVpSsm9Z7Io92BpaKSCpB4V2
nInbiRS0FOs7hh39kIyv0RuBhWuqAvVj3VnAg2EdMVWdl0IISKzU1V/uEg6oma+g
QSkStzKmPA1+eY2xOyYkAdcoJMg4SZ4dR4pCUDeJlff2BChzjxAY/fNYhIjwND2A
eePKmgt6OyRdKmjDL1DMN/Z9AjzTCn/N77TflBj7c96wmceiyRWePSu9fiuxPjJh
CICpnfEkHZodti0Feb8fP1NKAWHdIYVTugla2+8Ih7PBRnsHm03xYecfMTFiNsQp
HVpC1OnUXBN9SQa7JYTUAH0YWr8kEGzAPVYUDidTGC/QmJwYrvsPSpGOxui9J+T7
hkC+oVeSBnb8+vrqDTSdgtPCsWAYjMjkpPJiqb1+3tIDOYXJY6kfgGnxSiwNpEjN
dn5V7gp3jW9UB98G9SVX/jsQKuwY0YcaJnKIuv4VcC7EesiGn35KummZ+CeKlC7t
dOnQ3W5P9hdA+bHyixoJzgb7VXKp+KIapz4YtiqUVqEAQTzNoVjbl9YheApPzCxw
9Xx8e1paeYaW7BwifVDeoKevk25+1k+H69wgyGrKwYdghUIdztPDH2c/Vrs/W6DQ
H4VldQWiZLqYA6Vu1MR5pXDRr8KKfygCbFF8oTjE8N6RJUB23HamkAqSDxoAWWWt
yCyAQ11PIVi6Cif0Hgd7TmDPdorwZrv9zq9TzAUIjC6dgdELBo0F45tBwYDT6JDx
SceMz5OZPHZIu6dBHxxTmPkButirRAlINc/4+IYj9MIAQV6dj2NNDAY8AUOP1fmD
UOpRh0P2Dmc5a4w94IqNBNEaNoxAJ8xJsF6qqKdizFhb35MdQCtxY4XjryBpi5Hu
jgnmi4sKThkhHt4TEux/kQX9Zfno2UhznbA63oHvRG8BA12BgkhB3n1KC8zQjrea
lrsc+wrdJmvLjyrNqpg73TZyEZ4IyOUdLxj+PLDq4sQVfLNs4wTWK2eZdV6NptfI
pKVm0tZcmn0yBLlkc5xf2c5qE8pNXVJh4T76QPM5phalTduKtId6jNPegL8xRNaw
uI+Pgr/1v31e2gYA6tLiIeJJsj8peX7j0IH2if+wGPXM3WbkWGuFaxZJeWFIHHM6
mfqA8damE15smEqHUjv/TEZckPXweR1p49uHEU3pelB5OubpBxnHeRFKQPpGqny3
szhb4NWMBUxAZ0m0LUSYA/ilCzNwyw0TeG+a1V7AIHmUR6zVswHs1QHzXBLyhXtu
NtZEGYSw6YlnQyDe6IokoLxY1WKl6Lzwk/AAb8mXLkt894ibXrwhgLbXMDgrExHi
fjKiiX2G1Eoyh/ZhUXWp9k1ts3MJ7wU7jFhoPBxp9xJ+BdVbAl4QOdil6iDey7Hh
WnYPUuvbkH7ALmz1OUNglQMMyAioYGtbp2saz3a0KuEFzyEJ4VntJmPyW5OgQOcG
g26YaP5E1ezTMYX+M4plHcCDPcWr0LMbL3SWkXOAoNBzUgyo5tZdxqARn5oGpSQy
WFQE2IMRoy5LMPt9DhOwblLzSdv21rcVS50NxJ6yVcykXhAFuJrO2HMU96ZRwACE
wmWgMEf4c7kQgalFyyPYaeanSaEx2WJp070wR7GEX2yKK83Qw08LL5t3vaLRFjCW
3AtTPxyE1b39b3gpo2THYW78Dbt2OLu9wyJMYKf+Uez4VBtmftW8/dXT1O4pf8zK
Uks57Ce4ugxcPHO2A/TzQGayWY0uyr9P0Ly16lkySS2pw/CuhylH9e37IEldG1CV
xcmWW/QLucy5yL0/oZSPWuSOQStVqxlRJWAJ31wiiL5yvB1pEJi5f+vithqtZ31q
x82jgXx+UbP7bQtUysOoNN3fx/WhEnyUsd3kmc5uYrTPGj6MYzKWNh3Mn5HtzG0J
iM0wZJgdR2VJCqh4uKw6px2uHYgB2xGOkmwg6eHZrYGKRle8O3E523IJkw2ovbf6
AEBbDzFwo/5AIdKDVAnHlUN48cTawZiG+dH/+L6icikE+IF7rlw9NiYrNmFLQye1
m+zs5S1GQjS0QgiEenUKBobSVGBD4yq6aqK5HCBKWJ4xCkxhTAgFa1KzkVuERxJn
PqlMeKCAbwRopZw357xevarXSnnCX2uj79ECl9ETacyxJTONXA77/afaYm6lc+wh
nYE6QHSO0+gL4+BhIfhr1RjiDybfFgGo5vG4BBAoXuY22fNF3cQ5e9kdRPCNRS9n
1VZpequ20A8NhudLiwQepWdQb+mkJR7YMoJt7FkGFd0yIF4uD2vtWZ0YUC/fFx5c
9QLFm3mL4U48mqNEuVFOhuLv/hoin17AgDHvpB+CP2Sc+1UtFWJJZiSvd69lFVJC
vvNR0MzqkMYdy9LkK2tUle5x5EATC+aNmOu5CXBGq4jmCLN29mX1kuXex7M61frm
1TryxYDfQ9dMEhxqqQEfPDOljK+I+LXW+Jq4fEXMEviyMIcpV/zaSPva6jdpvTiE
SRXzSBTQMYJ68q6CoyT9Cu8H1qDwrpfvVptt/fM2or7VOeB0xVonummlL6CJTbdR
Jy/q0mun4YdSHLovAJdLpeYhVTJa5qqFklLYg7KwW0/t/UbxbffauZAz9oL11axD
1rR6m0xgR7Yv0TtaytW8KfZPjAUwHzq0zepNLq+eOyvGbBB6xoS87rGO+R7TxRg4
BztLeVmxSsea9z5h9kfTq5BMZLyLilHbmpSsxbv8VCHgbKQTYRTC+nxNTm9LmNp8
UoJCr1Pb13OYqX9zI2xA2J+dAigSev8uPr3xTlOr21Iu3WOo7DBvU6N6/9q6TgSd
QddE+UWnJW7yIHlEhRvmSBsCaksLjXyVO3my6tkv7s6xB3O2cqzcxv95XsEujQJq
+aOp5RdECzQEtFCWoM+r+w2N5hoSEkV5tpWunhoFClu6ul1obHS2iuWuxUJomsCw
50Zg78Udq0IygAd8vns+yC1LTw18JsF9LqUNr3vKj8M/dmO0QbPYFwvuGd/+D7vQ
bwQ2vNHNEN8BLt1p3c7LZOgCsfvVZHuUTANfgTFlWoosWCeV7dmB2leO0NHbhMkE
yEbuSJ231ys6WoiIFf3gyn1zsGOSHy7VB/mt84X4/T2e5mTXt5LFje1xu7kS0W9S
mh61xQACN2wOX9JqraBOaVtpUPButtx5RkQj2w4F3Q2noXcQ9fWeRuoKU9NUtyBu
b41DnwurRBdJehZSTdoxjQgEkkYoKxXQuLi7OTeGmDrVEampNxI0WBTyhvmrWAA0
vZrocHIfoOdaHJVoSTJcM2T7tPvcPj5o0sgdvCuwwyoAMZgY74FD+chhVQSnuYgf
LgQrXbarRoWwePaBt499KPL6KVDU1BwZVPDciL9ipmOPPgl5HAlcCdPPT0w10YBd
oybBnoG2QOO+MaF1TGNMXjwiBqxuMRC0RqvR16tSzdNQkjrF0/y7eXxyYfKW6+81
SLjZ2Hl8US53qnZSiGFKTiipQSPNldeY78hlkP37H1HxFfp4a2OXYEpmW7CjoLww
aELLkWT79HjWGKPAKZmxIaHu3kLuNlRHfo+MSFh6b1w10tFchZw0dpTsbuEexSRa
zfXJ/WU1+nqyyGvuBwrmbsXKy/Dy8d49Uvnv8b5F1zqifxQImxegdH97zypllIea
nYr/VdnlMBol6JZ9m81x6rmw/Hl9GusvYKYFmD44mR0+cIQvPSCgZwgIsQjKomv6
8LQbCCseA+ZKrpErC5ztKgW03kp99sJ2r6qcLdjDUY1a6gkgFjlMPuMn9nH5Ci0u
eZ7n8ItnFHiD7Jzhosgb58FE8OyosPZ6FEZkCWKSamWe5NxCpyueEtEKM4qyS++q
4v2O/sk5CbjzQlVWvHX5gMb5X3G+MdBrvsAndhHyYcT57yeuDbnnZZ+FPLCmDsZg
PBh8mp0kIo3N6Xgyoe63k9xqFvmmemBTiz57A7I98W9kbxgs/WYyAdQGIX7jQeEk
EmTxSykVAwQ08POa6rekMbSvmRMHrxVxxvjN5AaZwz0bMCFt9j0ZKulCAXGSQsnD
tzverrb6D7+y3Z6WNsZ1m/UMHqe84ekEmTVrg2e/NMbLrYuYpwisuIe7bVMnIeeW
0Ea+7nKWv1ngqk/Ey2b0/Jxtwosh3mkiAoqt5jMSwxa2FaKwQmh5N46yFGFr2d/E
ztOkpyeO3aeeirbQ0wRoPSNCrZE3CF/Qc2f/xi4S5Mewz2aatla/blm7lJNr3u0c
bWApXefDqAzu9qlcCZMZvQtx1tgWd9rsIPtBtZaA4p5947V6234Y4vSsiKNkLCVu
AQCHb2ntMV9nAr291aLFO6y4TZxvmXeADdptTdBcxX8qpV0o+N3NTWTA+Q5Mx4WC
M1klER7kurnqJt1USbKGgGDiL9sq4dAeAp35ry8trvleBObKzKmO4xoTe1BAXsmU
BAa7aWYfe4ezt+ld216tJ3zUI3BbbZLLgCiP7RnqdslcBpd/Sr2s9oVIPGkvN/SI
KNn2KWK5Fy30AqBX++g4jJpthYhmBA8CPZ0FkJi4ie5/khynG/grwBQZlk/eO8dH
Sjgrdo4xuGLSnCqxUroAxcRWi/AiTh4bxZ39dOIUXqttM2/FPtwf8WLA9gzrz20T
HtdBE0XqKIxvrx/uEcft/cOIlNkswIH/NcurHSzHrWmaNmQTuOCdQCbo0aKoxIIM
f3ziQKCnIHPAnuV9ddLwGTLxzkSAYfhoI/4rVbKU3UXvTaUJ/62uO/4mBHs4sme1
pkG3vEGWgchV6YBXmNFx+4sCoc2LSaBWhsSMZUgGdhGy52lEqp9V9wrFhgB++FSA
EzwoR4lvCwpNedgk/MLJdYr3pRQ5MhYiaLgTHEaZvdS1z0u20PC2s1Z/hMUeVphP
cwHl6EFDqh+x7ZQz097hoWsm8fTUqfQ3fEbsdlnvSopehiUniDDAxZfcOL9n6Hwd
1ZC0egfdzfrx2bAP8zraUGVwETC7DRP//ipo2xh38lfM+ywPxYVqsG6X3zHGqpXA
aCsI3cCKn+KbEiY6CPFZBl2JtBgdzDFHZAf1olWxD9699/n8SLFwFPpl/xstDvjP
ylQ0iPzKCVi1bqDaG9QMcX+3h9z4sHRJD8rjg1S9vr6d00dhHvdMzW+Ny4E2MqGi
XJS5y5O727ngMg0/mq0YLpyVrOulolP5BqWdHg880mPZs4dod2N5Nmz7SMCLTQGY
tOf1sj7M8YS7xM+vxbOb4ZAicUGvMm3QTLhgbEl0/zrcP+SHfd801pQV2u3rPKK0
rXnkvJGlo9jPyp4YoGCKlevfLw2a7nnK3ev/MI4WRFySNhufaqXk0sYkcaqI7JKq
UnTD5FEE3M1JZR507KqX/XVbkk5V1WJITCpmbCPnj3S6MHwR93pwadaq1w7bFxZ5
ou9psLGGrnR+Nir31wNfymvbIjNImhP8MNXUAZvOUqK7rqsMqffuymA9reeD/xHW
DY+qwRiAQy23jHjoHFixKHd5kNOiMJsY5D8hOlwsDmrJkHl7X5TdN6aSj9B17a0s
CyMQinh+TsgbnmxfpHhfR+68KXZpCZxJJjwA0WMUo6ScMqwb5OYVwxmzrqveRB0m
/PJHm1fU3iZwafE5xCqGhFdO2fuM2Erjuh3rsAY1lEUmVfMrOQqMOZCY2NLBHtxw
qFISn8R5MyUXz5AJcUXIc+WTDyVUaBA49gGIXMTXck64EhIdtZPY5gvweNx/perR
Azj2vPCOPjtvK1KQXuARVlu50Mk/aoQcYs60dlPzy6XIIXCUmGlCcI1iGJ7CgqnN
09nm5A23V1jsx1KDnGjDyMMmB9YM/8RVtbqscB4+/9enK2LGpahPgp7C0myAZrt5
D2JU+OC8ljy3F4x1cK7FbKI0YOydezoXHr7ShEe4HhvnY/xIeRF7zz2xAfRj78OT
mW01yt2cSkR1j7pvdy/OgBh1wLyD5vBPps+Xs0bL5Lb0AMuWamNziNlLgusy1U7X
pkjlKRjFRvW2sFtnKZ5tI0HL1jmAWzXpmUafs1RUzJXNipgKpnOUl/gaJ8aNfgh3
7W4HaO8ewj55CJI42Gkx21sZ3mI9mQPQvf+snU95GKeDNYGZKER/35BidZo2ocrs
bI6oLWFlXvvKBolfpyaHdzb3BtvQIwvnhIeyW6Tq1m+TpcUiE4HPn73v2XHRAm+3
4z50fIorcq5vjWH7mnVREJWFgSwzfDFf1avwHJiGPyRTZOOYK/2bDf4LAi5AVYk+
qJh1zduhLiurNj5h8c3tty8D2hwge05Sja1kh57ezXN0Hjx/F49lJvBsCYJMDuc5
eBtqJvbxcusf/3sOBHIpg1rHNjMbegAeSEjtlRgt4wMfFIa7pfYOHYnHg1vK9KLa
G1X1WT7FOkA1jweQ46ZPwS9w8GCELzeWU7zqqBcOo1fB/3qISsK+W8y2kedELVBZ
1b4l/4vjiMtqlL1EhFdaEWfBXGXcl8YK2AGyMPgEiQ2XGyxVKB9ZqCLQfavsrMmW
L1oGAzDoZEzSSQG/V86fDLZ4P8mdfW8FgfuzKlfPuh+NPbDvEMtL7h2DsqScoUJI
gXSdLCuGWJYPwaeeZIV8N+JD3ValzS/Q+pbuUT5YcaaJ5JK74F/4TsEeudE3QAwz
caG48aKRg0Jp8n62RVLYGrkvIJOmwSx1VLBkP1Vn/3keB493rg2KJTGGq13lhRPG
GOXVIPfhaXS/lutK7ErfFP9Q6ibSXNOC8lNfo+OypeITvAWqknGpzXQAMpuzFKiK
Z7ymDZwvFLjg7eJbyFZa0wJ8wU6aX/WdQWL53n3hXeejg35pzwFZJH6Ur5Ave60j
FWnql3XX36A86ySQZAu0kHwx4k9weAQSh72euh/H1vyAO0ncMJdE0ib5D8xxcsxq
3uPF8rkIQjBZNRsilheXIh8xJZyV2DWcQccWgEiKhclBa31wedTo6D4HIsJg72ss
KuiF5dt8y5onOzmcLGQpLI/e3qR3XSr9yben6E9UR6huHtroQezCOSLF9U1i3xYH
tDnlWmYYhvwfERZ84IfkpLE6kndylZD0qJ6Aer7gv5N/dDbtYBvyZo9tq/PQhJ4S
BtGPTQnVgt1RUC+rcDgcomen3mgON2Qtcq3SiTAdHhQ+fyjIa1bfAjoUAYbt0NJC
vHuapSGEoSL78CW1TU8VHbHX4vdxawOaxIdqU4IFi/60jqqdDuUR4UFxZNkqXdm7
FX42u0slZAhJPvrsU8BhTfEugcdxFaN2+71oK6oZ83KmUMfUsvLjKZIFdbrlcZBj
eSUvCPGKGMhifDJx7GSW7ITT8VZ4PdFqHXq4JRb/jp3RtAdHyXe14vVFZ7F90xEH
Z8/rV+X44r/8MYrHhHSvACbTKxUZ7VNRH5pNlWmTBKxkaNer7+YSRABOp5pl+rOs
f1Q5Dd74bbLS8bGnsNxJkRRlpKlK5S7WNfqABh2FGOcq9atVXPhg9fGwyTJtEcxF
fBVgvXcJ9AXn4Vu5nO9Xg2WQNFt7Jd+bKh5OHIXJEWvsZRdnKA5044RCAreFQRjI
3ZcK82N6/BbbvhWnlhvxLMlht6ruDigmavOTnN9TsUxpeWhQl8rOONKdx98KGmUf
XDt+MyyJN7nzjSzjnhAJbUUl8TPONjvh2XVuG4aMsQQ+WdIb2IAA8UIfj020KVx0
LnPlae2tWkGHUcwEev0MzeEbt6TBX420gyTtg5dKxRJZwfJfj5yGv40dICyQwZl5
7o+huJdNfJWQuJ2z3PFXYjCq8OcH7O7V75cG72VQoVzQA+BPouKmQ0BthGQ5j0Tn
7zl4z+gPDPQQcLWKZiv9n/DizjiRGRh/tpjGpVDJsKyND6YK9uirsEyRuDqgJjUq
po98GHFd9Qlse/Yh3S2MSAMJisivsmdAlRMh5i2mvOvdjbTIgRs3molFV4XEQyA7
nKTvy6mrej3EyONJS85h4hARJPsbBE/+99XWUubA1s27W6UBBdVgyVQ78QXcwxVF
qQmR42lsfYsvuxQb43SlPQRxyzCVoJl6GTaeLp2Mp30dXXjYZCaxwqi3lY1edl3r
H5KKofjAHMsE4UNstvfLRSziOuWnp+KzsO/asEz4koMYzhO5TP7AQGe280B2rLDO
yNA0V2/c/tc1SS8a9eBMsEYqatZ1gJSQR3F7YxFuUAbWZu+aoby6h7vbVB+qaRTX
Vv3surKfZ1JWvdUeQwAApv0n8JitDtGiQxbm5qQx9f0GGm7LaQgel7BEdAr9sQ0Q
r5UUTgOUdrC1NuBmKc4H92l6JvjLNHehFsOFj21yTGeXOruubtCraSeCnaQhqXHK
Kbd1J21hfsnyyZCFJ2haFhNvZjwJ7nrOjiAzQY1U/1pVtniQJNhVPYhDUE2AxO0+
5zuSNfXXtD1/EeJnUb8PQk6XTmTeePNfRu/nH69HXPh2+IIbGZM21uzvZ7T/hnF0
DtQATIIxd4U8+zF+ILNHIgo87wqKDQFmk40sZyeUbmzumSJ335/bwEMj1e2Ff7eG
fpGtjf5aP2T2E8qr912cobvr2+c+aWG17xspWMlfh9bcbgV3nOrQ6VowmE62a2Us
rgyfJ34iFtbrRYtXh5VyIz1SaDSvk+Axbkun5Ra9owSPR7mUY7dWN/lwz6vrBlwO
o55p12dkOHirZYJyyBEK3EbxK5LQAmKqvXSL66rMe1qcbwhctjyaSu2UPnSb/Jvc
nzoyR3l6RwFa/vQ8dzyB3M7a5xpL7Usy2l/RFn7IIzEEzDs+84NJiSuSY1RoABIS
Bx3+gHC7z9qq7nzSld1oS37mvrSrEU3HHCdy6z0SB8X4Y5wPa6qjvttiR1SWCasU
IDAFOJb8Nsoed+oT8FtDwh8zJ0Qd23jJA2YH2Az+8J3Kj9U0JoZoHADVPV45Wv7+
qdnRNkzQjx2Ezu/qbZw9kBgac419FkI4yyhjJgMfVfGzAmWwwntgZX5x4JVJhF9i
zYL0QEe1xPa2RDm48aUaJCa9DxXrtRUzoAELzGd76F2uTrIudyjI463WIWhM5y58
8BCdQU5wcr0rgo5hCsP4KOynepQSgWCkIeEw7R7PTC9LwJTMlnkTpCU5rVxyVIDn
/IQbAK+jjp/CUWUORjFGpS4NTgGRwfXL5KrKQOzxDeYxpJD9CJQC1VNXpHSrZlFP
fuBNJaZnIcqyGOP/OqDsfEgZXG22gNxU2ZxnfFCA88u0udQj5k73uMKnmr1CsF+k
6EKminOrs/rcv/ABmoiitUmKJQwzPiT4oAJPjmQhGHNDIYQQeMPhcZ1+DX66R+6z
DuSKvZenGfW/tQqDMaSDeJ8+ei8Hi1s09xbPxQl17g2BJBSE2YXIhNiv+mAtzkQN
NR7NbDgWs2gBLlDraXtmg5kpvUHep9/hD51o+3PfomAy42y+TopOEwosFrKjLpYk
1Ji81BMb03HfqvgMz31mxLJ6suirNpQ1yB0n/N9OW22Pi92DULZJVKdWCDL4drp4
W/gWgz2EOawm0H3HklvZ/3xUk5qpQgXkdYFRn5N/0p7N+8ySMM6a4yGAdNnQs97S
YI4z87Uip/jb6mcx2bMjZ4SdHlX9nB7H3JqSFDaxeWi3/2nBn6MngIm3zrL0TNwy
581+WMgvV1J+Ws4uCJoNW/8tWq8VU/4za3+UQ9zCRVNUTv9oxPBfqH+JsIdheLk1
XHCf22UwNvFv3Wj2VLeH7RFU/tqgzCjYcb4t3EHiNssmCouO0+f64GQC7kTXGlZJ
JZrX3G+3DN2OlZqvz4BKCtHAo4wm9O1uKqiZPLLx9Xuy48WT9wTGRmaMIAMRDgrU
rupOqYJg8Pw+IiIOn7GmlC5l4iCdFPW7jrx6pGGVG7LBM2k4T7dEdnF/O5mYaJxr
UoZUpb6lk4St7WCx/ynhUenP4Y835XJV+RdBnEkSA7ctSUrUd9h7cLJRUdv/qYxC
2PTMukeLi47BjXrcAYpuoijhW3pegyslcNdqQhlz58AgsBnv786E6msC5m2ifr0C
m6MXCR8hTmU+O0VAjffgrw7r6VZlYcpFQcrfUZNRm+vatpkr6m9rxrEvqIeq6iGe
VlcTF5TPtfDAAufzxa+LqVU8zuap05aQYpUiwcb7s0/1UrJtO7uOlwDjovRv45YR
vWjrVhtCuB5USa5C+EcjYjupxABXswSCioNhx8cXJ8SDQcB0TuxUu2laAQIHLbwA
YazO8Ek6RQ8QToyWy3x/h1cH3xzR2iJNgw/mwuKeGAcpzDVqQlQkrCDdaEdjSce/
+nnAQnoG03nJUON3JI0HvK9OmD37zibrk4/v7u9od/EdEZTiNE66wKfgnYTyofCf
eX3wniGaSRAYy6kKrhns2j40HwoY8H0TX32089hOf3ey5TcuNXcZYsznS1AFq/ws
rl99zUZphehT+mGaG9B+aDZS7eh7eX1c7AAs0z7MA0ueIt7znoTvkJ2DqNYcO4dB
zu62Ct9P+/gj2c+2eYmXaF8RAk2AwewB6039b7pAfxwoCuYivk3kYcD0qaqzGvTX
j32nRnBD0i/n8D6qTJ+5acdE1fHAxzQPwh+4lSvnleO3gzeC0p87u7aqWDSDG9ql
Lujs9ADbu23L/dDQVF+DKcqgzEaBj3LcfIb1baDsjyhboM1vdkkMcy/I2XyQ10d4
eaH+hwOVipC1mBBIz1VjjMBxx5BbRP49+HyqMohsVLT1gKbjtoDtdysz2Pv1uEdJ
T3axTaV5/a9SHDz6k1u8y5HNSHb9/FYItNK6F/oH9ym6LAAWyzO/cFTZlJeJxcog
+xu9ZWccEhBK1dTDcprB/qRmMKrDFOWdqFW5HDvlVXxM0MPbMYr2HZiJ35CZFS+h
janH78TZT0yHupZre+SJB1BojyZmSzeF5Qy/1V+fYEjIQ1iIK4DYw064mX/fPA46
87vqamI/Srh5MP4q6136cTISwNRoF8eJigO++NCnPROK35c0/carUYbavPVB/bZL
mpnTCbr3vcPUvwuptfU1IwbimAml3kwSr3H+zY2qHjvl5sVZKfQNLVKW5EQQMQJ3
ZWm+JM72tFRWKGtoIzt8Z/9acPoOu+MDtv+2vG0nasqxC4GLMoLoNd12K3+qOBl3
wj9blhKlFBxjg7Ag0/OBU28RXSb0EEOQaM2nf6V+0UQMpItqTy8Roc3NtEHoQvb8
vlGL6ieTb8yxr7hVU6AL0Dtvv8gPHKEnV56dxZF3tFTMmoZiXwe8vppc2RULHLjS
EYGfQg9vGVeHvJF+flwqh0REsrXSz3TcuYSsYAKKVDHRTj0k+A1KwSvZPDoYH+Co
wVz6LpMglOSkVURQY43949k8PTXhw6R56imTwF03WqF3oLG/bG4sXnCfsRJx6tYa
ouS6rzVBE5YJT8dDR0NGHnU4FazhnisjL5cAln5Ijfu5yDWt2tUw/Ypk3YyOYQX5
pyC++4KEXwl4BFNh8rbJPBpg/QcTBGT3ryLypY7kTgJ8bQRkcrtHiMYjlRWgk6Fl
SmopcNSV+8vqqJ192cffdZRHNR/59SYvE4uG/D8Pmt4ZFW/m4kZtFAXnJeQE1fjd
0XrFBXkZoKjVqeaPmzp2FRJ2Z4mAi9451shPLRSfgzXNtqEbVWkEN8lS6+B/eHPp
aHUQVST/ZbDzSSW5NLf6e0PMl9NPhDxS4In71yMk7fXFAi1ok1txWVb2wCmaWFpq
zMKf5JXfARKkkeo0kfLuBLxUWD/nFG8laZzdwSGJ2cvVn7rkUzdqZgZwXVeMSa7G
d0lY0Mc3rP+ZiTKlfB2rQwXdS0ycKVtRIdMUx5MqtI8OdrzQIbdYt1ybMNIwlGmq
4pxJJRt/vuEro2tKVQEtp2geer7ddFaPI4sFcBzQCc8=
`protect END_PROTECTED
