`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
heRy0ry6yzsXLjvBB/D9SIiMiUdV0CnxF6wu2CHmpy8AWimqLy+I8gpqfQC5yDOS
MycwJ/Bji6lnVm5G54uAtNVO0BuQxQ9r9b4nb8n3AF3BpAQBaVtLmZYBCag8NAqO
uxFKpVTk/ewX8SOxleawv6bB2SzNmWoZZUoWhHnJC0B5iws8juYIWoUs4+PsMXBT
NBGTeHQaz/e5KtGdOud2rsR4/M/VxtXN3R+V7W0d66mofA3BqqAEZ7d3P0PAHPWP
eELj9ESvIpVgMYfGImRKRdeNcO/+xIUpC9SQyaulPOmd2Yckqi0BO7NdbYwP0FA3
t3IithQ7MJWwkDyrExRJdIi7brLSMduHNGREaelaN732ElFCr4Dyyh34ERBWIupv
Aww49dsYw2VYvPxQoATF4aY3O0r/FsyGnKCaVOQc+cLpEIB/nu5X0p1Ot+w+ujNx
2x3q5zGAxlY6lhSP/WZOfLfxGSwehfqDzjjaOOANhjaTjoWfslsXYZuMzC+bUZlr
Q66KM7xbiAqPEYy67zyghphY9VpsCB7aJ/89zwb9U8h5ff40gZKPgZbqnJ2FpZ00
`protect END_PROTECTED
