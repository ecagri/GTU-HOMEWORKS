`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CXf1ACilmuktuF6X+qOJcoWPVceos78QUfgWyjvfB/kEKasM066aI4V4WqOjAg1u
Z6w5RY2sYSxZceRsZY3QhpCAWMFl3RL9ILYyeLrsKkpnldapI2hizCGqE25KAc4L
Bko5LzBd2hD8wXIZnI+K2+NppQ/UvdhLqa4q/L68cJ779yS1dvEOCld5xPElYVTj
5OqadhX0nikAnB6kuJhjnQKVXWkvuTudmuK3eAkyo0hvZe1vE2AFMIBGO7Sfr0F/
Wpuri5BgMa45nQlnCAIeaVs07fY8B3ZkiJc0sBgckQM5I/B3ZcTxi5JflC9yMFIU
iFZGX46J7SNEvemqMc2+VaAHXDdrHx3+7Dvhvs/b05Q4opbYHKfoHOzgKKZfax/c
zs5arTk7Y7buzx6zSlAcsUVVsZCW3EVe+KNEO6Akzhc5mh7MVEGSWGHJJiEo6oR0
U87B+y7fMfdVonG9Z/KAHZZQHDV29nqos6zvCypKfyvj3+UmmSBVCRFSGnXDIhl/
su/jRFuPxvBsXUB4JZ2gkB7DmugSXVMwx1X0ulwo+QiYUs9daf4m9o9kAHXLZd1i
RNtjrhggwI60HnhxPJPPEVH2VWe7JXJl0jpMA+FA/Khr98RC5PJnEJTyVDpIiamF
4ivdOqweKaih73pYvrr4t+BWga3Yz42xBxM1lkClFMsG7ruES2nj0wXUS8tL5ETm
G2cLKCzeGIZ3XdXHe1sxLRv/kXyc+ayLZwPV976EsIbQ1WE2cC9l8A2sHDoejIDS
k8OShyeqJDizcScUP2S15pHFXuCswPaAF3nIzFj2xuaXZqbP0eFQXMhzSwUuUg10
GnV9Mewn5kifPX1A7L2ZfQHGKZxCsMDYnFvcFBAd7ZN0RjQTTs/Zs0jntqrx9Vt5
dtFzMwnKmwycfxe86JUuKH8tnTpEdxZM+v6HbQMyTYFsPy0N7pY+F31jJaU8QqCz
JDMRjDOk6jQGB3+vcJ21N3nwo4D0BVkC64x37z/jVdA4Qw6bS8yBZI5Au6MG8Qjg
MZXaiZxLdvK5vZ1nEAN7djnMuV3WEgqmT9HaUwXpYY43PNvLP/1f/m1qNPgu1wP8
QREg1DgtMTml89AsRP8bwY5pnFYgLloBqhOo9PnyMUJhe3RlB0B5YOpAjRy1Pjwu
FXSFBkvTLsRn/8G5GhvTaNMDWOEdUdR5Z/xSFS1pItUfGqOy1WcLUBbTWxA06FkY
UikGSXZVnmieTOpNGY94WMbgcMLSZavkbbPw5qjklCyBuZgj0lLl4CT7JZslGZa9
DoJC1lm7glWnVqG7C2l2P1QE8yNSOnuwXIHU1inBvZJryKgXIbxMjLyyTA4l94i8
piIFtHGm6zbP97ePngN52WMcVrPJixVUmJOsA967xpf0OqGTuxF61IMSyacK9gAw
G4OtfvlJy4ehlMIt/TgGnMqdjkUxiZ9JO6BbBf8iFYph8c8xArRc+jfLaNQLwB5P
dapwxe/Zek8nfhBvRSwuCSrSaawoUB5JI91Lxe0Seg8JgVFtoGqmCim7+yU9NIss
yZzsRVrpaJuoPBQix5mrt5TpqxRGJodRj+9m/t9BcnLJ0VjY/fG6UxXFyszvTTT0
82lLfafbr/nyI68Oera5A0b3cT7/rAcMDDscZL52m696/s5GrX891Y0Fb+tOqysc
7eRPKr++/fDk4llQc72USuUhrRjiGQenLTQhkQq4+NY=
`protect END_PROTECTED
