`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gmSNMedf0XtLeqLlraVgfbpAdQN1hFAtBo6vFZBN1hMRKWxJn28iw+5EVTHkuc9v
aA2rmsJ8/O2ySwiB8+EWSnAbe/eDUCGqT44C7UwNsdzl4pNj87G3KdX8gKkBB8Df
DW3Emp1puG9i9g3W05W8so3IrCtQKNOjGJXFDIGdcukB41h4waFkbEjQJaEkcBi0
J980bvPNijJDuV5BwvM2fXpJsiCvF9IKhGH/IfUnZGnP2UZAcAjXuhHR29KM8AVo
KW7ynkWoSOLdViwphw3y5NvA/HvqW5YaQ8BW1AYUvZ9ellz8dw8qCh2xRxmizrAO
rSTptpTvB+i3Vn8vVoKsibhwuNbUdOQItcl8B8C1H4nzfc5uTTY4ToHC8bLwy0zG
DFWivWkE6UBzcFjgUBGAI8rvu5IcBZBx91IaD891RJp2afTSM9RWbVIiD9tm+xh0
IQH5WQylRP5nU0VF7MFHAOdIgqQ6KMCegrshniLOPBnjBwxfCn5tGjWVw3Xw9mzc
MbHm66AACr0CTvu6/fXqUqfhm2cc/E2nn9LH6bwpZbiKsA14Qp39FQcWjnUqzyi1
yof4UGV7hi9O3PzUXH9/fQIMcmGSsiJANmWwk8n2E/kf1+pLpJLETcailh14MBps
RUB/9H6hJ/eJsQYQgAqZespbdGvS3RRNLT3pHNYJTrGYkjA1QwBOZS4y5e8rPdER
D4Qq+7RIvKuRJweZKOSGHzT+PrAY+FaU1ygtN5j3+aZoTGDAZx/uBGCsxuf6Py+/
BWbtx59V8ipZNQD4BrJJhw8XUJCdMjhBU+f0J/P73NG+p8cQsxhBZEuTT7YwqHLc
umMTtlwteVeqza/I8mLQSAgU+lGlGaAOt+zHZpcGiSQzsu5T46MfvyIsciT0HhKz
gRyFiLmEsqst3ghKozYTBcGGRPq6+E66vJcxe2F5hm4RBRIr8122d7EfBqqNDSRF
78HlJmjHsS1ePdWgD7m6zsa7epFwBDruJPW9MPNlbqNDer9fKYl60Fm6WBwJsYpI
fjtMiDN+htsGeyk1RtHMYA6/lJByx+r328PMKKx6ZSTuebKvp7JV8Xqg6e7loKRl
f4EyuYb5SD/IdTwpROyZuc7KDWFFxUAqUAD08EDvMUMe5UTVzkeEBZjs0WckNOpr
h9fMVXvaocaZn0gC5r4GEy8F4OqB/r3qF5wuZK2qkQdTy62O/K9gakLtOZIgZvaX
pO8mJlB/3okpP0f7DJBVKWWghWsz9RMjPQ4v+pDydo0q8eFr3LZIeOu7veq3gdVw
xqdfnhD0fm6av7Lmxe0HemBdycI920J3gl9oHgAvojq5QaEClIFGdcDG70MZAphk
p05gW86i2vNW4gDTsMWI59vGbME0xeX6ioRx3Ch5+vQ8kJ8wXoc6Cb7mTzT18BPn
IHa1/nBWMdTP7qYanKRZywMlx0BGphfqswtsXCv7er4+yQuEZIP9iabud1WEyn9g
LIvC2H+ZJSgfhl0nWQf1zUjeJK6bgA2lcgBEGZbw5zzM+ZeqdGZzYFL9GnaUBz44
YHkyO30MvAVAu5heLNyeG6sW6qZLqWOeT9EP8e6997Q2b7aG4wqEOuJrRMOF4Leq
6UQFeyXEhifC/08dadjddLK87eTAu4Q95sy8N3yHBbQ9mF/7POIwgGyAkqa0Xy4z
2ObmvtFiM2I/M6heVluC7WrAv83mWwx6Id6PBt6R/BBSroO+1mw0+iUhQdq7WNWZ
1XZ2uQK7RFiL7RZ50lAHOqA00pT9A7XLa8HrD2Luse0C8b6kNU2cfvfenc8rsvqr
zfm9z4IeBhIRw+Z4GPQKgsjA8bfqXOoDMOUg6DgdTyXdAvSe0w2GnzNT9jfzohsX
PzPms7DqjrVIAYjqFLFMm6WzOCMVvVPFLcPi0nhZr/ajxO6iGmoZqW0x7xFoSd94
I8Bfu0hA5r2Az7B0cGdj+tv/b08N403fXVNpIJ8ppI3bR+o7VPMsGquUsc9BEKgO
T0KzBB0FvbZN3lOiY/PDesRHxRkj29JGTOiWPRlK6fOn5vsl7sz9afxufvKxTL8W
+skcDXrP3mhCKsPBgbIhzaKuK6O6jexgKX/0W+hJ64x3F3YEoxmjfEVPI+upUARg
peMhDMnQaVJ+Z5w/tbv9J7eYojdBXCQN8GJ1ukxvCpecc7N8qKH6UWsv17vbGf+X
LDUfpcnUPHJcCFJ8GVwG/Yoow8D6bghXqnWsaNt2nanwH71K155qOUqIKJNie6qF
Eu1pQ9173KcnG9ifjyRgv+hOOJu/5l1OueR4RtAyrWR7xxM5e9oLU9migEfDs2eE
3AQneoFJTZTckqQlU1tufEkNGNFSnQEKcAEm/5HO4XD7jrYLKGIIJYz0so3SO+tl
FXHs0k9zPz1IB5EGGne+Tbmz+F7hzquEr3I9OY9Uk0XEYHdb9blQ8ptiHrgznjbZ
v/Anp1A0HW+zX8m0Odmox1XoZ+Y+f8CBTyETxuQjuGO8EehJYdZR2q395YktMEz4
QotXNiOJKvHt38KgwFrGd8dorbplyBXsTu6sWh0vGTVzB72r/uEO2kGKJ6rV6Omj
XdsNi+xZ6CZY0COCI99oTlbfw4Nag2I/Nu1H0DDpt8gxVjH8vPRk39KCr0LLSFFO
QtUNcEh4LnlrOq6h3riFMPZhdhWK3O7IAhpZ0qJR3ZJDOTEg5g5C3ulKMNoaluiA
9poPWbo+nPisRlqkZbFuRu3M5HWRFIcDb1eQcd7qCSGSz4qmejzhA7jWY+FaHvpq
uik60rBOh4WRxfEVWwJCvJjzDy2L2jNlMefeoaPYumGgI7/cXIZ7nWNcELVyeFet
EKzINnqpOKboOkvvi0iE+Ia8DSkPEor4MN3uj7nBdVm3zIPYACGivlufzEnNodeF
u/0NGYbFx/Fgek4jgYtL94ePebd6PUCMr2gMgnqXfD6Tq+rJaZsUhJI0tuDeCKiN
P96E8hDqiWc3OvMcZWU/61WMr5vL89qKUqapsmc4mvFKtJyOgCz4n+qqj8urK6AY
yFcfxBZiN2V72+9E9MHgYrwZWijtKEILOMLSbHGJcxvw+tnB9dkFCvq9ZevNoC73
l8iIlJni3IJlGK9V4PFMSHcPu/31mbPAuItszJ9fddS8Qgem+V627uvWwPU8LXs1
34XLG+84TQz+7nYiPuam7LFyGdtClb0wF6KdZogDbT+CnBMgiQm3SYZZsN1Yf9O6
FFmaSWxxn1cz4d3EQqYpUgNRIYlT5F0kjrpLh6/h3O3hdh4D9HwgKfZm85O5nTPV
0h3owuKBkJ313fcfc63698ecm5LtAaSkUXdsO2plTDUP+s/3xEvxg7uOcUxCi2Xb
/QgWbEyuFq3fb4XpMC4MC5egwpW3Ppa/0G4iVYCkz5qJZ93/05caJKjLbtdN9RmV
klq/vNplBHe5tMF6auO2SBBm5AlBOBYg89s0TNKOQC3coMloMljlltXdvvnhdVsG
kFPfkoJaN49/GEs6WXrZMiz/0kVpgedGd/9HJ5leI14LapZohJdQxDiF1UdMsORh
6yhcxhNiBPNLDUVilCJFl4uzvdyKSu0rmsVM1gUGL0JRuZp0h17IL1ZWEcsCWNjc
9EMrHr8ulF4P2BIrkMFDDYogRkBBxYnxwt5vwi+2v0epvBhDNONVUbC9+ku2D8Qy
1P/dtTxiakVnQQsekepjc3Uta7ix4jSvTrkcBkXH54+i6mweG7fKX2InonXR2b1c
W+7pZzrat4aGIwXTgmm/6v90LAXNJe+CZG3ahWXO5Dz982vnpTacbvazv5k7g1C1
khfZRADycALTQqvKwf/jho9u84VZYoRL0tjCGub2Vf5pbg7dIT9Obpg7/TuvZHAr
qPMw0qGfuxD0IfRwe0mLYTnhjWcuOR3kDw0Vut2SIOR89QjGfMqfFJ3OQ5CYEr4o
rJ++peFJSAhrBGehU2xN1Qs7xqV4Hzvdi3bNLgpym0eEKuqtgKUEpf0XwrvOs/bE
8lClRwF8i4AFt91fPghR7N05myqXGcmSn8ry2fsGXLDkCwZSKQ/Iqhd3J7B+AJex
to1zzfJGnt/Enh0TpuX5L0kQWi0xbWN3yZZlyeyEZw3BKtw1fmEjQ3C7AcgzgrIW
gXveG6qlbSCN231fGJhQ89up/O6tmPuRPzQxI3Ra6RHCCwUBnXD2fmSQW8lnpNa9
loYgqCuxP2S+AW0gUzqEBpYHaiLKp9ORbo3mCiCYVOauPD0IM97VGKliZsv+qXCX
UpeOVgIJTIS7jXbNH164RceXHuliWRIgBi8A/OyR+p7It4nLD55L/o/TDClcbjXP
ma01CXVH+dzZdadHkJssYQ5fSHxT7dkP18pogBA9jq3GKGieV1stwP4GrZ2cYvft
C2MFQhh4Jb4AN/dCK/fbuBRLV5T1FSMZDmyY5eDTnqWK/RJgy5WzQBI/lZ08zlZ0
xEj0kfvWCQdNDABCJozkB7dTDXgKM/d3f/IN0J0irmRn8bXjIyz0K/EdA7f8poUk
+ybr6QYJprQdauFTkX4AyMefxRZNdME0QxHePfgvBQQTbk4eK8qSOB4CcHzea8MA
dJhdGcI9HYE6ov6sc80AogIELw0dmNFk3oC2QyRQCgi2KHvlXSczxKm2badb2j71
Wt+TqYPat9G88PA0ZZHDIOdxtEI31yUtdIHKP5yjy+tm1oNL1m9DHieA8ERMUDwm
xvKxQzj6XAgwVI6alP8FwtkDptogjyTtTR44200q0ODcm7j2z02uKlZOuJ7m0MMW
Y2KYGtcRAZiw8BbdmVn//j8Nv5MaEhUvbNzvGBl4BihEZt8X/2lZ8GGGnTAbrZzR
ilfh9KGt33t6O/ZiYEOQIZuuSupQvKPP3tq78LQS5vz0QqYEJd7L/hd5gohPqvT3
PYIqruGxtmpeyS2PsvgUNSS6imudqGm7qjIA1ZGOLomKf8T14ksHR+8/um+BZaz9
skdbUnNPhCyQymNxwd6dVjVBTnuxVakLnGRQMCwzYutmrgu3u+QzIyF5ldlm7vyL
W8BYc4w7nKswgWmNUTyH83gFMAJmW+lOWa0hYccHnrFECbN780ZJVae6l97sliIr
feHO6BUtJ3nyHwQ6wXSEr5hINsNJTp2SFBRO0bJl08e21YNWC2syvIVGf8zhJIxU
0zhUf4jKtWrpFm7eMRW9QUitMbYqLdpli4mJQzkDCkoYjVcXPu3VnjW0eCEAQdR4
MHQOpcANMBpawO4cK9zNoP87IB7iSUzTKALja1+prFAZHGPBYnTicJJOB/E/FXGM
TUqpFCV/wYW/vtuM2pO60DvY/pUxzx6P8aLu6ZeRojGLwVZbnh9iLheSdI9UyLA8
fnpEXPtcAmF0XQzCko5mcgcOV78NE6hYkOCQlnpMfb9LeCJvydBwJGk8qtQyYBLG
b93yIk/qQ244wAOPTlcIlQXj/EyGfehXzGjb2A1km/i6I4qTlfG8mm36c+c/4SoP
w3mrGAkDDsb57zDXdm0mlK9C6o+zB1GN5fV8S/VtvfmiRNKJt6ALEX8+MdspZd95
wXlTATz6tXAtBTrDWeO8JCOcVxaWNa1moWdtrLpa9an2hkE6ABmXOGsolAc4kPJL
comKYG82Xmc4PfR/PikSzwqTLCMPsTMutdSyMGXtkLkvt0W1Irzt3BQBW+FyzSOS
7od9a/DWiV/Wz3gdNCIrB+hvUi41iYHxCjzbrXFvSwruTl7zvZ39DAWDNkpABx+Z
FDuSbVVnmndLFYo3biUI0xHT/LJyDYyV8ok5S0tNJ80+Q3CfeBDh38mTCSAka5i3
bhuTtoCbDxMF6lkI6tQrXqz0HtFdfJcQN4ozFRsF014uoRpBFKJYJZ1dLD+9ax+5
aMwBQkrvIu2IMkYIkS5+VqOQ38dM1wVQZy84/h0+dejGguzoacgy0GwmzqKOvSz/
VPNHZS67qiV7mAZdEIgNMkMSranhFHwKY/DCptpnRwac5Kdk/RiWBsp2cjHBm7bq
6TEEcgDkcbNetT9PkP1L7T+AXlQFzhjxPF470GhlhpoL1loLZjFxtkW/A2ftvSLr
uDIdJ5At9C5BDkByi0sw1NhDfjCW/q55w0XO2hZRAWakRY5rQGQ45YX2NlYv6jTx
koKDlvsiE48JzfXpv+T+UWBl8uM1juIcovv5pH4RQ4J7yJxt5kwIhOp9ax9rV8w3
SNCmi26Ot9g/bvat5GH+QD40EmFi3QSj5LazlC/TE2O/fqploCVEXcvkFNqbD/y6
xp+gLbNRFDX1YUgImI92fHdIYZsxFsHXEOwfUjr6/OquD/htSoIcaN5B/MqAg1Cd
VK6lz9EX9Ybg0V39YZvjn3r4jbuCeK4CW8BcrSKKlkE3Z6Q3Tg6PxAjZX5g3JKXR
dMCQat5knuVsUt/HbHVMYlvdrazNKgwA4jYbNaBGeGrnfXdb6S100zfyJuFECVVF
neEGgjA2badbJgtdRpVsc3PZJ5S18iyjKX1MlpR5yo+YugV+LAy0XhvWR8ElvU84
RM/X2cAYzxaloyW+YDvkT189eXGiIlhsLU6J1KVwOpU2PahvGDyGv2WrzThCTFlX
Cj8yxnaTVeFJ1habksp6ipNOGBaZUfysTB0wkxbPLyLtp1IpvZYBIZD+bcGjCJZq
Rkhx5tYveuhEIDOCbs9L2TctoSWIj8h6lM7NJRS9Fht0qimZq6A9WZxtHMSnOjRI
WkLvp71YcEM7uhDBuO/6N/aQQAZfGQaMoAyPYEQMmvkM4jn/vgNkUCILvsrJsP8B
RvScU45zemtIoE14wMCGEJijUHiN15xKurOLHEfAViQjIWc5dg/bMiXFi1gDqCbe
+68eCjgQv7oKK7MCqPYNqZRlRNmFAyCjWbKKP6VhHbO+ZNB5r6Q2MpzSRcjgSMBb
XgPDIkuV+XIJ8Z1+zPYY15rn73i8ii4TOROfoWb9s5F3N1g/8C5Tz15OnwqJHcU0
/q0wwCJL0V9/peDroYz/DaXuO7y+ou+CNaHSOO3oviXMOuf/eFJHcD07pSRcy3Mk
UI/Y09/aJLLXYmHo+EpRoFXU0CQQJtwJ3wMZJ15q+fieqx9Q1TNLkX3Q/3SW9R07
Q3pTDAYw53hP731H7la2i3KcvH7KTpWujif312bq6E3tRQqsBIQGBqc60vS96+Hu
exR2TOHqG0QPSOpApx3x0FzNX+Q1UIPx0WFRb5plIZTKpNYra/iUEGi4F3fcyWBU
msRrVvCMl5YcdokzdKO9Uuu5voAi1eeh36hDqiIowNQRrazRm04z2QvnDJhyyxWG
mj0Q/UfoqCVwcBIA9C1UqP2htCWkOcATIqSmAJIj33qPWsZvMY8R9KRAMsy3LqI+
4swm/tNODdvgJGMj6pWFL3vxun03DJEkrsQH4Bj4ZX6cWC4wSzWwCIYgaFu7liI+
orEd6jKrmd0W2XLN9bMB0M+GbbcoXGGI+Fc2UCD2uJ+oI54ZDF/3cdrSt5pPG1Xm
KynqZgwLrlmHVvE9yAQPx63S13OK3JalGnzrW1oDMNpvZKOgGqp8kBqQOKmNjP5F
fOTDtvrZ0vzIbkwSew05NZ5Yn/RzZywzJcCQzkmxdCqmWKq6MBEqMaTdIYsdnEbw
LlMAOnzre7+mzsKEZYjDTZiS2I8gzsfYRKzL3BOJ6rEIkal88A402WJUxdg6HsEX
LxwE1kDwKdV6bDiIcdpb2NBo3MLMk/Ihjbz8VnToZJ5Gh1tAGbvUy0sSJScQvGiM
02ZDODxjP25Qs/S09+jbRMEpU3pi8kLQg6+XYEIsL4/C085bttgrbl4U+zD1ke9m
E6vvPtAaH7YESHBXVlHVUHQOsy5Zq9uI14vPAeoV0TInfsnvs/Wk4vl+iInVd7EL
ETA3adtSBo9yMXQiZlSxB6hkwKaSXhwWzOehzzMtsfbHFwMWcEHhJFgJONBK9rX5
nSVVPHJrkXzOLaSIaonjyl/cBf17zFhdF6SfWIMKmuPY3VUNafKjRCHQtk09goWH
iIK/+REEhB+Q84funv+0G9+SFnd/FMK5zFcFeHRFv4onAMGvnghFEigb1+DZD6cD
Om35jSSezDXdS3SJo3YFeNGk05vJGohd7wBY2sojo0u9ldmh6A5n9GMpXfjHzlGA
vJ0ulNhS/g1y7X6STu+IIS94s8Himp7lNFiuq5uOKtd2F84BGnEAdKfnu/kBQDC7
Lziat3Sif2ZPkxEceLzhanMi/0Ph8DsBV03vjroHwpeuYwQ3/KBLyBUyJee0CvN3
Kyi+/aGm7NJPW41+NTI+ITYFgjr5hc108Qq6p6ibcrpu7PXerQCug83Isq0kdjbE
kzPDhxB3ZTmwOMkjp+bOeWUX9lyyAeo8iukDe4HDy37knpkRWbbYHryjvdKDZKOU
1S8gfPNnS4o0vGYsdsufm0XZWVHXPZ08rBMfqYWxz798tP0KDTZPn/rK8jUl2TT2
l7GWXOP+Nmr+QfIrq8xK9Ho/n4rlBX0qLmIDoDS+5apyyJH65NTrz4yo+rTmDMsu
W09jcjs/ac+/Ro7/m+mvoZvoyfANF1v54A8lFGFp0TRnFTl9sSZjM7736TUg88fj
Ro3CUWBnzqK1XXcI3BlblVucoR0jAv01hbFEcrgo90C1Ug8vDkSHIjap+xOv2pCq
21pLa1wnk0Rmu/IPjP2dXk/ItuIo4QxhMfvVkQjr7Yus1vsGiq7O2NoS+dK8WcZV
VJQtIG957ZOwOjPolWCOoBvXxiAjwL+GcDp+NLlyk920+hG+4Yn++f/LbkQuPVWX
Ihvky4IWUDtT5cPdStMs2YXKmMHB6aysDOCZ06whEDWqlo66HpUGwJHAMlbDUhV+
gzH1j7v+5+6RSeiXdLagBFuW+dAMwbi198oB6t4DHoaA9IvOUdA3uRPAtmtnwuNH
z/jU4o/Xjz6MkLpIRFiJ+fLpEjLhTXWpTr77GVLeCgZ5gaQY7buALP1afvJxDW/q
QYJWeZBXD4sP0eEp1YtutS37FJYboKrSiPDaOYVpBMAcQyQETEK9RYSFWC7noUP7
UuEHGCi94nsiZ3+OzkAwyQiLhxrydhwnJ9yI5KaZJzjejP/bZS8w9cryDLOYmeT2
mCkuGkRR4YtQcA0F3zwTZ1F1Xf/sUG92Ri4hAmLBGehU4/wnHnfzksaheiYcHNyc
GKs9DrPDC1zCBlUiLGXSc/jgqYy7XwbDHO/ZvjeWyZR9N7K0tlDuDED+M+KBb61P
8Q8BEuCZdoYm0FQ8B/zKUsFjCv11e/Z3EUAI5fnGi3nP9gch39TgVShkWo9kcF+E
1D6QNSv/S7ffBLrv2ltuIo1je8gaWl73QswE3DurnrGzbwU31yCoDzUGDqfJf72d
boo9QWd5NN+OqXCm2vtDkK56FDvbvz+K9Kyx7tnOQ/tKECmY0F3yTRTg8a+LwGKG
RhMRqJzBMdmMtdR5HDxF7cmgpKnmh+BHPnfgnO+ragQG+P1nG4Dv+b0MJNGRGhth
onXv6SkNuLlm0pVWJwNR+RHVZM34lStEFSJktEehrVw7W6KFh2F6wWlTvx6q1TMF
vmePvYMBzsF6ekAzhv+qHJrswPSWNDIK7YF9Kn/b/qa8qOYM++ohHax0M0hUz/T4
jNf8jSqxh+H7tDNEMPnBeA2n/x7gaF6moOboHARNqb/rBGbu6zCEGr56bHtPlxel
9yYHD708tCjZdQUCqoPNOr2hZYQLOu7yC/JJ+W12TVnh3dgmlM9hrS8QI7irY30u
LNzqglr5R84yeiDDfyzusXozqzX2veZEZNYxbGlbmVF3hQ2g2uv72ZmmCzowgODb
jIRwFtvxB7lLViYJi51Ky5gm0cAS6xrGbaEpokK2n0GUxB2NErUcO8UWFZOFLoaz
cFAcNG1ZhuzzlEHSjEKCEPFZxr3hqacwFx77PdDbnWIsClSZp5bFvcPm4d4M9hbL
dg1Mylq9e/qpo0VJDLvFdP5YPt5CGlrAttEskBkF3/KS7V4Uq2osYEmmxTdw5X4d
xh48NSePM3Dta79aUYZ+cepEzswHGkeYG0p+4ja8bnYqgLwIwka4B3QpQ04bxHBG
SSXkdWhqbAM6Jeh/Xz+Lyrhaz8jjSr6PZuApEMCwi12ZXDyiAZy3KXLt2WgCL+KC
aI6pe4y5KENBEQ4QGkBWdS4eUkOXVjLpZvz+7kbOV8qiZF+06VwJKlqJU7fagNg4
sXOziKIjKQWJteZ+2Z4DrCq0cQz4FYUwR/FG3kSe92GoQ4yCMwjvDXOKLBLqm0np
pxXAZlNZzC33+PIqp3OneP1toF5e8dL4FRUkifuqw+6MryRSSsSDMSTq67Z0mLym
NISPXvu9Vd5ZLbk71oE6Y8EY1M2EgAunkzkPPXStJte+AGMnVMC68d0Q8c2Pw0Y4
vazKBDteiW4hoodhYnBYNgBPNtGw8Vn+QQMtQYVIye6uyD1T5mDsALwgThdySn71
zN2vrF+ygMgICTMNz92wvFkjKx071zYLGkMKaytGsA+nWZ7aUyh27D2W82cHk6RR
wHcZSw6dSO3ENEhOgPGIK0Ci3lpb57mHUPkk+LIeIDm1sMeRqXW+3xhAdCM3+qXA
LdCLeaQHvmkXmoY9xzAe4G3qNmsWtWlUUSYTL9SI/IQt1/6v8tCPDIJLr1r/1Gfs
6ge+ebx9a08zNzBTMgP+zvrXMOzL41eqab7/7/nZNr6D73fkUf8CU3FNblSYzJ/C
xcVzd0IDPhXiJa/JnaOSAmTBBM1x3Qs4xVPO/BHyRvRL0Niy5xBqtkFhZrjLeP7H
pyt+7TBo7RczgbjXLjiPBd+NNK0f/U1sFJH14IDFLP9AtI+45yxf3j+Nx2JNBDp6
meZjCLdClmmywwIrA5gErQgKsd2gj5I6LNM9A4vY4Mn80Ub05GQA0DsLrDmIA4th
EOKqyDoMveOkLPlyamtM6bkEfEBLTF+mmbaUE3eTADIHVtIVnP9OaLqempdnUqRS
EKlKeehd1RTFl0aPiFuY/ZCvRxCxd/UnqhfKzJBcTe61IQOSqh8KrPmzGNuRFBde
GNWhI1Cp/oKtZXO/Iq5MMGmMOe9w3Cb1TuxcuREbmM8y+ojZTs3CSv7TdNRXmne6
zL47xhTLPp8zTloCI3YALVXZ5/E/d/EG4tlj39hXGvbGJfAqa74sbdEGWlcOV9dC
4O18KmepDydPss98qcIIo3tk2pWcIqkQB9cFkY86jzn/1ElwmVQOlICT8Y9eoWAl
HnJK70jxZ7ou+TA5sheGNyWlkXgEoS9ckDgAgU8ZPUr5Kzjs0TvgjT6b3qRQRFuC
YbYJmtZ8NkMwySrSVtMlbTrzYILW+YUtAOnk+DaoGZIWPuDIdjEvzMzBfus1MsTm
Do7BOVwSJzB/m4kWCNzEHEN/kGlDFsa/To1uAA0R7RgS7tw4MG09RTHHWVfj85FA
4MDx4/jG85WCR6oN5QB2aZ2EPCDseeSZ2cRDeq1l/CAUOo5ccFZBGZ0bcL37mEyd
MgQIqeeiKsJnLERUnhLFWZw8JHHqTObjpzvJn5yS7uE45/9JW0XvK6+OE1adzCsz
MUvnZjpVWQ986y/Xhll/Z2FnWpY41zyacJpykHQJO3uJtUAmBEvJheFdEw2fUawg
sylF6xYTOI6VEvRbUiKvxYXaXmT7xFuadnl6n0g1be0hq3w9lXpMBvPSDJog/5Bl
EmNR22AHOgxDgZE7D+lZPca8c0Dd+lXXqAuneyHtIFOGFWyY1Rigxe4zyAcGjtQX
q0Ffd5S6xShavW8ZNP/BiE74ONLEOtziu7U1bYc+es2Wxp+5fmNS25lGPH5zI75g
+lqoFgKwd9N31n3d48AvYLQCoBpIPpqdGafw3RJjTtIoi+eCnOwO+gmCHWk+DEdd
fNIeaE74dID045Ngpb9BahF62UXxAK7Ncw8OK2Xfzni5CHlNVAilW1xxEJm5yvjA
ihF0RmmEO7f2BgbsMiO5pJ4q6UBqfFmZC2s0NzXK8+Ik6hN5wEGXGDRQjkMhgDdy
TlU1UxwR+kFImmpwzgZ2dMxywIXy8u+ccGKSZ+5f6+60MeYHntMblYT+LHARRDtS
SbKDy2W/8OSPoemBGcrvtCh1+daXuDHBXEU1WFMOWrWTOXCrGWZaJElH1ffzD5K4
h6WiuVaupvBayB4ybE3PBayx+XNc+K0h7vrPivu5V/O+euybVxkoY6AYVVJpTeL7
WhedvzqcuKbGDsiLmd2BnCQPRQWLsNuk/3qeTvvhJlvCKC9IJYgHzBDPjqB/GmuJ
xuLgYbNYeQUGvA27jpSzLoyvfomkPpDxRB51h6EqFyCq+HiTb+sCRGMtHBmm8O6g
y7LqHD9ALdi8VI0ZFplEF+6U82yxwY0GwnuovTHKsIMFndFsadMQijqJUKwPqW01
n1HxrSwC6yYrP9og5aRNX71NHeMb1+qOUar82qq027TFVZJivbMkWlYwT47vFMkN
lQu7HIAPez8KfbL4xhDN1UhdkgsJXjdQWkTedaWlPSZa2TlZxqa8iPBXpFkOeTOu
h3e6BEWk/MdkLPb15/mYyZwgeA1Iixbe4oph/UozGt+gGo/btyv4b+aT9dXhuF3f
/gOT8PHUEuMzZL1vP6zaYVY8nAaI26cwcaUiua2GJus9Vn+rqI9Gd/8ZkquJk4kR
k4odX17NWmqB6aafJ1MI7nij65z2XH5QKeuzcvVl0DluIJLUfnxl8VumrjLF32/5
d+S8ZbXurdjGr+8OIAoyIfbSWHlf7/1mUVPyP2O8R/ujE7AM7szoQKI0pEomDgS+
t6y3qgUeEOx1qhsSvuP8TsbvUpbfmW+ER2v+eI9NlbrAWYzrIPMdVXvMoCudcP94
5zwxKcnJHywZew8apRoYo/Q6v6xl6OF5qiXCe/4Mf1xjhwfIZzpi7u5RxZTv+Ada
wd+DEjwf42RnnhfP221PEa+8xdaYb/vxyM66zV7jUU+qbmvbCi/FQPEA0I140g7O
ZIppYZRV+kQVx69X0UivuTQPceXJO2eTT1y2ai33TWSb8KWWNSIHFQ8FwOsLKMIT
NFHzCWzx+JTZHmelH7L6kPTqmRhzk0Q4/IGzUu0ZIWgNv3giUN437OtNEX2/Bzai
OBftk9Dn7WDRV0rIQ+CGncfzizJ0tqtERdSVat1jSTxT2SyFRYbq0sL3e5vWj/uN
n8ixHHjPdNgJ71KOxu3v+4NBtk6RcewwmHJ9l+C42PsEkGBJYfW7pGTvsaLIeVeT
dy8syPyBDelQsJh94tKfq34TK3H1HIZgmGfvFetveNwP5vkz1GP6KOI/X+H+jpHg
NTuy77BKO7Gx8BP6/L/HulZQeCnLNhpQz18GUfQfZE02XVqa7BBMRoZhB4hRIqQ7
Nx8SubkWktuErzAjawuUYqWbv489dWAf6hWuMQm105gNFk1/YV0QSv7bviLnb+K/
AOQO23oGZMZM4ByoX4UA0vpUVZG0U3nu0kOYMGEk2SZj5/H8o/L1CA5i0uCU45tk
w6EkcADwe1S38yoKfoP/XyP7HPoJf5K1qMvHCwJWdXQeZU53iMDTRUEs58NCXzjd
R3Yvn1+pY9GP3FM8VjNDVBgFlrwxhHKV6p76x50fBa+ojyhpSFquq0PkOq8p85cr
bLeLn/qqrz+m1qr4xopd2s+5I87WEENHRlTm1ZGp+lzHBUkercwu6UQPro8vx7Fv
Hw9nDNPWtLmXRf+2r+DSxxTsKOqy4t/Z/t+ZqkoqDpIYVY/BexAz2MJr1D1Iw0XJ
+qvZgI8GWnD+xvmpeGaSZGYKuyBIfxhkGNF3EikgC0Eo8waldjxRYeR3ZycWCwxt
gb8433THW82w+qIpcIo9fmNAm/sKDaP9VOaXyJMJ14XUsbuuxFThO0ClLaagEg4D
qFjxuQU9AUXTJtrFdsWtZpLmRyPDMdwnOzMqL9KEItUbpY7J93iQUZnqcJrp+6ER
KPeH+FxhWKCh7NPTCr/TmyllWeFWkegESMYkAEoNgj5VufdfoFWrfSqaBDmt+9Sv
Q5DuRRGvqVSiCzzaRJ2aZLqVOrrrE8hmzEXWN+vCguomV1B4d9gdNT+XZ9WGZ4uQ
gTyJH+EJ9juyEN0zAidc9ojfO6CQd1ODKyffSKJZJNjpTlK+i43H1O+jI2i65Elg
yAkqiLFTLUkFSdWtXVQv7BhEe8GF1kAMHImYjuaB5miyJah7ODfu+lZaXETuhZkH
ha9rZkaWnOWdjgKKwEfEwc01nZoTpJ/cFqWzSqm8KWlS/9bDMg6nFc+ErIxnD07X
6A3RknKBsokKpLFnOHnwxU3kuoG+RG2GuIJ7gCyJ0NXHx/S8vLhV01/AxpSX2gqz
aUeNyrSlQKFWu3bkjAd7nEU6fWfS5HiGxmp3QJMGCQiV17E2QxtviIgkAXGvCV3L
kFHofHXbatx5SQt1mFkFq4Z8kVt0R24w4/GNQJAEmJVuFBEJ9L9oeD9CRHn9l39m
T5xnsTNBPnm+0audlu5YgNrXYU3WjKnVbxreFhucrq8j7HB+zZGB2wPLuxE4gtsH
T7r/C20AAym+znbtHCdUJPRGJn+QDB4GV8ytfGYTPyAAwiQ87Yt72ggjvqcuZwXy
vvBcrludjtr1YvtVvrt43X7ulURas5jzpDQH+bKoGcc8m/MHHuiYv5Dbe7KDzU2i
5UfMahZd46dU6mO+WKA3XGKNJOePXfUeDmwJ1xV/wMh5ufRxOjnOlRaBlmRNiJRL
+XlQCISczcfnh2OPuUtU0Rmhn+ehLb/RtNMEIutXv3Q1Qk/vD/HU5iF/CYCT8HHA
Wk/zRXg6YlxhR2rQw2MJ8B5qFi1mjkePZ3WXO/q7tSq4kN4CL2Eb7JQvPNX9ixub
pLBulvY99fJ82o21DBE5O0hXtouT6ay6BJg5EuNjuO76k4pIWtR7e9SLLn7cN4aO
adZ6O9PKoatzlFj+SSH5ybLT8ZHkY5xEWeClR6/du7YbHtiMA0djynBt42ZBVXPh
f6AgexRe5H9UOGkXuxIPxk5ybMBKvVs9HYGIsFJbxKVXcAIK8nv6BnFaY1EyMIxo
jWRitHDEhVMEW6H53PCqOj1sAH9RXYeGLb9ZpdBXuJf/vcEI1g/0CDZUsHeP/ZVq
pdyzTvk+Bc786N/hjQZ4CMHTZ4ul+Vd2GjtaRcE+xpSq3NwQG36BaAN0kme9UXI4
U/BdqUlyhulx8gilIjeqFFTWnCz/FQ7ZMdk0Es5PzZGuZVVHNKGGAV5zb96aXHwU
r3wF3c5rOt+4wgfqNGejRLDjZYq5z0E6pAJ71VsnwdpZFS5AwkjHLopSWjc602ea
9qhY/jMJmcc1KXsY1Q8/xJ6E4VrOVUChIf2uV078pZbMV1Aw4mmETk1esdmf+Oq+
9sOrZMh//TtxHB+PM0gkSFAyWwqUvXx8+DGgEcK6/KEXYZzrCUA3IzrHD5lXrfX7
V8lqMeGXNg2XJoSjuHipnL3PpXIYdswSTEd8N5Qy1G7wTogdM+XFMsL8tR+Z9UUG
6wK1I/PSo4J7kREOcAj2mTyJT3+ADRBhODegfUKfiIDkAAtZIDgCxZEy3nq1XalG
KCoOOfiepyY0sN0/xyRZaq/nciK1O42svo7QDAkMN5sBQJn3LE+QTOYRGlB9wEpC
cK5tLW4aERHnSZxKSFQ5KxIN+LP5krxnAeyCbekb94m02smQCIBhncWUlXXw0rYA
hIcEzAl5lkqVKFC/J/BwmCa48NYahxpXeORWvBYuxnCLGwORyhMqW20TrzCXLWBn
mpa9K1N/M0hX9wgRA7/yh2m3Z2cuXTmgZ+S/Em4rvU+lXiUL8Nn6vcicJOx5xsbt
Jepwi/Gzthil2lQ/cw+hXkjRCUV5PrzOrjkswzWK+wdQH1npr3JsGv0DnoiAjTP1
MKoykB5gh5/a9OCvkl3GjczMDYxxg05k5g2vy/WXdKE4LtXpOxi5UqvH4D7FK04F
GD/1bkAOqBfk3X+19k2UVwKqg2uYmVTaiR9EWOH9PcIBNyVrPk6qcKdaegU3nNMV
tJzCcKCo6S7BujMQ9LZ7bToF0Ls2v7paLSEW+fwDhlOd81vCEKwdLYyP64RBDlux
t7g+4/jQjlF+seKxCe6kpf7fuFJ3H2nGRCjtQ6+vOEfEcyT6PSFH9Sna0QvbxAmI
DDj+0rlDmv9/K/mREaEKepfKnPK15gfR+Np9IjcXxfelkjURSAbwxkfWZJR3pRTJ
YmlBcQ+bl4WVMUjZ9YNEA8m4MKRni5m9AxAx3NxMBE0TNI9UEJmzoi/IL0r4R9uy
3lke0h8jV7qOtn0oiwkMX/doki/Udm7/O2rYSd+h4Vz/9dRqe9Tw9c585YbK+lz4
yWUDGiu5/M2x9dKwJC7vPZgrHPjarDhXogzs3KkTdZSnD0I4GMI80IDLjxY9zEBE
ecN4eQnZSXk9mVzL63nRfen6bIcc+EAKbqhYEiCFgB0b4qhsVaPVssZFyRMdX2C/
JScqkQPERRRmopdIw4YgkJJqfNhC548RG69SWP9EQBGt+7Q8ubt2XmaEQTrOO3ki
lAySb9VChUH32DAknbeZ0gQZ+bf1aVjc9NAQ/TtggKjUvNitQsgyE8hXvAY2VuEx
l3sPM704OHoJRlLjhWU5ECjYFHSRbBtUSVWw7+lSQ4lssxhqHM0cTpO2O/C6bNsM
aAB/1VMKyGlxGsbrdam1LzhAnJzTJbMQbb3NFlpGHHIs8SALzj46l4GNeJJqeRes
03tHv6Zsoq60MGEB6V2THs1WtWCpWdvjpVS56jt+hCoAk6r8dZ5zVvO0nOm/Ilx8
UPToaJvTkwjGcmcnhzi4WScQj4CkMurAg0gAoP6K2rlz2nK4IK7wYzAesuB+NlCb
n+epHTVs20MD/AjKjLdAsz8c8zVV7pkqLsimzDmqBqHDOyHLeWFqzn/7mPlyh5m/
Zu4Oaf9En68FcJVqs2UYxkT+6fK6oBGsN4lxkOLJyr6BmaIKyvG4EhtEi8wMQ0yf
ODHFqoakli588rDct+/ne+lLmF/0iONfSdRDaf4YeZcM6gF4kCgFd7fkCh7Pquf8
8Dq9aM1hjgvLutjTiPOmDFB32zRsM+DxPIpEJrBAtHbaw7xlZnuLyJreGJuqfEFL
KX8fDKH6+efV77CzvOGhgXdrb2ScPusIlU6InGNYHfXW472HQ9MYGN1TqsYNmQ+s
7eVD9MFZKtFpWb1jsZNU0S1EICN9V2sIumz8V5WIWjBqYpeH7iNJX/1Z150Y9t68
JyrNdC4Pu8k0NOt7aKbpLk3xVBce89w1WlEC6YHvV45bVaBDfdsSwMqi5dlsIcsy
Ng2MRUZaEmaZrag9Gl7Ds6IfamCLXYqXMR8/95si9A+mqDtHjiNkTOlHJNglm0AS
P5NRFlIGx4h+qpcH42Ls/wmVrH6Yuwu3WmqZQSQXug2LCD6upzJzv5dGW+Fn+nFN
kyxfthn7VSqVDXbt8s+K3dfLdEyKIE9AGpynAlIYtseHL3iJYfsgiYvWZWf9kprj
ieX8HTAr3xSrs5h6jN5eVviDtKkarzJ4I4sDipguVlf+L0WX+jmkl2Dtda2btR1L
cd8Ww5b7PnB6trPRJ1BFoWEQQjxO2DpkW9rIkdpNHASN+5UCq6YC2VsjRKE5tYrq
Msat3f5cczEwj0OZ6soeZfu1zmkLgozDl3qcWMnM0+3zPuQKSXodOA4JbDHfafMA
qQO5O5Ny8ZsCnmiwLnM/95dJvztW12UfymVefJ02WEXwFGrBjjn4J6wW4jtNIXur
+3ZDxYzip3rnJdUuxAmDACR9Dx6EZF248TwLz7Eb05whwVG/4znV0s9MjknAjT8t
/EXz1ZI1YZUhfb8ReIbRDrKAKKj4GLE8o/q/ksXSrfyIoLbb6AiBZ/Zq6eujwEyl
C1LBiRs4/aw81ZIdQZj0Dy8WtEznHfjm6lNLOpq0xu2oBrb3pRmsSlSG0OVNv14G
+6Inch7JUawRaaWcaoDpVrxvdu+ys7XQAghsswQrNCU2h1n7NfdyRsPGiYBluQTV
nMNlpA1qVsxrRREi7KoX95B+dclpk/v1hIJwRHejnXayIXVSajK1pqJ43c0Tewvh
z+8DY4lVbY/Zr2+nDG1sUZeV25xxNivsKlUTuYdNEzrupbdM/kTLKFnb224pcnG4
KkbqhcfXKrOleQ9PAgTOkH6iLc4FKkYvlmLQk8eqWstzBYszx5Y0rl8t0BokIdhA
fl6G8gdeyNEFLXC867OR4fAISd2yFY/b0zPy8EmKDaAuSiVrYsLRTfxEsEMaqz+h
57K8dewwROnZ5KKB9zS5v0lFkwwvWsRkfVqvSuCzXSE6MesAqyjDFzeeLzzSik6q
ShqUuu/aeHfCsWta0M1pPyENBrE9rELpuJkXz2QJozWQWiyBj+ZYZ1ulfRU+q6CV
NcUSP7TUV3CJy+rgalabgc2u69lp9fW9FD28tU8r5wyHmcCmtS5P3PwgRGcp8m2k
/GSU8qGqsfkwS/c1Hy2gcsV0A2wQ0knmwykOAl5sLalkKufHIr9OKjisVzk/gD3H
1tr8ubVF9oLw+nBLMWzLTVYV9NUMOaexezcI0l22V787EuFcp0S94yod2Gr1nf75
sTyqtMhzdJvahp5tl9LrqAILe5r9NnzzT3m35NKj/LcUrosLMsHg4bpaJdibIMHL
RKw2RU944ZmXXqBu4/ljfdIz4E5nXxdsmxQ6y2zwVMkr6Z32MfJlVAoZHxIl78uS
UJagBaiGtMBZ98Zu7oJgucoFpWORMImUvWXHQHI13hbR2RR+ovoyYk4cIeCE4vof
dKdkEMjKMsHAaxuUjBeoZxFSZgw5CZPX7TXPXm/JeEGoOVo0YNWdcG6k9oaCNDxg
qOIBrUXCLYh9dIKNHL7mQPg1mY4k4NMpgaHm2nUxGQJ3tp5U9Pf/a681lEsLFjjY
wcX3EC1i2apZM6hZtFHe7Y8+7UFRB45cO5Sc3KBsywy89TJLc7R+GFxJxz86w9AJ
HO6x3FH3o7kWhOBbV/P3MOpDlcRt8ay87ygAC2Q4dRz/fVs6qDNx2y0erJdlTyDZ
//xJOMfNv4B0DHHwOt7RerCglJ+jJXl95+jdsc1SUwy206LzG/OxmsvHpBwMC9jI
rsvLkALmX2igUlkB7ybw8TxMWnJFRK+zPgYhoxC+SKgAr2cBYNS3QCavlqQgliiU
jeYhvXVI8sLV8oxiXGaWbJe+fX3KSbzrjV3DDCH6Y3zoyu/RbAj2YP+G0vJOHOjZ
GZBZZxcNwdF6YSA0Kem180gpaGBMVWYfLabyIScQMylCC99X/gcR4v/zC04sCMwW
vlxC1w1nTYqKYGD5oM6Kfunjf/mTf1V6Wp4IfliT1bwVl6M6DCOr7vJLj82+yCLq
7hG4aaRbrPm1BQW5fG1XabWlHWo09/wdyoQV8B83JW6HbROP1pU3D7CI8d/MIwMx
ugsiuCY6VPDbw3wPU2ITsgpa0U5UmB9zKcloZDRdIsYR3J1jEtSrz7wevxyrkPKn
T1Ma0Y2yq1W/0c0YKqLCBGlvEn95N0jL19CxD9pRPl/IkJRxGJIHuafO9NIMmg3x
yCvnzqmS1oxdwVM8mDxKEhB53rmDndYjT82WTr9vPvOAMW9chEdRgvAkcM/hZkeX
YztrHtQFU87M/r89K26jkvFQ7G8Z13tp/Sdv7U56fdOX+f0GP+TyGwSoZvH0Btri
JgbRiqFBT69XseB8+ZjW5N38JsxlTWjfmZcI+t/VA/aRhF60TSZkwO+ufxQXMR1n
D2wVpyOkKAUk/xWhKfUZGyhSjDkSZ6tvvoxrosOTGz2IpPA/6oIDg+QS0OK/yyE2
yWZrZSqq9vAmfwZmG3LFQQMbDnL45gskyRtboW1lQyxENEwpZTXnSAAf71vdnmhQ
kfW8eo7/vSnONbd4C8ICXeaiBvqaszpdZteMpkYpxE/t5n52JsirTtC9TeFEBdL0
mL+Q8QW2Um4nt311rH/GjsyVJStC3iB+ni5+178rL2Kt++TyUhre0rzX6WSM44NU
xkzWDrMw7SwXTA45MP1Rih8xc+gB7a8Zgb8uphDYkRiFz2QJ54FoyOHxqD12h/KC
YNOkeDhO4Fg2SLgC1zbaaBXsW9VPLkqHA3qJLo+r6KqqinCZgdLCRYEl3IE65ZPo
ZNoFDNwy+UuszLZC7nG7PxYsuSsAAm0PUg24OnBJDGBJcIWU4eZ60t/+CaDNlllQ
zUnNsJ1uqs2ezz3lnPjpKTFPYKpjj/G9Gu8og6B4XhQ7cFIQMeefYYcZXP4S9RUY
AeRsgWsa6N84DoFtOTIqOLcrG8dmxKVdiEMwU5zvLGF/37hIjcUpO3ekKhSkm9oL
gzaQN4vCIU5a3q9MGh8oiCsTUB/E1QpIKw+8zKVQYRfyRF9bMpPTOTBrOfKvo7bS
/8ZY9G+Ar+cNv8TeZhAHpXufeSfzwZe1o9GMyEZIEgV+TNhPk+S0vn6bjs3hQJWV
+P6j532GukQ3zbX7pkU0vX6MK7EZ9ucKOmh7d8QlDvnaZO9S9HJtE8JLd6L4yZhz
i2dWQFknslKoQFiyp+OkQa6XV4leZXlQ0u3YrFj5pBhrln5XlKKOcaYT9lfTPJ8z
HNkcQ1HtLXPQ+/WHUAgrSCbC5/62iQN1r1qDwo7q838Oav7THvmvYu9SGe97Yd7P
TwJqj36ghRE8Hhs1RBEM3p3mbk46QXJ/9hnYiQfSvDi2avx7EAGL0lrRj6L6CCH6
fVnxcckHFb+v+zUZl7sYbfscGoBxTYcngZA2GW1hm9vk4jVmpG1KQZ4bKk2rIX0D
auVfBgle9ioozVH8fjN3bL+oDsZqqrEqMR/YNQtcuojY5ZrEK20L4FAHSyNsAk2a
E3CpnLv0YN8y9G+5OBHwqHyCdXhv/5Tt1Xa1OWWy9E5Vg9kCucEyv8eAY+jqESEd
dDzGjmZC4ZS7m0bA4Rd54DAMYSkhIVV7fPWf/q9aApHlwjhdwpH/UAOIYpf6OHT6
twP1UkOF9zLT2i1uXGMCn13KemyZ5jakeNCdUH++RIDewSnVvXqs3s2xQ645rDEV
BdgmVBu/lQT4LSkCh5stskr5R/F0Kyfq7K/gOg2i5C1AQq4SBWMYFaU2eZ4ww3fj
2Vg34rHpSiJudGum+h1PFgUt5fOC6Tc3FBdc4l7UGY6Ekzs1L6acDkac9c9MPmXs
zSDb6gOdSiPLTGHxthgiUM+vXsaPrRdFak3hnAsshs41y2BEuTEfiIByje4rvJaW
Qf1EQ1JzMo0aelhrHigki837IILnXwfU5Ljq1yo6Pf1Lf8ryKDVIRgTOF8I9XYV+
JAZx/hquX5ZDdp3yH7DGEJ8xdh2mw6/Bd3ErQoUVnh82VrTkwmZQsO8aq+/3jK43
LEezc2cZJmvvHQnwzoK3t4Zj5EDEwVM6b4JCjRbUie2rn4RsbWs0QUc/CM2gGXX/
TT24/EsjHILHeNf6W2bjY8BHCaisNzpENVP3y49npFxLSbkRJRuQmv7sYdTkzu/E
gszu3vV6j9THc0YsVBHivGE6EhzRovcgmGMq9JesGx+mcI8YKGLSPQp8D50x4tuJ
+MugxsKpD0J8t20glnxcqs3RDM6g0DzDSJ9ySAT7xr6yZmPi2NjYllHknTyYB/iK
05BWFnmiRE26zwxBsvnPk8vkwP6iOMTUgoxs84wDLxDB/SrSu/ECyGwOVfZwKmgU
kDfGxNm7g6GNIR8Wo/fiv0NlK+T7lL90oSFsL7Yn84+mDJ2v8Fc7JCAOwyS0a9UY
lRcMQ8noLriF0QjMWZyWS19NtFVSi3KAj/M77Ml9bqnmSVLhKclEmDXd4EivhvyW
Btg9aChCHsRVUJzU72Zh0QJflIgGTvR8C9HLb4mZFvNAY55k+suMiGS3Rsobrkuh
ikvfPXhJQPbX1AClCUK8w8ZqpUPTUfiRLfgA84EBfZZQ3H73u8Fnr/wE9tdsa5mO
WupThjBT6A0nNs2o3JlM8WbvUegKD2AfQHahCKmRIuoc3fIXkQN6poaa9bU/Yd6G
51IWMu4TCHP5hXXYClRUtzQC5nF7g1VClSxrDkSPAwFlV0xGyNh6M/OXk2ujkm7S
EI/t+53snpdw4sKqWB0SZorI90Gm3X6U27PuiHyHad2WhXRl8PhC2v+MBmwxhphV
dxHh49AvGLz+fesEZR+2SZi6Gksa5bj4k4g4LnXBJ8Qg2oNfhnfZwSERuIqpmdes
XdG6gX5sJ4WrnXhP1wgKEoS9FTnvqGysZgKb8pZksSdw0a4crI0gh6TKBgzlNNvG
Mwt+d4+1fZCPxwqKRv1SiBWW2hu2D0ALlCileF7xXrzIjc2s7Sr7BQj3FlRIFSwE
ASDhZAyf9SCKURStZcix6pYctH5dyD8sPPfkPBj1gx/t9ePRw3JzQdc0yXpoQVUq
4GkIk2JAwOXMgcLQ9e1Vs22ywGPfn2j8Bfm1zPsO3AGEUpQOjlLv3sqLX91oFz1b
QdAqIu4ovSj6S3FqtgkdXKPKHrWos96WU+Wa3Uhq7hQ1LLqXr7uW7Qm/0f0rBX6R
BACbkic6UNoVEU0lUY7iyyNmhWpiF/+hn4XrFAtKmi1erFRVi4Pl9k4wveukSakt
6Av+G+o0NnjUzJm8JUYv8TjlyeHj938bgy3yDbuY7CAzfJQuwdWd4gW2TidMY20U
rFCkFDVB/lQrGdt2WFkTyfxj48ePgy0FjK1Y29ZzcUymkNl+dJT2+rRa17qtixxx
CYPs4WhpAch795CfYNb38/J90HsRbVuPjwj23ODFWSVHTIFKrcxBnVrY2YQV3/CF
YhjaiMOvlyWc6MDblLQczAyJIv+NhEB/U0gPYcuVHulyu+N4uf6pRRjm6sYgB7ia
53dqcWfcPpy8NOOQg2ebtr/6xIU8iDXHdz0ZLpGZDNGhRu7THrrmCVhWQyPbBnIh
LIVhQSYXMh/MJRj2jvV5Nb8nmPo3Y1kbI39SWopZMKTuvvZhuP04IiobW76+GCog
VIadYgaCs+QyrbOgtQPaPKmm4CtHEw93hOMO6RVV/xp2R/pQtq1jsA2RcKHR3EzU
cfEuYeQQ/7wifQKTOMbebwqdviLZpSFDG22ULNVuZ+YZ8CTzHZBUQ4Xy2bYHLGNo
RyMIi7pvPbZa+XW85kRttmyuxmfyreg56B4D9d0X73iRO2yIUX8Fapwwtko47lcm
Bh9a87853fLDfxtuCQMPJEAghdw65Q6lorc381fUqG1G80FVkCRSavk7f5QJfHjl
t4/ZIhMvzukfHoqUPkWV5njq/tYE4A72V8I+LLLVFE4McqCFKFu9QqqReOYBG3oJ
DTuN+6fdDP3U65AYnglTDmwrUeTmsvZ1fc3n/TTqMgAuDvhIfjcDCQprzRRq7oeG
pVN1GNxjvxU+5KreAVvGC2evp3lzhRT9vH/Im5mykyfT7V/hdAqVEVHLqhno85OV
9Ugz68c3v8ISq2i9rqS5vO68DiCmzsuSYzGUQjOqcI9Eqydef0wPOQaavCL+JRa0
Uu4FxziHIB6NTGS5bCbVJEO5u6KeJJ+W42F1YlI5ewz6Ny1Plo3/IzU4fHTjRzxJ
B2UqDQw16I8/pWFPp9nUTAszV4kZFx8MhlRsoclOlptLOEEsUT3brf4I1VhBQxxu
kZ2owQECvuXEj5iweuS9xKU8/+wTdNWCZA+tPQ9QJRB1QbqCwlPEKfXF1Y5rOrCf
MXpWl1EFdSLVLTR4w5C845AUmET/MpkwQMuD+E2cFOPujtgR4vfwjF7MpjHGX3/w
WiZrPq2aPVWC6IlTKDOOHC39WGE2sn4mlaFNx4EDKVb6V2p0bNLekhwmNaAVqDaF
430Od6ej++QeZUry5Ac0a2JpHqwMOmiemUBQx5bkcqQgQHvdonFx3VVKcYXy4zIp
HMTVrV7rW0qi2ToeivGayTFu5Vbdu5PmfGPiolQmIqLfUsTD4ZxE+6fMMrN55K7R
BLwqK7k22baQ5FzIbPe/MuQo3MC0s7iDVotki+HPvM3Z7JojJTWxxVpWa62cI5Jd
z+3YKn01INigyFS6NEF/nkXfO6l3nTsu94WOPCDCjkO0TGrUr4c08IQMto/rz1dN
2pVYmf8oDVbOYc01IV2zv4a625wN1Rh7fcnVdIbcwwSbXD4lqpSsP7El7gYEyQRS
sZYe5LyyZsFCQ5Uv2scggt7nQS6Cp7dbc5akKFalyPAm8J3WVui4o7+ei1zVnPL+
ax7vVUE9VqRXQbs1w4vZYbITk5bW6AbaX08Q4bOjBjkR/C0jYzrwRSzlwX/CXuYX
D/enUzPcjNi8iNdJUyMql1tpOm4rq5jVKoZBQYs0YXknaFHK1BQNEH9jEU7VP+44
6+3+VTbJi8effyE4P4xkNL00CofRvGSbcni1kaMWOfkz5zyBfB59ctdwEPWfujcg
gu6OiDxNwV/ST6es8RUM7qGakyBX6LkwC7i0CA5kuCkDir0gOEsiXVtmLxBkFQUL
T/ufI6Xgvf39SmRSd5XnDZtnZE6z3bqcCUPOciIaA6IcA9qFiYj/SLV0qBkupvjU
tmu7xce3XMiCWtJj2F9jjX3zTPNH5dt5bW1i6iHknq5WINCkwrVCfr4tNL8rHVgW
XPznWj0Zcmjqn65x6KwDWOjNR+BDmATWTakha573q12mMFqFRnIeCBGXzYnWpsTT
oaqpv2yHoSqBWlQ4T7MtcfniZ8gqa60I9Sq0Zto+jmbb2mpMuY6zsb8gkD69IOHE
7h9YRH+LwW+RjCu2kBqEDPx8WRgko/2y+mLBoyRuYGjX4SHl4JyH8A9nizGkPeqe
6yTNSSbSZ9ARsR7HRqku5BNAjzqVRLTC/AE7hxjlUQupSGO98piZ8Fw8zN5jKyEd
x6jUrGh7E1mxdlKQ/gmG0LuEwr7amVUPyERWDUQdvpyxOJPmE8RDD6/vgicxqWzE
U+fsWnsc8i076+EX9Srs4BibdoossvFPuXnPXnHxj+BjaFCcJtx+upqhBmgnciqN
oGDHhJi3rzQotTFByWeCbZm6gKYJSDp1R4uvVqnJ0ru0K2vmQ82aUvz9LjLwTSPA
inpTvkO8Y6HdRcN9DQ00/P2CApu6JNiKVTyrWaqI6C91l25Pitl4eKia0ft9vofc
g3HyZKYTfRVreLQqj8eR31cI9S9OTVneHLIfte5stU1ljfx6YjQwiFOz7Licszdn
+HtqD2FBWk44W3FA8wRskCckLpXJAFp4ndBw+rmNGnRevdWvMosEXDc44UMmwo55
RhF9JrPTEdogq2LS/myUJmSqtW6RgBul9dG/BuRSmfZPWEErILsW4YNcn3NjKrey
ansfSF55dRqUJQNQnnPJa68HyVF36W5xe/snAi6a8ucutosLaE5UrzzCEHFeUILn
dVIC/cY+Ex6lBgf6MhKdWCstKPSxvcCVvrBsO/oG+j1QWV/P14s/oNoHHjsKTBSB
LXQ3peHCfvg76n0KDIUXGlRDpq73AlhqbN9iO34wdTSrdE5V1DXeroz6tIE6eg0z
DFMtKgGbWeJXgGeEmHsgg167Ibr4+dlNOe7dtBXQ8tOvYxxGWYFaScYjEJVvdOtX
9FuuK93xMU9kRS1PRntHfggEfLm9jwGctQu7pzek1yCrDyq4ecoeIsAWhC+nmVe4
iXezyu//ATQh3iNdVKBEnLSkuxZUJ4ipX0A6MSzxb2IXPCI4JVgPCqrDu5zLohgj
GocuihARil23M4gQQU/G3GsJFp543sQ9S04mVVP9nBqXtfSygV8BiHFgel3Oz9YT
a/kFPqEzpBNP11px4MrkL1xh+9CJsQcJjTZOuMx+UsA8aasQLtmte8nmhIAaxZKn
jsZIhnfeZazVbj1h7h1GQpa5jwuoMEiYkAeaz9Y57g50H9ZDHAe1x3MKKPnJd2Qu
XOe24yK5ijJONbaq80bGUicDUSGd5Zc62naN1YY1DPQwmBdinSJWP6sAokcNL4V5
9HfHC5sVPqubfO7Dl3hnbxxVSNmNgjj0sUeDRcOOmWYeBxJIN0OFQttiaJzjqbxG
Bt6uecfz/e+LbCbxugOhQMYYuekhorN3lD+plZRqLpQoTlri4uFHZqINAEupZnxe
FOdgzr25GDVwOBJT6z42BBjRAsIlK5lbbez9ey0uT1uuad7XuZXYDWDpYNxf6W+w
ZuWcasRBHXRwiCYDXVJ48CmSiqys3ujDGksVbeG0loCF9W1kG0ZBbknxFG7v3toy
j6X2HpNAW9iI+n6mLexafwPCp5+wtQX3TYOKXge49cNpMOMKx+AAQdmBPjwjF8Bk
TUtGLgeI4B/s/4RVJhAG2vAyKuElwHtrjVT+yGLqQj9RSrs9gxTmWYO6c04j3QHo
Us4cyJf0agtZXynwTPaILYVNIo/Zi5M7XWJpVtofuGbBdgwaYZ0gB1v4t3eOQtG3
AH5H6/nRALsF/1ygxgoqr7Wt2Wf1oZOtGqjJT43LuSfg/EoTM6QmfcwyZjqZxyqb
VJ3M/XBTzufR3OZYj6EnO4lgGv6nRDylR546xIYbX01QRLM+CU9B+eUCYTuqtU0c
LmPu9YETyb9Bq3DDaZ3+TcQrvy+acyOmHyHaezIsBgAGo6+Ak3EjXVLXirGsag9l
LNHOEbhLmRevlL0a7M2ljG73SupcU0V2hqQ4ZPfgwsWajgSCodQnol8DJtE2lFhY
7dKsy//3BVs7SGs0T/+75LbfHxlFTiKwVJXzOnTm/VDkfI2HXh2vmE2OEwsHpVv6
A6FzUV3cUcenXl3sAsuUsFKhF7nKYmCojnQLY7OCEvZokYVGwNJBO6C9csvgBywx
M3kIfKhkwvaa271tRzzhl5ABSrbWBwqZJuloI9sWCdah53bQQuawxhIvFNKFVLZx
tmmy6S9j2YO8i8zNMWHRLFTK+43nJy1YWtpOIhn7G/j958nYGLh5Wz9d4Ho7SPD8
J0v/uHvqP9m7P2oVEGXVwK3wpTaW/J19f7kXqYbvNdxN+D/oXiGNnkjl3PbZM9so
58jbG2ErUDWwstVBYJ+dV7HTR8gvsR/oequLDWaglhs28SZBm8UUI9WP+1xtcAV8
tUJTE1fFhe/97baG0sWXOCITfH9qLgMkuKJnMwU/ZNL9sP1udfdlYPKEPhZ9hoV9
g/KS83IRVg50AqfaqYuYwTvBwvxo0Qd07UC9EivVHGJRlI1og5bW0/iyvWYqLitx
Z7CILY4q4krRZ1cXpsnuGh61+MSv0NYIo3yKTG8PVeO62H2xPsL1uoBx0NDij1oH
TbEeGX9pyGM/Nc6V4Qt23+tMQPWkZc6rJ+KvKGhaBnTcHs4vpw9fsQDy1+zKEgev
bhDZPwXcZ1fRjvYb2SWs/DSrXgM/mHpC34llOoYGVfFPox6j0wPLnHUGghVFeNL+
hHr7iMNalIWirAqfBHUP1W80/IDWnfarecnVK3+nTzIsh9GEsLBMQLoDcQym2hNe
b/wompUwrIJV/wb4o8iZznp37mgoJCJOXrL3VTr5bxklG61D1MZX0Jd+UgaNrrBd
18uYQ2LHm3ESKeO08zxt/D3/HfOyUyUkJDzIGqBRB4l3b3VBeU1h/76aUAsxyfxD
9P8k8B5dMQZnMF+uIkOXuDRxsKM9mqw+VuosgdR7623JHV0fZi6Cl9N0/CrGmhqR
fpgz/N5FuyPju1YL4H7yeV5hDfMJ0XUc8JySx4nRLBWldrzqS7HH7x/RWYp7mcsu
jwtDkwtDl/LJhsTHStwkTPrg63XARKMiRvHqxGlBEN3xs2SBSBIWuKP7/mVeCxQR
ZuISUktVF+J741K9aUEHlcIX6ewnNdtVQD836KiyH2EnywrNvqtThyxCZEAjOydz
Fc4orWpzVvRSmVb0kdR8yt+iG/V4kqaYXp1gGvLDbet2BdJEH1AINDYhYWgKgsEv
nsicjPNNXyti8PBfmCLpi8Is8QBN4pPHS9goQcQhb6FQ5KFyn5JzDnsvnaviWs1s
EtVEUe24FTPYIQfkR2SwC1a2JgkBmD/mWhbwRQTKvEuNWlz3ykHOo9ESw6XWoydP
cgeAzQWGHHGAAHuYWDELPCYaItwKtfx2Hm5hJqyekyfXEcBlp4WuYQN1pVfN+qxw
9dIxKlehRk3qWhjrrMryuheKO58bTePa9Xi68Fg6clqbf+I+uGDC514b8z/+YuH0
P0u5Y88AoDU1EZ5BsHf3IByMm+uMhPYbs4feoMAoOd8dnlCudonJirHQ3z1njK1b
1mn0k5ikkvcKp7h3j7KuCVS0kuEPmiajFcp73upLjq7chQgiO/x0CZOHUM33vr3b
erBBEP0F35dveBUSoBB3NTfxjuXC8Jyj1v5vopxu2E/5xRbqZTRKHsfC8/Pq14Ka
nobtpqXcVaOayF2v5ir12pFzM9VC9fRMUYnLWZbDP9WdLiozM+RA3lE/YxawGv6x
cQ5Ivs8AuNGZU0NMt28nicPHNyorZ1eMcX4BeUArDhQGh0Mgruyr1fMMwPIq1Aq+
SXpFBZg/lH2X8kkEvlWgXIF6NOdmdSfDqxUv/d/jLcx48KN82qEZgAuy0nofuDCV
irBgKEClrc4S32+lVefcDdwh7lMTJh7bT1L3UlbamocO+kkXbkR5RpiHgyMVG/Te
AWmT+gkA14zSk8ZThvuT3NtQOubXES2JYLFocjrUrRLzOEhnF2Y7Km6aD/AuSufG
2HLfejM2Jqw9Wbde/LCmqPLNdlWpf7zdBwcCCO37yMTUxUs5gtQWRuu0DQkWFUGA
4LA1wuHrffSOocqGbHWKhu5YJPgywA8nj4Q5kGvAQ7aAsAIb7UjVRa2MXs3vYTfL
Ksv/MjXu66HCU7Akoie9aNCx1BUkYyVnfU2nyh2l5J8PbYS0/F7myQ9FSQJ/4CKl
h56anSKJv88C/vlylj5MDijt3X1o32fZzYqG1DGV8Po99e2goRbGqqrX3sQsXOFP
ImYUi5l4fpOYGnttJ7XGYfeYMf1005k22BHo5CjcKFjSFYyfl+DtClYrcsxg6jac
m90OlY5T69I4hSpnZnaxR3lON/MuoH1vZF7MbNO12OnPOP3iaAbe5uBnN4lfB2LK
ZA51qn7cpVXcSsY07vEceMxlKgns9Gp7MztVZIU/HAQNjInxWrJ8Z6aKcU98C2P2
n82b3mB7ieHn6YrTyfRxtOM1vcCiONAlroG/dTWi9d1bAo4laqiB1Odd3fuQXO6j
GM20XR8VxdeDJvK84SUfaTZEAV6yOnXip+zczfwuZ7fj6CfQicyu678oNwQ5yup0
2LgjpjzdDX+3QjG/+tcgA8rj2AxsClQRUfFPvtkRMdak9IlecKfQG0k0m+8W8OaU
398mw3eQlhhCKGkXLbIuMaOT/kLsOnfBnSEtCn91s0cSz7kqBDcmBATYV5hp/ffe
3EhivHuRO6wWNxNRxcHVw+POX1ICbW9xA8inbS1DbEqfuIIbAWrvh6ZvKiB5B4xv
Qe25ix+FHUF1nrYcYdC0x9PS99zJtzNzoNxJCxTjCCYAhA0AUzueoezor56ifooJ
Wd4NjGJ/0DepjPIYZhRDFDX5uU9kwDXdPeDGk0uIAeXKCITNB9ynIdWSaAGP1x2C
R95rqFjN3CXZ8C4jaqE8dTvTs4opwo6izS4zWWZ4H9nHYXw4CTFcyIdcQAND4kpT
YR+JHPhZDSCKx6G9zO1gaVsDho2+DbVx0xJKnowcA68iXkYI21dEke7Zio9m0F3D
hmE3F5s+hmMoSK/BRsxSZVcOOtaqwwHDH/DWGCOWaFfOJtc5iErBsiz2Zt9dc14D
kbO4hh0dZVhqYU93sKX1Ej1zDrDC1OHkcFpsBLFnBAM8BMButcqQ8XEfZukBvz+R
OdMOr8vkYBKM5MQkPclcQ8/UM9dCaON8GonK2eYKpFDK0FUtBik4302ga/lHI88M
dvmb1RezjJFFqOnXbvM7gZfKSukkNDX3yuiwP4vcEsNcsMo4XlZeRl2cSnSjnTSw
Vs+yhoo9HtN9TX9rCVRznjZnKNsWWBF64ZIHCi8fNQAwjUuytcO6/Krao+fsYMAp
go2FHRegTb7jX3WkKEfgukq3E//lbvgWeYxRZ0vEb5NYVWnvTKPP/i7AjudKvcuh
UqKdy5IxbUZnkW//T+XUKGH+fVCCoKSTIDSv9im9BJFfrv7zDsqtlIMQeHsPCTBc
4/ic/vhM3O4yurJ7sSKCZgFV5ZFYQXHcH9bni5pEbKDDH81vlmA/5R0pxdunbyAy
AP4ZHAvpchEQuc8Qa/ZsIrAdQY22ov3F6PU10hoBX/GrnALkVUCpLePkJwH/mQ72
VsYmI1nYoT2A/ndE2Goo1AlxX5lvasbzF8DFr/QDY6WYjR93hGOyLYGWJwfvpb3o
w1kNSYgF71wJr3T7lrko8fFnhuItk3o+gGZrcfxbCQS+ZuPXBRFXIRmRbHcCPhKI
eKmNs8FmFLOhc0iIXZCk4EjHb9ew7Qn+jQvqgXodnMYg+28Yw6/lDuDruVaWz4Ox
h0rZfrnn9a88LKRFRyaNM7Lb948x+dRZ0w0dGyR9RZBZ64fWQi7d5uldyrsOV0Zl
xP6WusvQYp9xaMWP4tjsH/f0HiX2ZxdE5y9h1Cc0ahA6qX6yDNzEyCoIM+u7rVdq
rCGASOak5VhE6vYtm88lX8+TGEhNUM0AyOU8YIzISt4KwyvEkBX9aaYvkPvqe1cv
hiRH6t/knrPkMGDQlfJ3xbJBopq8ThLentchHERp4D4bTDY4sSu3yvPLQArrZSp3
fJ1Lww388RUyRWDjHYu355wAX1Kwe1b+peW1pBG0iBOkGNykZ4bYxktrAhJFqTPN
ETMdqS5igbZizzYoiCSqJKczTkeZLcnbhgHnS51uOIEof7N/zz4A0NM1oLkDq/Dk
ia+aS+UM+87xtFJf6Y0FomCmZsqVeRHhuiihS5B3NjUoe+wRb84T27grVWM8D5iU
/rH8uYggn4ZK7BppuK+bGIW4EVFHZDRDa38DE91ugzBfMGblPTihK3FKbTKPSLh8
KRpga2Fm6WiM5VkKUMnUNFGyGt3zjtw4tXkv+71OWg1+NiCInLWxU5oASGEn1m6X
YQC9lNx+daU9mpDsS7d8TaGOB+9l5Lvq4QQoNm3K0GAb7TFELznqruez/0YV9p4X
loPrLHqGz5rDRbgOD/GdYmhO4RyVw1GBdUmEHjpVJtFrGEyhgkHqlgdgWDnu0p/U
CgE84mEvRjZhfhB6NEzkbHwfPumA802ZTtWUIM563XZmaW4liWOP5AQx4VjHY7Tv
xP2HYQbN2H2gCGK54ley0RcYSTLy2Q1RiadRg9KAx477Lyo58LQU9MQRWa3TgfJ0
Ii9HEJxtTfVtQ7C1ZDcD/ggs1SxlRcDTMY9x42kbgCnjQRDYErDf67j4GTZPaG4Q
xn6kNsXtlpBsKUbiD7nphENol/tYHwFtytmA1qSjr1Ibz/rQsrwYiKujovM/Ia7B
nfx7J+tcltmEkCDWMy7UsIxQlMQYcBRXeuZscZJhu7Amlnxfz6EfPqTAIgEA4O0P
G1eFPLWxKH+54/aDnXFiYqsTyGnu+FS2Bte9kOz6nF9x0NrT0Yg9geHO5TY0vd5F
YcI5v2MmKi5h9wa9Zg6L3c6l/JQEVToTNQ5X9+8dTdShgczAj9qEok3nZgi8Kgu2
dwf4gpa0BpIjQefy6dgdcka4cICY6C8DFF3S8W/AOXULpZhGzbMpEgpO+6ShAC0m
7bjC/Js41PHyz1h7lzr6b69CvVTVw0gXUTi/KmT0fWU69CHCSTmxj7tpK8E25jv3
T9VKY8YMCEVFN5Q0EcEwIu6zM/CDOAsbDUaN1axX7Gr+SX6FPRwmyk9+LeNPptZn
lVh12KHkdCuhprdc+rU3hTjW2cEdYW+P6FqPP0hPQxPEqzbOLy89QFlfcXKqXTFI
+pW5KmycbuNblfKeZPo2Omw918l0JM58M4l38GUda3ogs0tdjio3hMyiJaIsBznk
i5+spvvaP5M4KHvDE5WywWxBZ3+gFdpzvtb/JPSJU3pMeXv7faVepZc7jAuQ1pqc
BZpm4Lx4EOE1vEasNHVCq8RNv2/1vbQFDENJ9wCjo2olsnFBQ/8apRVjzxFrYXT+
2Qme6MnydWW4q2d46C1wS+2T+N3H52Tx9gJ1eGrQEGsCvYQP8t+VNt40kc+3D4Er
IO+AuAIoShHY8ZH2wCa8HrZPrT/Z2ffhYjM8Xp+vwP/WWcZVd3biaDFwuIwMkNnv
kXssfgWRrs4/cYkxzLNV6jPRXs6saDsiF3riyxFwspIySw8GfkaNodS7IzDv0ocE
BaUD/BGHmHhtSWkxwiDVosqF7vw14kArGpluZwHiSvpMie+5Q2wgY9E7OA1uEL7z
rhdeIa6FKwugTGgjkBn91OMCghaTWaoSBE7YGO1ax61izZAo2RQ8ixMgJx1L1wpK
dGRYp0WguTMe4QgnrRCOG8SaBCE0FVGCcoo11w8zJ1U3YXgzOxUb8hVnIGHA2wYI
a2VWU36FaRTZkposGxNFoVOcq76OQN1wJdQGB5MKRKgnxnD5ByNQmarUu8JdMa0O
D6EYuW/0QHbbjYhFZrxNB/ra9+yzoktPsRMkwo6d0oQOs2SCvipZHDYRgmoDjYD2
94xXzrAjoNYptF/NX5F4V7Oa9CFT6+FEW57PJh115nC1wqI3CTYGqfPkbzRUI4Bt
9W9CyDSbEECZ/nEoZKk3mtYuxGgvNb0UY3V8vPDjcJ8ttfcOzy7QWvzeotBwO59V
ylm7vZ7Gj1TFspc5bQg8B8AObDZRWEGmp54saXlnX5vahA+1WhCTlAFGkp+JOgKS
9cHWgcayoxz0e9SBCtqAATxB7v3BY4E49jQLFJspQfl0buRfj7SAeXO4uJlz/xlC
bClsFB+7mcDfSteQwwknNwxApzKw9qS2m2qlS/4Y3kKvsnund67O4Z5HeWnL8A+V
2cTcePrRtPMDxWmxcwoqlX9RDvFy7QqZVvQJ1EvQLq0aHuls63PvZyYp7rm06UZ5
RE5a8o5sEuCnKnw6bHll9AaFpqwsCt95UHP2cJHo6sAjzoLmxit3ryvsf+xiK9DU
/T5V8RBtdslioN87Brk+Dug3LxOT3BF2NgC/bt6p92TOgwMUUApi5jkeUizXsLWE
LSBsuvLVWkTNrESItGdFUo/WEjou1FA69XHSzfZSAT/b6IdE/aJ4OgCmpTUEIPyn
TRq/3uqUtNG5cFT3bENp1XfxdRLur7jGR67dex16QW3RAkKIsPJL9k6jfCwNeTbR
ZPU+U6BuX9e8zcqP5fcCjHCljIXpw/ceAGT0ZqfsZC70eISysWQSwnHyKF26M3UI
9rELcfPxElp94K61ypNRas9t0KrDHI/2++gGPQKP03OoQ1Psqna9W2mUR9AMu3Cv
/0AWBG6aqiio3qQ6oWXnO3G5IoSqEWRPxoa7Ptzn1JiznbLV2Zncd9JavsEAapcC
K8ZSDF+TG6Suf1mZbJkbBpMiY2on38zdeG7HC+yzDu6FWkTBAeoSboqkHQDtWLHU
yoCqH+c1fUHAjzlqbtqMG2WdPGCT73i/q6V2WfD1ghZocQnrn52wde427u3Qxkp3
nL6xo8g9pZXIjWz2LKs6fdn7nusVCnwQo80e9ZRsOTgqnqs/Cs3WVdGCs5z13a8/
tkpQdQ+ckmWGu+rqk0h6j+RLAznS/kLYJCcgvp+YxBtZ9I4BT8ZojOZXF9R2MBvX
Ru3IueocqQ1Vrl/nawKedetHz2aZhOU9JqQNUjH2tVFreF5NmXW10LX5T4SD/AUm
vvKU5hVRdkHfgZiEdom6Qw7cXBbc0oRCSD0nYGPllpcTXw0t9tp8uZ6CFvCplKlx
3cL/tcZMeMe04dPlwgB7WqphV5+jeIN+Rz1aaLYj8Wu+XPaZt5B2osqylr+HyFLG
unkFBMYiygHcowbwLIJF7p6YI1n+PA4t5fyHfkJ+0PqFYQDuyHYCN+vroIJaIAHD
jisTunx8QghBiPOrW7oB8kTrxRWWXy1Nq+je0bCzm74z6rLzu5+7qouAIf3go46q
eOr1jjX4Wj1L1f6cj/6g8SJ/2Iz83KUJ8Ru7XEsCW7B7DQZ2rFt0Ucsxd5fym62/
iygCGrH54wRO8IVor/6M5XkG+K7OOid+o1nKgd4hiORKEPETioJnkoQyQ+t4no/0
KUF/iqBUbLIUWjAL5KTCm+aJs/qKhiAUswD9VoA1jaaeuOkPi4HpLj/18EZBgumL
VFpDI+YTzzzeLjf2tNcAuUwU15EaXgCWgnnNuptSRrr7pDIzBQu9Q+X/KTrUolT9
LRpRgnYRPDiMlijf1eUpbOO3csGK7ls/x6uoNm9KbLUgSO7jv3iYfLBImcbojNYm
X03o4wU2X0XzxuTy1WNWY7EbYK1weqsjWFTkZ+z+SNIA7xiKOnuirT8UcocRgQJf
CKLz4uPoWJiL3JhTiOYo2uuiQJmOdW7rBBwzmzd2bCqFhXUOBcEzubCkoApvURWc
OYaY6YPzHYTnOr8Wgscu10Fnr55uZbNAcjc490/jhfSVIi0KZlfLka72QSWPrVga
I5Qx1hFziC5NigK9vHB0NnEB9CP4c4+kmIiIXs4qVtzhjk1vN8aBjjWmAaXIGajU
os6guac7lY+ZK6UBdfkVvfs6esTsqpuXkMfsOiD7/8b80mKgnFAIgVpFqOHLP9G2
BJPoc6Y4bD2MMcdCc1DbepQE/GyFM2JORKxL+f2UV2CMP+NgTs/ntMSNPgyIZXId
b+yPpWTQdqnhXF4R9rSxASqx9/w47B9DIg7vm4/4MRh1zQcwdMVQWPknpyd/QW4U
pYcrOzZn8B02dX7LooGq9E/rtTIBfpdUrq4QMT7Swz60LLuZeBrBw93gk7Yj+9VK
kHZ9XLTHSXCfBJew5w1Dy90FzFSv+Nm0o1unf+dqMaQqhkTr2klvq4ZrQciqLX8N
vwp1SwDpqI5wBY8Q9tmgADLkfKw6bf6IP11FCmyPzDDaZ4tNKCDM4l/wy/sGXSpH
GPJ5l8/kyXqUJsIGhfLw6pLVe/ubuqF6q2rV4SZR7C9o1GmjVLNUT/qFpJItwRT+
sifIb3VsBqbJyoqJciVXfBkUCR+YnrnqA6YYjTJyG5msaBIf8HKY8mBXfL075c1+
vjtP99GPwTcG23qqBsU7aktgh4Ab9IVrPmgazBAbRpf+JYiXqy1jxEADOCImH1dE
IjVvpxIaySsOKE1Az6s/u2hHtz0HvlU2zk6FRN110/44Fy3pL5Z+tp05e5hDcTix
H1EoPtoKbCFduZgni0wkEzWYC3f/xgJNkDUFeRbpLNMveDpfOje5ao3qu7Kc6TaD
sPb4+26t+PS1BeY9c2pTvH2kXUhzx9u/a1DGXcOHMiYdetWRTXCa6DyKWaIZ0stn
3UMQ8EdjrHOK5OM0rrr0kNP7O017ysb9XAajIEG/Z7qc+dvbC+dVqM3GHPAXaN5A
GNU9X+UMFQw1egvkEARpB0JoITnJd6TWDyS/M/hltfIIGpd6nNRbtxNxYQY8MOo5
uqffOEsC+NbZihRT7PefgR7x8dn1XDvOSj/VMnpd+jcYEXD/i50T5bVa66Wts6Cj
0+cK3Otvv0+8gadYjLaaAZVdA+VJt292KTmZo9cMQu1URERrojaaAk2smo6ZGHcu
Qvmpu7q/XddcCprb7mE0vq23lilkOJWMyoyJoCjxmbfo09xmrHh0Hbq3ICiYpK5A
e0LoJAvp77nR9us3WqiOk6ZyT50Ldw8+8SEW05X4bjElr2/qHX/unSmJTHoSaqpo
L/J9ljUIl24DpY16hIOEWzGnu+GZc2R+PprnVCSbOMs7ZIW2Bkyb7RHVWB43hKk1
fQqMgaev/jm0VazUusxJ9GsNwBT2c6KscY8IzYPAEmIHY5CI7CxKqoKDCKJF1TkU
2EbNgw9oPvMFILJfrmLxlX95Xr8K8VhSnvxKzZ7UzNhFFMgs+URefk+wdNDNSCHT
zNKrKZ/pTPNw2YxQRyGSkKqacXhfjEUB0fjA7N+kT4FvzyMxgg+EwDVK9xwaY7GO
Shp3VBA9zMfzip33GePDfjUlMlfNY0LiptpycTIug/aZymqQ6GI0erJAeHbojNQF
M5SoDINa4bGc/KlqciFEVBSMwTAmoiWQ7zpy2JQrYuf6dkRozqLCOvi8HX5ocpTw
uwISyiHd3gAhlEZQnYWpXsn5rUZC2zZtuDTn0z4lC5O9EwELPmB6gDPXASA2Df8v
3TlpVzERJ3HcQbwtSILKP8LZSdso4TRRcKlxQBhL3nJpGIrkFzOwVnO4yUEuB5GV
NSiQ02Icjx3XVvU39dKHhOvE9cZGQV5P2bsD33o15v3yXwrYTuudMdCswU4b5nej
7A8o49RzWtvL305QuS5Bl9nm0BmPFSlZx948vRtmyGu94QJcTDvZGErN+FMy2JuU
f5KLQMgdz4Sa42ZneUNhyEVvaIeKXete1cBqj3b/8xbLzLU0Onptu1jyExl8AFZ0
barqVidjqe4dDSnn8PpqvAx04DEv0xuG5fL+bXMdSQxzAwxoLoB1/MBBvHF5s151
tp3puHQ60aD03re3t0tF3cSBin4q1rh3T9OvC+1oqwQBQfnLuS4SwMFM+g/LSr9z
ym9zb40lQD/mZMhsr6sV1f1CiwQPDlbQ4OpR5DDhRDj2dZdRFUXX/1G6VwWl3qub
AiPvxZ4HraaSc5YS1eCeOlXMUNxsiLtMQbphIuAc9Ytk3vAf34zbaSqKkHLM74cK
pW6vhSwtqA4t9mq+oxSNqSi9mic0pnHPIy2EL0hY2aGi7YtA+h5HnI5ReV4+Su95
c2K2e96VIFmlbQUfzdAG5b+YOlNRKCu4WNqbFcJt/d5El9XfTQEd3LiqzeipqCUf
CNJygp065goLC+jO8boBcmLVr8TpY6bAvxOVELBJfbjVBbdCe/u+VkcxwJoiPjEb
Z4SOxXlI2IWTECT3/j/wZ8LeJVpstkC6YjPOrYcRX14VNfwXjOvxG3iPSWDJ7q1G
vio0umyCDO2MQyGq2xGegbiqoOW7tu/ZAs1VcL50pHLUVa9EMpI0ZYZ5w7RP7cOH
243+LnHHDfYMSvcmht5y4fxabC8vrkdL5iaqRfWvRNBS+eymzj4TYMEgQFoAYR/b
NaQTIsPld4eQScVJWsSUg+xkXWF4sQdt5AxKszTpebY=
`protect END_PROTECTED
