`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a9pW3QYCfxjvvTHNcW/Vc0HL8sEkUHDIoBfNb3B6G7NrXenmfHI12NNkoUdfo9Li
OE0mxGOribQ904CTaqboFt60qUrYr426MRvHdC1qur+rtHMTZ/2ybk8OufNMv3UX
GDQKQwZNfqJdbKrKqjAh5TjiPFR+bcbphbbKqftGiaMfGiGMklIvfoEnyPk8y0/s
0r3GGYlbY6VAWRzgmoM1YhgXpwy1h3cj74RCxG/nho8HuCerKiYn1TBm+78bNuct
t3KiOkCL5YZS9M60CuTXLkO+vvoQdqnyijSN3j4/v7mZKizUiTF6ABYUrTJTeVnD
QwL4AYxMvOPF6oBzKHT8dTwyzMdxNyjUqBEueYjzrdFH/9WF8IIeHW5FhbrrX/F5
FhJe1ysJdRQXCdtMJ0bIF8/0v2soEiO6gKkip5LCTmiHL3zWPtmTvKr8sySppMxO
C1TDe4IHozPIYfM1+N2taI390RapLezkWPbzM+7xpzAQPpNhMuS64XL7QloyO9dn
Nz9gHx34NJU+b+jxrNxvqsENGj7zPBNVQ7NMcy35oyUTNi/mtHUdjtU1G5bwZiUq
qWIU4xbYJxVq9FzyeTDv2ks/iGhOi3EVcAYIbxpBBRcG/L9oxlGHPqoFRVxUXhrg
u1agJMvD9hBHKMVeG9dyksx8TekIEO5q/UQhVaBGa12RrNhgTTJrZxNH8zHpMtB6
5JXHkfO9W5AP/qh2yYc0TMmKz7GBQNLWjtQu7zncrKQM8lrtTs7RUWkSBHxvfyOG
v7orO5aP3UiJg7BGnq4fdQKx3vS16MGT2kBDQ7YfN9FCGa5lZ85POALYAKQstMVx
AChnzzxLMXTdzhu3nQrcoru1BqgqiWoa950KSGyByrJ8IjAX+/XJdXijkdmk1A/k
44OSxsxs6jF9ziG5PwgpO4/E52SzNkMHymmXvzZr4OoMKcldbM9nFxrEBlDoDYqp
yCzrC7NVisANgeWTvJj7TdKhdDEY5CZDs0OFC3nDCrD2V0yae5zGswo8WORtOkI8
yeNKWTdHEdO4M8nDqdY4U0mbM1m5AuBcJFq72vUqHNUZuy2SGp41EvbQWyY7OKKO
k3urUYx8KkH5hrqV7SpclPbxtH1IABPB1TPKmNL9bA2xGEbx42GVhz/zzjnUN7VH
4wXqHz5TbuVIJcKfjfe8oYivazdeuFlWDq2v0Nmy3l6zOYBwT3h34l75f20xWUNm
2BwJ55Cn5Jtm+J23CBrzHPwT4BS/sSzfaFpSxN0wCOu1vLX3J5/J9NFU9deiilRV
K7GD4KReAIS3MUjT4THVrjdI3Vv8mIVm+5PSIihV1neJLTKkiW5L6ZbarZObdXos
52/6RfGhq1+MrxNbY2Uol89VtzCh7WU1y0h/+6UNJhybMBZdNhgNVOGapg9YAOQ7
7vGWg/KB0GwO5pj0pAlaRygeDN8xCw166lXQOA9vmmuDBvrgap8/L5RdxDATcZDy
nE2C9A7nqUe4FEcS2L5UC65ginGWa8KZNwaQuqesnooQlw6hvRWWgf/DLt+nBXt/
MP6jiVCT8TT4W5pglTefIBwIDoKwKREJAZ8jVbeidLfLAFNnsE4MUDQRywqroeWj
Aevlk6t6Yq/gDuRqv3CiG0PFrfjhkPnjf9KA6O9t8+xiG7XQtCXJiV5l/qmGc0TO
8nPLSfFmcOF63cT4IJo/MEE1BkNENvY7Y5YieQwnehuUNb7efrQNjHRYHe/8pOh+
k1MD0yWBubA6CtFIHOmPbG+B482V0zWASJoWgnfc8Ts+CsdiQNvVq3ljtC+n8mxp
lDUSwNCqP+L9SUKj72VayyDx7MN57cf29szNKlgkdiOVqYg5xmDGrvNmqQXwFZ8G
Nf1xbBoDGuq+hHvZUe030eD/xJEVgkTsUy4PrsYbYiCadYOfsUKIrHIadVpzXx+G
LjlErosKl0T3BltUEukByPMfNT4WZ8+/rQRwg0KfpMCH1lReWtu25YlnjIh0xxOL
dLGoI6IQH2O9ul9Mk3wFHgIjc9sYTyprD56n9Rzfzy/8oxi6nVzhSCRM18dr3hV9
zGzgPbcK9BrthDdCKzMMel/hjQSCGiLWoLb/qL2cifKCkdO8cBKU1pGXYAphZHwM
4yi4X57whLS52gU0ogRQocqwEwraipzWmcYnlrkdyf2XdD7QGhLxi4lJHoAueuBy
B8RVqmjtHJMfWHHFn93R/1wdMM6qDk8jebva7xupzgb7RvDLYMKGW9xv0r354U88
jj30fq5wz8PTMBNW2zdJ2lDmwxZ3691CQdiZOqD+VirpEWUxoxFjIN6jfh7Qf+CE
AupEJj26OFW4W52PKfvAbALN6v/ksjAu1dMRkcbALp94YKKnUDIxiKajpVNsCIiz
urRqRxgacO1wxQwQBdkQJmvz+lZMy8Vlelk9MipiDAgtADV8T5GXgwBlXEctGksO
Gnm/oKqDy65umR56DvFhgoxKKpCDqfm0xuUpNdq+y8S7Wbr+VxdR+5vrQlAovVT9
M5Ekqb0HrJEGzCoT4iCXh27UcxDu0shHce/XGDuOL5sUD3nmcmXhYpfpVhgURm8e
KuQfOgt6zN55M7Bou1rxH1H88FSyKQ0+CVXpeZvVNH5B1s/6sUY4IH4PkcHx62id
/bBpb+BpScYfWZ3GyIlkuoFI11IPMX+LuV2v5wE33ZIdEgl7fd8/2EMCyqBaIEOV
9WsGEYEq8Wei+w+ANxDjiyItKW58esThEM3/XO3GqpL24/7nLwzZMnu3pSHIDa+r
+JIw0GFaJAmWbu1CkqrHosLCkNPIXsgnmuZztmQ83bXG681LU+m3mlzgttYcktAf
TxBQ5uv0JEbsSbhvVQjcXx7J4O7OzWaYaNnxGgJmi7uBL7ZZsAH5K7Y1gzSwU38e
89JZW77F3/LjZXK4Yl0y5brQ0mUWfhBSRWYy6X+P8PQ=
`protect END_PROTECTED
