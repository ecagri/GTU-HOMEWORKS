`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rhhsfyBuOOssdQa1QntGNlJn8bOPfKjL+o3k/5bR8NeVKTvdRzhSNYnEQo4nayXk
DTQUeSM6SeohszPTfapGNMIKDHB/pYtlnF+TlKNkFpx5BrDVwaNj7wzIioGEaX9L
fFsfecbgxsx55/5U03xKqNWNvujHQAzmGWX4P5tmOucgVuCHrUtPF4Uj24SDAhqS
avW+Q4SG8QQ6gmVcnH4GT8HidUzVMVhjoAHZKS7ApT13YpmoFPn1AH2YBc1LRFgn
Odw4irZ4y5Arq8P21RR6C3wBp1UwcbczlaYLOwFwztuNFWLrWKCXZhCd1iDZ7IVm
PmI8sQ0YW5lrOvavKWqd+wXIRGyTJtar0YXEQIwfKEIcr8xAlIQREk+djksDU+EJ
zpij6FbobUC79U6G8BoaOSRh609A3CLnWbtBlExCA37Du+Fq7paA5SafOS429QhN
CBEum0Cna3DvGPeL90uoGxpTBKdEQ8IggFZjd4zqj5BBH1QVWPxtwGE6EXyiSJNP
jAJHQO0Hc+NK9jr6iKDFCU4D5MyozX89AtTPUMlgnNg3KNU7VUtDffuvVcMBTrk6
AoWN0uNICNdDcWM0a0hAdwlV3kbwpTGwQH6sU3hca2+RT3Txyd5Vb1Nuikuo4U3J
ldHfokkLgKfCF3Yd5301VsF02F7hpuPAynax+0SlJa1mEz6RzKVtyGuHIwuQ0eoU
qokWBPRzTv7RFh2/vn7V3A9v8AfSVGFIg7OnCs8IoP6Rqg9A7fCl9yR3v0SEsArW
+k7yNcPKp2Hb+jliC0VIRA==
`protect END_PROTECTED
