`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h/RB3x7d89H9U4Q08qFDeHekM3DvVlWdmULwq+esz3029cetIfb/2u+mdDpgrAux
iOG9X+QuqcFMX5dwa8TcfzR7S62Wxo3xYby4OyYR2V0hTdx/O3VU8kmDwbOU7c34
tPWoHVIbKp6ZAdigQkqU+z3Z6hOL053szHCigSRmMVCGsxy6i5g0fwg64x1LBTyI
ce8O5lLe76y3N3pW+gMBZ8qrh1npPeUchWaox+VmwgFMtFTBe5GqNhS+ssy5aiNU
qmMSUVA6DcP5EgZVFuOZpYj0nC8Pm5hq3v46b++9VRkdZc+7diOTMrVNHda1vrPm
lBa5QNfsfwbbDZ+KEYgvIGpHjINoZe3aiifoSrNXA4ZxudqhPacnHGi+pTryAN+7
`protect END_PROTECTED
