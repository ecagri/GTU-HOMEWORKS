`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4c2rxFwKP+lte7U9wDKPR0teRdw2QBgmR7tUpCy2yZ7dH5ziuU7t7e664gX8XHAe
RU0Wt84BpiM/yFA8XE+aBUHQJnof16UMxSbkxXlkXbQhdovxdNwvdcC5vdv4KIuR
H+am12ELoSMhbGbPkbXDBGUxDlUEIXKG12ikCpyk93ItSqfURpadxC2HdlFr03bh
1onvhmXmCSj4d4IeS7qdSgvUnoBNwY9dJ0EaM3nbqKMRMGLmPGD7ZM/byLbrCUMs
og1PmS6i36Q3F/XgSW9sDlFu+vaJx8fgBMR5xbO83V5rcJcoYSrSDJ5WSDLy4V63
XfNj+ou8wxLhCsWSf0JOFoV7uCwYqeLDNYd6GHpIzjbBc3617AXa/7PD1KZDUdMf
XH6I5RfYi2B1kpIyJA4Q7A51nRwPPDeV68wKcoKOlnE=
`protect END_PROTECTED
