`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dZXWjDEG0itdJcyyiKH5RXfFjfTrK5ZeAZJn0urNmxJDnCtFMaB3IGsr8y9U4wm+
02sz+TW5K89y9WAJFprckXfGXK8vPqOel2gRbE+oN5kR1sHxBVHC1sTBcZW77jbh
D9wgspoxoeeswgyIY+MThDVGWUeJBKhRt09WzcuakpwrX88bT9YGgoWMPtzYFGxZ
1J+9plypGzUJZNquJ4C+MD/6t70hQ0FAzMn7L3l6IvH6ePLKXeGhESDxG5rSViBd
CDAd8QmaNF6HaMsOhNff8xf+tvO4644VT+TeuPYBrvjJY3y0zV48sAf+6JFWOPp+
8yiBWDNCe6oXLbIfA9rEfBK9q5o69cy8Qe5TuMqXXq+VV6IDuef5//B0OGf+ys9m
xEjwqhhYTF0rMetDet7e3qXkQLqfgwePMCw4pOTL26Yh00b9hKkAeKzB1fA7uzeV
TV25vQZcj7DK+tICNaBIUZc0W0s7IaafUpneP97cbnb8VJSpC9z/ZIF8mKd3nIJQ
KPP2JK/9HIXV53lF8X1mqm4cfg7pgmS2Dog+amlH9gVplenNVxuaQtNP/eR1uy6P
UXg3c6JAEp49dPuM9Qblvv0UlZHHtVFflsIiZySUeHVIo77yybo1qKWn50Rfn0pl
LTzsCgNxMx5DvU0lQz2AL33WqocV7zpyboMHmj44kTtREZj9I/f4muKgZvN/HBK8
UV2gVohkLpeE/hzkukmqAcis/JEG5cbQKbnpR/c2melkU2SL5zNG1gM9jQsHtJkV
D3I3yQPcuIulAjvm/bptQyeBosMqrLCzw2zlplKpQRo=
`protect END_PROTECTED
