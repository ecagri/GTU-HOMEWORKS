`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lZUMzwvwviS71PRtZ0rXntjT0N6+scH+HQbZu/h8YO08lOZePPVfWfsB6ZEusgrD
EkfN7Q7Bsx8FiSa20FEt6XtWvkAnBuKNJyupXt9AxW24QYrx8sx2AAdhL8fXENj9
54BswliEm376gFRJyC2v86KWJA+0jHWX8w8hSDYYjjC2TzAHkL9sN8cuDQ7FBrHf
IuTGBAcluH+0/QuMv3uh0crjk7Jb9ijF252OpHamskTKcl0DDhAVCnus06A8bxl+
YtV3h1CNQP5NT+O0UmxkzMlZi3fy7BQYF+DAq8qxyudmVpkosnuVskF9vm7vyqQS
stHxkLtGXyfSs9nAITYZxkEZ3OcTpiUYjrzckZPl+EFIkHRj2WT26ccs+jbPxRUD
T3nuo891V4ld6Mt4Soqr7sZwPPXnJiMjBI0sXmRvKhOR03b/LsCG4k4oesq1JqDS
tPw5YfsDLSUv+Epe2yZ4NOL2dpFAjZuSyn6odmpcYPGmYPjnZiFS7g+13yPJWw4a
EppLhAAsGG5F+du4iU5Qjx0vm7GrMlD1+qZpqTKcyqW3kGmgk8MNInnWgwSbE6rf
hN3vxWUJBxOFNoaKrDa1Np1/BGbUvu1K9C/VI/hum7kLmd7kELCjAzmE1xPFVhNS
QU404PnOJtEb7CD2/94rdoULx9QFLzk2TBREMzFejs7PcRlot215/zjaqtTFb501
TnInOdRzHJHNiEJIPWb5amGy0k0mcjDH67KeSExpH7hVVdhi+E3Za8BdHwTwF0T1
NKdvCuCAkai6Qkw6fnJ/jXtcH9/YlI+aTTAOrMR2CQPan1gLUaTWTzkWdHzYVrbD
82ROGAmpGmwPpbZHEd68VFb6rqbVPjlyVkcGGpazNVtIAnx5rnr5jDsfLAF/3f6e
G/jb4nqcH5EgSzsEKpX3ccPd4yxZu/ovCPLGBIfJW2EtY5Eo9HUPjy9DIXInQi2n
zUTJLfFVxVGRmWw901g2ikSUIvB+htE7Pq/1fRVyI4zJTpoWB/HcWq8hCxWagoWY
ftaTt7S5d4X5oynBSZnyjNeUt8Kld54PmnONc9uzKekrHW9blltubSZH7AlZ1zbG
73YzlyarIeDQu/4y+MYR5per9YgN+UTM+lQdfaXNumqx9yZ3NXxjejdrn/rUWY5p
IzCpGnyV4LPoNnOiLSQpHWalztDEBVkSno5hGPYFCcwMjD6WJWlGcR/PF5IB8TMQ
44ZbZ02B85FsYJzcU8+16BYtAFJnKAh/XFNtBDUvsOqQgSLJFObAfrTFYa0BOpmv
0GOtULrRoGY7KdStEtF5h7gTuPvdZYTuSdU3Jw3ShMpB6uIHwkzzlqXolkKagPJp
7QCpNNkc7fcuQigKig9rcn4oexIhuo0YokGJcDRaLZFqLYWCbKmZEPBW5YQgByZU
wmC3HUcSBPOus3AJZ/iv0YQ5W9S7qXCmdCrwWoQj5jQBzRmnbtH4hBEXUYfO8JJG
`protect END_PROTECTED
