`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NoXr/FPax8ygq+01t24Z8AtpFS9o6o0PfKwS+QuPKImCegz3pRFmQMc7AfhTvk6K
h8Gzesb5w/w60GcGE5vXst1080Iyo2UONtSkifoCEgf1tbgO/IgxK9o5BDpILFp6
/s5NQ+UWjTMpfmey36dBq3O2SCrN4LnivEIjsmfHWocecyaMVJt2ywzOxSHPbm5c
GXglGw6IJew2yDEHRa/kXMnFdm7wQPpES/WxC2OgNF9V928NVnCFEd+R2uuiNrnT
CfelALwfwQh898nBQSusSXpOwk1iN6SfhgDzaz5tFS0Rcj3CRZ83fT2mAEIPi/Mw
egDCvnadOCCzATrdMZ2OVsexx3/oMrW/gBmxPjw5BOncq1z0aD1V+ZI4n9AsnpQn
pBeeWGpMOI8rN/qf6MZ2LZUeca6HxDa73WnnoeKJkpvkvjjF7Ny12cwuqwk3yLRD
JBFOk7FlsO61bTTDNavLwwtJrhOXZgQUWkR7d2q49V3INyVm73A+JoC1a1O+XM10
HfjUnRtoo7miSQdc0XSTCqypH6BuzSYgvOnxs6tjJc1dgt+dhvDnUEZf7ZwIM3PL
nxpkGLTZSZv8Fb5s3jquDytvWLB7lgB4hcZr6TbJj02hE6JnjLgRvTHLPeeno8xw
XmZXpjLcBWpTy6hOyOYcYxxsiFUXH8SolDB6vKdb0dzkFmxKNmdMPSKiKn0GuwzR
B15bcPTgkcPbf5et/43bBdW0wtd3oIVRRc4zPZcfpi1EBaaP4LiAyHUwjKlMXbUK
Z5O0nqFUxyZcObVRw8T854sBzyAEE4q8rAnXrYiMHtFm8QNC/C0I9VISOmGxERf6
1FpUMhLXWPhsYU3mCTHsg2MVK2OM4qAvQ+pYaY2s9JnQ9wHhQJaYcz7S+WlIe49w
t8rRFBCSKq5sI8YOz4hzGq8ggRUoNeHE3jt1UlYmodOBAIJjFxP4lYrpr4+ibmHm
lBAwO8WuBJRZqtb8mITGbCg75ROmCxHCHOtnKvEvxZR88UqIjW3zf7f1d7amdSnC
q4CcBQ4qIEGFMpZtxNQDTmpktg9DN74uUBzIr3tw8O6n6HbUVvAYwDBOcD+t6B4X
w5ANSYDVxmSPyK6Go2Gf7IkAZWcrDjHuuAgrr1yEGkjGlGbKPxN55++OchEpkecN
EmvJ4Ay5+9lYE4sRrRWntUdb86zmthG8wFSh1JR/ohFK2p5FOYPMryd0VvMWk9cw
GoZOBOSmkei4637u3YhzkQ3ZAB31vKvItkSVpj2FlAGE/XGUZf/Kdoy78eU5NS03
y53vBNLM7Icx1+ls6Yfk4v3O4g3FWobbUORWrL6oEPxrNXEu7ii2S3F/kKPRvcdb
JIBgs/bNsZn24XjU/HP0sw==
`protect END_PROTECTED
