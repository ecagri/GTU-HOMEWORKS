`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6eSoX4pri+MFAzVoTcZMtM0ofXtROOa6IOyzJEIPbTv1e9vVSOn+pNU17LUHO61C
nQtfEseCfs5KWBiBHyzgQ83dIc2fg9eVb/TCDRZOITI4QwUlFCYryi8mqFiaPots
EpVusBOfOdui+u8p82CQxDArLqP0wq/CBxNGmxpoozI/Qss7D8kNMK1MaXImdb7X
3v2zp6YCHO/EAjGk7IyWm7XSrlmbiIcVSdVIK4Syk058u8XnWWEVONyyXZt4uQrq
7Jp7nd+ueEyTOfCXa2bm2ASqvqQFBE4eNzklm8+Zu4B9XVMpUvndx3eKZaWR0HuE
GDV62vq7on22BQWJJpWE0hvZyXOHJfArdiJDDg4S0XUMkn5/NOfr1ct213AzA8gV
9UvbXtqdL3gO1fPK6P2BXSFXBdNNIhBjBjvtQ40rF/nIt9r7zvuBTV+2ScB5Y85P
VcruUHng33FQtmG/n903O8PNQPA5gBp6/EhK/HVD5PcuPbKWI/djDYSm6RpBGJBO
k0sBXIABcfeiAyVTZ0WqK/sOVcZiZnvH2vGhiymJ/zvjAISKH7c/jkCcUgLTrBwD
nZEZ6tgCJddIX7wM7octduYgIV1fSJXCStHKw/5xN6z609fig64AVjlMOXVa+mLF
LSg6fvdw8iN46hnS4FXCMRw2JpzE+s3i/qAHBwz1XS2EnSWQvQYY977TtNzn5d/l
TDZmNwdISSkP51QlasANswqn8gb00ObZBp1UPP4br9Q+Q9ink0PIVfa8BNPq9CPU
EK/jMJpz0tsEImFuWNC31sgRyEfWXZ3qHxc8ASxdLI+wDhxZy/s+WwoO2+HCY7ve
KVIkR6WpODzXglnyDX0gZXLbGpxip4kIFn3WJj+SXV1CHyPwSUIytuAyV2y/uKAy
eHDi9q7ZCv/LngZZWzz/IXyuXmIwqm7srvxKqdl+NMyg8Sj7BqRHHxAHUqfhn6vz
hkbPUJ1LmZ0e/TPhqxGy5v3x80OmqkQUtQ5UEHJqVG5pTyenHFBi+krGEiVSoiPU
0LKeyV15qDBP7UXy9DJhxjjR2PMpHV5zAdpz8BzNUdJejyr5FAMaJsJjEqL4BGk/
vUCJq4kISrTUij+FNTKlmhw1ExPu0w15HSiIui+mIddyDE7yBhvsRCw9o7tLWvaS
wgsTh2r1i6hNN/mtxwxv43hfZvYWmoCkM5hb52/J9X4fLhliQa7oNz2pqwjjHikm
EUkp7ZU+Y4cTPcYPM2PdIKXXGBOjpcnpDUeQWHLfX3gINq0ZqqRPXPO1VuXINmC4
n24s82ZtCEWKqWSsKauDS8Wj30IO6fLaxZX5ad35x/j7MD8bUBhKU+Qd1NXknD+Y
EBp+5DB+dca1qaaZyS5yqO+OiKMq3wtdx9kaBjHCG903u9t0weeo0rsSOzQB7RiD
mhIyRxH+5hDuDd+KqEMl5wlGvYQtKMqXW2iC27IT08MzH3479dh3eaPzXOeuwg66
cqBMEStI5NcIqntqh5SSlhv8YJ8g+/PnIVr4rfKdTnJW8qW82ECuQmg98WS//+t3
I74flS9u/RPuOpBZBnlTMqm3MZSV5qINq/8l0lxNUBpQIXm8xrEjWpQSUgMQQosS
Iea30FtGKAltHPO5AxYiNMqmVOJRPc9Iyq/aQb7k2WMhK2EkpeDWy9oIQ6SXqgI+
Ecpb5oi90jjEkSAJsJsu7PoGuHDMhvbp4b9DZH+e9CqdNpk+xTMeyt6kEJxLoDTZ
ap6qpSFOCrf7zUGMwANB+9SJ7tnwGStH16ObaYCuFktlJ2rmCy3OVXJC+SkO4LcC
9UkmJ1VasapXaGpas9QFyU3BU4FXGJiMGeeRhhIa2/9T0M0TSF1dn2n0MvoDaiks
usvMNzZTY8VEssg8/r+azju4295HKlSjLHExh17teM7J0j1tD4RtOwv4briB8ZKb
BEmaqUK/9Exh3Kh2OrFMej1Q8utkelyWCI9xdLSNnBH1fWcFu0Eq7PyLRaVJefNM
ov9qgglGn1iS30UIKoOyezdadWilNYCQ3BSnDkonKULsJJdDH2t+6LFivq7KbeVH
ufo1AyWbW1iTcBT2o+/I3YQdmckXdh5mWNmYnjXQb4G6cDOwSzrp5/xQ/V1yEOUe
DGSkWsu//qTZ+xmrYlwngPUxd6kbCMb8xNjj+IhqlooXMDq5Uzi3JLxjLcVioBKb
OiD1K/se8+ZnDGPsusEUGQKUYTcF3W14Vcph6lR9uKoGrR/Jn1f9XarZBwqSJ8M1
pE7m76O4Sx5tNlSN/IjW48Tdf9zpjZ9lDjOyAO0ZCm0pTqT9m/XAV/MUH1fO4Fnq
V92Xz02VFfQ3sWLbZBHErSOYnA5JLpKazUeSnIxtz85R8csItafLjjq9IgyRVzs+
qcE6X1EGK/vfKnd8SppvFzTMQKOwLZYM11fNODUoyMgrW7CCiv3kP3QfvVmxcHfL
q4warFpxadAQRHd6YktAO1v9Vs517xUsLa8Wutbn3feA/71ZtgIfghKekdneQHSy
Bl5Uyuhdwm8yga3OvwpJpcs+ukw2D4+lvkyYR7Fet1YEtOy6fCIUMc5R1xPP+WcV
yTk7KrMwFl1ej79Uiq7PNIgzMMMEl51d3e52ewXCoNPbr1Ufh5GBFYjsrYRq5DUb
jB6jgTL4g4Y18K1JnyR7YzMyIpficO7pF8X1hfYJiobP6N9Q0jPTp/dwESs6O71i
CKPXzqfXOq1y0hfiam73ZGkFJ5QEoOjmZH3oiXA6KppmIUNca61PxCtlwfq/8T+/
0Kf/B0y7qlzV1sJBJxny2/vACPYW4eR5MjefKY247rh6yIjlxMKl+MUf9x2IIY6P
FFLL+kYN6yIw8hSd2Lqw/RU1Q7rauRmQnMaF1sV71DYGKu/N12tXVw8MD3Itgiux
hL6j1KhAHBs8X2aA5pPgLNgRad2O2JUU9VmhubwRElGHoTZl8+BWHZU9WWiNNres
3mhO4/i3ndjH6hIeDyOLPkcQR9fYD9s4oi9XQNVDITm0Le4hEhgVcUzFVixPDjTo
OCNEQ/2znue1HSSe42Fk487XxgI0uezZxAMQf/5wvUyhQappsf31jKCW3qDsPGjj
SpkO5ETU1V8t1tYtesqo/B1hQs7lX8DfLXo7B2YofXO0UgB36N9n8BF10MLKlh1+
gYd7OjG6zD7RWogO7s02pjReqCqzHVTZrUximnLVAJbHo9i6vJwgp8UFhKov3ulc
F/mKeS+ZPa34tMMsf5Q0zE5M64mcLFX7M7J9M04YpZ6JQaZA93A14UMe919+/tAH
4Mm2+WHn/NNg8uJ3gFnrt3a7BQYBPVQLyRC0jZcEzwCpzrPQxWMhdIJ6qAhxGdwS
w9dlmzCBpTVVArQMIEHLpXErWKgCe8MBpf6nC6s2XQ1Ew2C19CTuYL6h+ExWFM4B
ZhmTRwUnppDHG0NZT+vfdszUPaViOHcfV59mi65tfgHqorMj3bMOz3+yX5L1b0d5
MIwtvXsFq7ZJyV+n+giGx2HUA64TAqfn57ZZ+aiihFwf2eCy3yYmGiZzHpuoWrbj
ak7KTE0Kj8TZDZorYRE3Z0jbHSXjar5yjRq5oM68TaGyQHehNT7VezqcAh4hk8pK
AxBDyVCyXgL8j11KMCBoiEqJ957FRKoRShEczF05tVld6cWzJE16lv4oLbBXpjvo
GJ47N/FFhPMwgNYAu8i4JJwWERqlt4Xxcyj5M641Or+bD68RtlFoO6f9l5lIMzbm
IvHm+pxlXijDKoMjrz0inSViDMtLiNf8Y1c1gpNYSZYq4rjpf4IOPDrPqfHttjga
mWTQ9YuNdQM6nrn8ksYH6cFO+mrFLqUFFGWzPTNKRgLEcknxNDGXWjOGabm/eChX
GDsrG0O4YOIM/1G5C/NABayzb1hs/Br4UgC++4mPBPLU0x0UOgTEPUTgyjSdB5xB
Z0QLluyatKtvrS/kwFTXjuSGqWZ2VRNIlmQwuHCjk/lr8tZHlkFiDm0WlTN/cfzd
4LUFjP0incLg3teMhiYrT4hiROX0P0ede6CodsLnKp0pGswgw0PYhywtYgRMCSaj
gm/Kj+FyHViwxiaFlTT8iXJNTIKoRcBF0P0qL/7uOqOri6QEYQPpoRTGjn9Dat/E
6Lhn/DGiUsy4FNnstRL5MXOB7vInHXqQbrQ6qdiuuj2V8H4Z3n1ko0Okqwq5/F42
tDXQlytjtt0abQxn+uBJ7E2SCoFtPwzvz0VILkTuFfRNpWHmjXAgop2i1S5RthFS
ZA6cRNwdzDRJsfoCFkVEXcSCCAS7VbipW1ZgH8Nz71gV60b6X/OJ5Ii+QUX6nqEI
A6NW1k/bi7wz5hL609TxQBe4Z32fl6sJVmx/OvKT6fwWjQkqXjTSuw6EElOVdHOw
vHKlCjRCDqoc3r54kXcZ48g2ZKpWZ6ZocWeYIp93sBCj32JB97GYDJQq/pDbNDkl
DWzbNKs6u0bvY18dcB+w06m4rgO/Bbzcxab9RuxAWE9RUtmIvbuG1IS5eVbgNCTP
eXduizT/kxSPmiIG+KAVn+8/r0nhgiybsjoKLSAUhlRmvocYXsA4ymWQ37qupmcq
mab3juXcsiqmwP+VFLgYnc2tjWPd96KUKdqBkcIRAPJeSQmX3LEfxGNwNNeYRxxv
6S9GjDUlsHySmASD+vHoh0Vq/8SBkH/iLuJg/DuLVeB71Tec9ofmrULVIaEG5THm
M/N4D4VtLah55iIHOCo3ouWWKviEINAd0bbmTIEQX2ayPhgxwu3t2yo2KaqZ8/cQ
jAPI19sWinGeldu2UxqISTwOZQwgXR8ISYpGbPwk3YEWs19LvJ04ms8+zuBdV7Jp
ihRoHdAZ0U+u3dIjtgM3YD+HpJ4na5w8DzzEgAI+RL0zHPwWMh+Jv6V9dG0cegkR
HvqZN3fqelBZooWJAm3c4Y3oEMhtKrCjkAtRHh7U/qhCyd8rzEeTtq69Qv2C8WBm
RTyOX2xnpyNLqLM8YiCmn2dwPzlkyecGNtVFkn6kNlf3ux3T5q6J9kJMPFDXNaze
LQ7MFC6PKl8JH6p1dfLyNcTFZgAnup8Fb1cZDh4luRckYdT/aLzMYSxLzOdyF3ZK
3mmhtW+fofQjgCD7SqaZyr1CL3nKdoPvnNC+MuMDuoLakT0pVyK0S4VvzB/mRtof
Cj0GOuKo6XoS7OYGAww2a081dRD/ulS4LPvm/i8hhGIwyOaJ8RmwQWQSktyjJ+bX
NPy3bOtqzKgNLDutbeKtL7fv6cgmTk2uQj0WKO8VrQoEldmdgekd+/ljpkZULpXR
pmpo8I0vfXXnYtPfKSnIZXiB2+HD4UTlwFQcqugDXyz/iKxva8E8laYZG5n8gfka
AYtX9PKwgvnFyNacZm0uPBlGiht//+KWr1Ofz3zeF2IQXb9iQmM77vrEbjL3h7Rg
DbJxq6XSvB4uhuXiMskPITvuC15B9sQ2TedXdUqyHSNq6M9cxHHhktQBa1u6XkNo
qnP9B2Pvp+FRQtNoL62gcExDOB5i9TWDAEyiEGTSx+waIIQnyJEXCacpTQoHf/Fz
0Fg9BYI5CUesz3IHL8PqFOq8Y4/eqSNbbdRi24/OsgXOYk3wymU4VwoePjZ6PEnv
MV9h0cWLeDDq3fq7tNL/MeiRHVS2CoqNDFQ+MYSxcPfFuk4WiZcO8yHGAwKbFx9V
29H7dB1dwkstcoMy9dgTIfoR4C6W8BAXeyzMBzhD/aeiKk2YgCRd88DLKoIgGXvy
WeGm9qsZ1pRWf4PnsimpU1JZe3ZCk/xXJUOUJtuaFjEYLwiIVoUgdOvyvm44JQbe
Q37LjIcJEejj9j+GPlis1PjbHaxJ/MVieVLhTfAyV5JXNudjeSlwO8x7M+SXUTWu
RqmiXOBMKYOJbAM6a4KPZmxpTFxBVpe9xzM8QDw405n7IbI1xIBer3p5rwoGbIxQ
vpGUbH9k+CfdXufLnvtf/8hHpWQx6GCpOLrFzk3huKvpAWOGGMYbNG2jz7IG40Zx
urPQ5Vcjs4WuSJfrbwtzDam5ezVkk3c0bNZWGaSD6yEl5/uy4YkijCGbPKEPVGr4
U36oYt074oJ1HP4kYNBko4sWoeBevp4rmv0h3S23ji6MszYkxAFqWiIBON0Y1Vna
S/j3EPt6AKhPdIQCrhQ1bCP1UN6NUZ6SqZoQB7yPmxOhBn1hGTrYn2gLdvgygKES
CbbqtaXp4s6qV7q75o51x/pBuKkwv+rmCIRpF7RJC9j009HIC7sz8RvCfnmkGWZz
aGEibEMm6J2gtxEAH+31WvvS7lRfn1RwEUZaPBfxKp4hoPORqjKzanLotCfWsvKB
8/Bd4bLcMK/v7oiGfsdYPDTsii/ZWYGd5H/z+QxiHLsOZTmE4C3l/nXUimdy4Hs4
ODDBO6+mT+fCZ27rBl9EZpko6qLRVST+daqB9UKOK9Q4e5s2yz7AjK0Q82idWyJa
81KFF9fJxYfuza6+YF2dyQV6rPv9pGJ1PVKi98h22uHykus9DROZ9LPXCiwH/0cX
r9tf9Vf4v4uld6l4TAynyRZRNXYs6GK/qoktnOjJKTUc6JpC0j0YTBmBqWZd/l8d
OuT4hbsOo8Sgl3+WHG+C9gFalWzEsIA9CX4zZbyqlnoBvNvIU6s+gQsxf67K9puU
4P/QGfy3shs/8M2PhsKe0iHHk2fe/Zd/c/JSakQY2cA8OznwwNT2hhOFnvO58X9D
sTD11ZE5c0Slf6zorCSM/dXCtFzm2zQWpYbtc0wa5Dz13Tp4kZmKSsiTflJB51fu
gJm1AAC4+y9T2DzzBsQLL/bYPnz7aBzxNIxCOaj07SwgHRzTg19AWSTRwpDZG1zU
HDcJs2bhzZyZXtE3gZHts5mTTawYZEPjcFeITDJaJiKCc5/c1/2bxPseEqN2Slh+
bvx58cVYw8qJLyCiICX+Z71LLjuYZqfxdHrHxdCgEeaqs60u4TZto9N+U8I/d0yo
yWQgERFBVwApCWuDMLNbsX/c6gElIEzRXQc5Lnkd50heqF1YX86FUeuGitbHiGnP
/JBkBOJusU+/uS6+8V3wiwXJxYoeo6UHw9uDwTzo+iyKl3s975AgC8k7iU2lXsCJ
yLLPlCmeelxPz+K3r0RiW+2tSS2BFL0vxNMjUOcyUzgnaUVsXtQqwZenY/UGXA2i
BXhcwK2KgzrqLzYZ/tHoxohR+BpPaeEPPf8+3P1S2aM/v5oKWE1DeXXALwEqLfRM
+Xs89zmh0hptlRyGkZY4y0sQhaNmCTbjSqQEBHhqWQoa2vGqoOJwhx/Mk9NF7xi6
aoYlNIWuJ/cafRo/Bl+ZpLqnJPbbpQY/wBJ33xMYV7mjEtNP0BB280AoOjI6LhkD
cs2Wt+PRny+S+RgqYsemq+1Hx0SdYiUkDmWtAJSYQFVYRpUJ56iEWjdl1/VI4dq1
pqzIZAZ6p73nSVunAChX6jz+OUAzO37uknSw0PxTrLDcTtgttznoaq2+41sO92nu
Mosj8R1uv79XjvdHodpkRAf/3sii4NHHJQiNX7nzmvbrRIPzJvtHw1FC1d9RSr1Q
ALcO/g5DNdVh7WrBGZJuRn0t+QQDEgf4XjY0KRdkcvrONwLoFdop0NpZ5iMzOhaD
tGRlzXZRpQ9pMZQALJ87CjGE889YJN23aLQWMwDx6Wc40RxH3jTf6vmHowwthXBN
7fnH6LBt7qE/YPvProRPvGp65EsIJcK/gzizddu8XKYNH39olxuxoyLP0DFfgDA2
vlj/q1wSghjXOPO//JkXkIvA3T/rxeOXx52zxCK3S07DaDbjYjpn4U0jFcVxjKFB
xa4bfMuzRl6E1Pe3zRSlK0e2ZhMSpZAupmCQI13e8OWlAzsvPrkbt9ywHeD1yjtQ
ZnlxDCI8Ivd7kHaQIu8m84b0aiaHhEVzC69/pNOQrpTsHHRjV+mZVC1+LAlyrsYC
ZSKPWCgmAUf3TOINTdq+lH96z/6hvpHed+xOVlQ/xvUXvWL5uJlIOBeCuJqkv//C
Ss8xuhDKEImx/a8jx0MPz5npwd5UDM2b1l7yAnpz4qQoqEX0qohUwDgJFaUjWGHU
8eurZS2PCdMFxqrUGa1tigD2eHp9ObzAE3AQkz1HSpaEDbqH7eMC+gKL4SjcIjfo
kmFTgADueo55fgyR/+QkTAprSb+TfdRRYPwq0RRt7/c7do17y9mF8tic7L2jpnql
/J3MDyshO3LvuYg/kbOKf/h/rUPeke7VSLpiNRDf+yt4L051NrovKsCrxnIc18rn
U/HHQV9/KYA5h53sThjMpfXL3qIL7pWnDtf3cxUvtqADq8oCiZFZBLwQVtnWa3Bw
t8vXKsuTLH6SEQ4CDRnUwDRbnRmA85dCfo0i3dzyiaTnQgcQGPdkNWbbGQsbOai7
twe9kZsv/pGclxgu+mzaWfGuBDmtlgzdUj9k9EpT72tGkyaknnOSJT0fzNhwmExM
lp4TZj2ZBMQAjcfj06OZqhqj49zwbNTr10yoPu4xrfoncCK3UEX3SJbqm0c17rM1
EIZhuuRvJi+3rzBXeRDC6bS88rEooVN2LdNZSChizZ6GGKU1JU10NUcV5SZqKt9a
keaSGXwAc43ve9gxHrs2WxHSNG/AljARXzbPPU+lfqWum1o1I6mpF2oEIqMq7LKe
VT/uBH8wQmg9vq+ZJQOYb5DJvrUlhbNxJc2tiq2Xa88fP0QiKKmvzxhaC3xtYIej
clPL1ENgXRBQ6uyVGUiA9lcErd73XIWwa9wx7q1z8asskeWBT3dEgRU3uhw9rVLA
mIag+nmwawpPgNnrlk/wwSVR23N7m71rcwqYHSliV9sJSnYsCFhEQCia05v4mbTR
OPhhDuDRigDta0ulZ6HVhkHSu0YPjcn7MpiiTYbPcXJAHG+DLIip6OMKJYSE8Xwa
bgwgW9FHNh7+jPVt9mhztPsaZ9m96QC08Es+avkKT6VXnDcoP2+eVUuJK9SNJXWJ
+cXj62CPGJMeZAjU/UGHQrSYlWGUappeSjVz8FtlpUyCcTwupYsqQI8kdFFYJzqt
1/qiVSvFciKgk0GoskvWdFWW403KQyloyR3b5cMmxRVYUryuO+WAgBhRs4ppznyv
Zm7admMqwF9NHYdt0zSqIZBwjOiNNNNi6TqQbmJmE+d9Xm5mOQr6ONx4y0J5a+Zb
sjV63KI1PpeaB9KbhfukP9PaD6rml+AirTAMyrJYQ/BueOEgt9zWxlk5/3VTcQ2v
Xf2NuxsWtH8tsVyR75HU+jzeVCMDkj6i+ndH0TFYK7xgs/A1MCzpow7S0SrRonyu
XWD25rZn1oTqfaHpVrI1zJ9ApMyoybektMVb3YBFoIv2nGtSw1azTrm0A1RC6Kq5
8ztN1dto2ubEp0KrqQ9dAnwWGao/wO06j5Ioamu6+vtAdSv/tkSq+TDN7Sdh+XFN
r3TBiXAHQSGf1NkyBQ5OsKRBRRnC0QSJ6e+ovBdxZDW5fWdy1uzDI6RBJaUUZCq3
281lJLUFGNfXSMVJLONJskc1W7Gz24Ec3YWuGLF+oTX0FWSq5zw9w49U27PjK5gn
Z/6PVm15RicV3cAS9BYo9+VyE3fLCTWkV50wPxiHH41NMXV+3AWKp3bVoI9c40hc
ZixNpiCTTwOlG4M4gB//20mu5cYSTWEzeZAmUZ2rozUGRMQwNYcZtDnQQ0D8O/Ie
X03/IAy89aGlQikER/+D63rdIetHg4wMFthrP7ozSvyddYVelNSaYvT0pDAMhNCA
SD1mGFyWsJTQN2zfgHa5p15l8ho4F4hV0418uuKWLYkCZqTY3fDz362kok/7b9J9
2xa3MAjfjTtT5cIoevWt2b0nTC/vw0fsdk/8MSuBFX3wZnaKgQ1FRqwDbcQgxdOH
N8LpVc3sV7lw1Zw3M9mkQphocGWUXylodqAPFekTAfpTxS6Gzxbs9YwmTBoNE3Qv
i7qMtutVdDMKFsDHJkcFpT4GlchcelQ/yZhEhebd7xzR/TeVVTrAvjCkCDONdBol
/dHLAfIv+j+t/RTE8bD6jvitDb9cr9vPguQvYDNARHYUxWzrD+5nwqroOhueCdGj
+nthDKzk3Brvwr+9Zlu9fmE1FOCLpl+ypxZMyg3+3OUGNfLrQefF0bTp+imLSkJ3
zLLwho3a5wUOWW6tM2ypkosCRvsmC/Q/Ok5CB0VjX1KvHOvgdq214cVxtL60qK5n
syAjQdlnmVZlhCYmU9Lvh/UroUq39Z1luTh5ujpwwoeSDO9IiRN+miLNlO/efI/N
dG3xX1RgE1CXY/8LBsaAgKzMMptMzlg3OcNjwN/gk0UhSYLoGitaoDnrYvwa91UU
WGsWnpmWe2NYwispEp/+ov0oRBLG80btxrPaqd2yRjX9fbt4nlnyut/yX2t0PlHA
ikmeOBY0SrUReXWeLKne061U6JzxoURZljq5mmvhIDKMhva9Es9fmt9H4AkfaLxP
KGKSsyF6Bhl7VACxsgGQr6Hmv9t75qaCh6vvTGRrcang2wQX0BOhWMniE8CegRw+
oNa6vAWtmoXbjNfTHUH/ZAjUWejjDz54SRUmP+KfKB33/HBvqels8eKIGzST04S4
536IU84kUElR2gBnkNVF0yK+Jas7chuaeupOXmsIkcykaiBgNrSOY79/sE34Ho9t
rlTTTwTfeR3S122bovR6neE0/z9C/4tF1mrt9RfDjACye3VHuIVqBUrdp61DJRQP
77Bx15J/UIPR5gI6ZjyDDsXkFDCyGy7FpYYwQgfbCOOvr5L5PjA+0pk6yuWgbQMw
wmcXrAShf3pRSrTGehr/1ahSry/OkuZubFJ24wfr326hkxwK04VHeY7umkDynVmm
og2+D23AJlqGc438RzfF2zhXfQ7r4yE1tO/njcZRX0PoLdqMcPPyx4SYOkobeDFR
aDoXNFWRGCmi409GwkYUzbydpEmi86/17/iu0fYmOffV5RXQY7euNHMMQAmd6nR0
4HP3YvbFX0D4F9UP/eALKoIfWtcEYr9yA6ivlWl6BmQtLELwETXO4LGfN173z2fD
ueBjZ1DN3WOscHoVT1UUx93QfC8vmuKFMqIvQTobWefvR0/6bMY70DdFcvfSTwgJ
6+x/K3+NtXv2Gy8I3v7vdUlP+JiyIB0hRef6uS1MAA5yqST8RYqfyn4603UerSmT
uGqDg71yhoM4DPibyfSz9M5UrGIJtu1mGXL49lmWq3W5yx5xjeoGPptlWJ6cRPqB
LBiBP3PPfEreJzrLBf4nOxpWQRnpbY6OoYqTZjDCyRxbNFBn77olIl+veHIB7riU
CEdQZQsAB3cAwsBFuZj4N5OLcriMfJPcYOJ+Y7EWLN5wFJqBRj54q3Z4LT2r1KHM
dG6uaKiPcmwp4Rrs1MeDDzGTvO4BVLuTUmjdLptUZund+v3uur09TvfRKs3oXEgT
IVi8h4jDiaX1mZzqkk8nY1uw8z9U3B7gOdlmV6Kzy/XHfqM9cm1i9dhe4p4+dxzR
HrFaoi3mYRgA0eg51x06Q+fmfbJ07PLFGlK8JxBSE7YMm2tzkVnwKPKL6k/7f1bx
z6yY5jK3U6myXfG0fkzRXn6ybeJYcHG+xcK+ivnSS06gs+4ROHFp4HrO+d++zj/q
f/06FyOFlZBPKsL3aMNGLXLUZFiADAhMh+6KQob/iBKSP1uSyZmZJOXhQeEinl46
qP773X0JTBsFqmqjL8HMwSITrU0xork8R4V5zuSXM5NRkeZu/4Ba9Vy/TAhh+gLK
z1zoZ72D5t7zAzumn9WoSHDVyByr9HFQ4wiachcXHOXCMQXQjVnl/YndXUnffddz
6sY8wc57h4wPnqb1lnqSMzRDN0dqUcZGWZvrGUn3VwTAGASNyy3ArFHy8gIO8IeZ
SdnTKx47Xf0GkUjAMcobKIZ0u7VjhlZLTPYpJHsmYTuqyUJ5gOeZ5EQwohTXFJDN
e214l1ga50RwJxull7Ym8SCiaG3dL4Xvau0PAIAvrUN30G+vonT72HYFTGX8NVBH
6Er4rVFCNgCrSj2TIrJnPnnwf3UlKO+RJEqms3ZD+qa5hYtfC0A5oQ9e8mHiDo3s
/mTuXigxguEdmbkssN7ZuWqCXCiM64+69VXn3kX/SdlTnmTv+KnMpIYRx3ylPPo9
qH1Oyc1aUwIgc9pevfkpO2n9NhktvtvlEnF2rw/NLtdQ7lw/xmVyRBEtsCZOkaYr
6gTD/Dl+b6tbydFs988oV2O1UlysiOMkBCRXPnP0QfpzV3B/FksMfcbdrQ0lssVM
j92ig5m4sjlEbjblvyJW9DLRR7CtftdUOiOmvu89Jtm0hXAur+7xXXvJ/RyBUgSB
KabFc1tXxRLuL8Azc3najMA9akFXBqoGhz8PW5Te0EPonK66+QqQHRml8SM0Z/DT
NaF3rPsp5XCdAAJz9e04kDQ3iNSLBhMO3k7j3c9ah583IoowigjGhMqkTSt9StPR
sLy8FvZUnYZ/WBEapvofBgdgqwEEokLV1C0YIl4wWncmeLU3+fl5SQ4UBpUEEeVG
cDfkv6CZVTOmQaYs4kk4czeKZJFiDC2UIVkriYlzHjFFQSK1HBo9RQtyD12ZZcut
3iTya3QZ1iexjq8zXb8+TIAZQhXihNumoi4q97KDYiYZiaD9jKS8IaGCAUJn9Jld
IPcGxHiaHNs0iEOpDyPEQH1EHtli+Og7EpvDaK8uVcxiiirtcrzLKHynv08ttgqd
hQ3XBVmkQa4fNLWcHdBLRZ5+98vZB6s4SDK6psABCEnBFLJoNCloQBd07FSsUYX2
9N+oGxUvoYncEktDGq7MbNhr9Bgqj78Pwmxa00kPHfNNxnIIZ4eqFPXiqAuGmnoU
atkOeZDXX/Ij31sRK9b8b4U74hD6XD8aYRq+feq84D7xuxAL7QIzcmq/HEpomJfz
m9PRBfZ994+g45TX3pPPovzxA+72PHRBOqFxkbDe5CGsSj20hwM29crqA/1qT1Zj
ZPGR/JG2qBp78FDv7PGijZCKrewcvlV5M0Ym9rJJkk+Rp1zy8yyW9U0t3JQ4zEU5
5ENH3BNDOnlLdTsqhqULGUzgvEGRdh4qfq/mSDjo2gDxPPyYNhm9AQ7h7yKO/LTA
c9ohrfyuCK5a8JLWEYNLv9ttESmGMVTvlb0NcYi9T4FgpsUfbagEH1Ew0X91db33
/4J6UtRYQXFlpw/GNzboOxAVY9ZFvLa/4+8IRCpSXk3p6zUgxhdP9PEQdEIp3vHo
NBMxe3EJnvjpWl0XKOwHCeZ7DvpMNi7KqvPh1oP2QTv0lrQW84JZbHx/03wXfY6s
7nvqK6g/xLxctw6e39qc5mQDEYnSFc7vsE5my1SlKBrJLKzSKc/c72FfYC97wylj
hlZhg1tWD9p/vy7FegfTcsgcLXHHNi6UWZVgC7s3xcvmMh6UF5WUHYu4tw5tUJ5M
T/FWFvNY3Lp7PWqzrUI4/lq7a+rJ+1HmIFUnYGcHPGbic2hwVibq84zEgjleOpO6
KtzeqtqqYcMjxt5L9ed1XduX5lrq8Jc+ELaaSA6XRd7meRrMN+udBgo5VsdoKaA3
97Dq50IFOH/z0Fx75AARxZgBJkJmX6oNYyF3cp62K0KJ6VEeuAZgvNZujLsOW/0F
ddsXRR2f5NqgqDtgECBugGiLqwd9PR9h6JeICP5lNI0oelWdnvOQlZvDQODxiu8L
maYrmjGVKS5tKAL7j0s0sib+bjwMT2MsdUXqDnYBPDpvOY9bC6JMeRF2VP/XBMyG
q6tsruz01bUN/3MTsrz7lVWJkV+bLhvIVwAgH35Q4uYQQ5VmCiuQkSsFkaiEqbuo
jJs2Jq+VsrHDAY2R7kxZ1W+jF5FTY6jRkSiWMDMuugKL+qiqitmvi002tg0VqbbZ
Elh6mfa+cnx3HY6n1cWqBs2ueKC4zaEtJxDGDDHCFhqxYPb3+CcQsM1pmmyqv9Zm
tKkWh8LzSk48h7RkAz1Fc82LLFKCeWa6X3cvp5hHVgQZ1eQI4LKRL3MfndLbzyxt
ehKnQTwzoKJwQl4knXuntaRwP5+Bay86A19Spxw3gxBz/+vzqjgMGTY10iF3/O9T
JjFEhJiFl3fm8xaQocXD/Gz2A8Mq0IoTrTJA3z5m1g2KbrpRUu71REOh75qpPCh7
hTorvesrUsjQBW5HMXf3gR9e2TkSPVET3SuTkO4Ya0NVWcDNRkBRmmdAdHfcD7Y9
jpCVqAjfG0U2OFXOEXsC/hxssqve0ctMUE7AmU4GEhdaegf/UguAGxjfJZi/vHRs
keTvOdeTvkIhdr3PtXZ2WEiGyADaICCm4/zKPshjyBuqOIcPxR7p9WiwNe9mhSXo
mk/VfnQGYUdxq42EiLnZQGJeB8wdrv5QHf+e7+8uqzMaFABhQpHe9/HCpMgHrWuF
9RQJlR2Fryr9NUcH8Kv7jutv2QD7EV2gPslIpD3c1Q858VClb5WbDZE8Emw+OPpq
IEN8zZ+8Atp2/Dophg98xhITqSm6U4/3WV6i0d1wWMKqQFY9du1xERbQYHN12P/f
JYYZtDCONDdhyvintCEjYcpnZhcRmmK6JETtKVokIxkBICmCHvZUIZZ9XeyvR+30
gdnCGPGFp7ez1ZXuBoUJQROpXV3P/wWiYhG3fMLA4r1SRUopQdmqwJMeT2LqlFn3
VVUzgBgbfLcSAvGlnnwBdjYQgoWp3RVbvwYzCdXsZfFSVonUe9HXo8fo2WcNqKq2
TJsS+AzAi2W64WbtyMRo8+RnizBOtxFuNJ8IMlY0uPBv4WYyCa0g3HbOOqhfjeEb
MqLQS5BkdUhuWkRLYSk5XIwnltOKD/wOhr85/2KgidOXOuw5rZcV0QGny7w+u1o2
+GeqCb6RyNzseyHd/9vGTahsER24sWccvThBngbu0E0+/vJpxRW7SJnWnXh1NWHP
FermFgM1zFuhApHRryQV7oBkC9gMbwlI9kS5ocJPPsFDYCApch7AgAQxOMyVCjji
lPhtkrobMv3fLSEh4TSZvNL3VFRUIpx7HovWIYeiPoOHkNXUpCvfVEPmO7xySiMA
Kypk9aHF80mWGCGPjQX371B3atQE/ZIw81pDyePqAOSMUf/xZGMUT7TpKn07Y8Lo
bihMd62NfaqrnIfTx6QEiMna2gkPceAYbOqaXV3hLT7RvoUX8GBVx6h+NrWyBpNp
qGkRytj/Vz4Btc/IwqIhSTq4lrUR096CoivswkhteKJ5ALLp0JV2jJHnFHic5s7A
txx3Pza2ASmi0Xre8/AKvQaEG6B+ll3APLNYvHNygidFcDKPCGBXKkg7hb21GVFI
EuwCBhO/oJI+JA51u5kytVoWYKFYbnTAxeD/2sA7h0dlJTEGflvo7FX7Rg5VUikS
NLmCMbbZEFK7ECTWI39/MOP1MQtBm6N4dqLaQ34ZDZPssoEl7+KEGc/xk3rupBt/
ZQPwnS+lN6om3Tl3Wk8hbLTYPL/90ya9m6Hzf6aQKTC5jiZ+TOY+GIPw15FuN1k+
Dl/8zr69CLyRd134wzqhvjHWlB7pkoiLQjt++Wlyvcpe6sCVx+7CpWeOiWyyZjbe
Ut/8KbZdngdPwIWC2nkKMRO824maIAeWCZdRSsHRVTXF/vzEUrEn83ceeRq99Mvy
uRh4aqcLLTn1kkw2zYE0RDaMuZDNtaVMGoArsjawqqSNYH8sh1cRENqkiBe1bg32
z65aSCEndUaJtL2nzQyypZq5sp1ermpsZthJemBkriRXA5/rPlDGDkyT/KF1/S6q
5MbgbZ8geTQCkWbyc1oG+eVdcvFM77pNQBDwBcRVNzaQKzeTBMmZEQGBJ2dpr7bu
9FNTFUIJICkoV2zJA5MDZuuzlg5P28oLccacprBnd9ssWL572GYWbKVA0RMVCiuJ
jKKcAXAjIeDJoyryX6RA26T4fsOXh1oDZ+dwgNCo1V5qqh3ay280Ib38Q7I3+tCR
ttAQTCM6LqFDkDeTPmkR5JhYRiv371SzEE2PugD5qeAIGn1x37PWg+lSmWzXTNEq
TCLznOyZ0e+T1j2N9Pg9OXCMJVVW7z++X8xwJkpkOtgOMWZdi5Ua2AKrxT8ZvF1X
1JYFAkVSLmJlEMqTHmtFOqmlecGnnsR/PXUX03d/QP9rPSbj3q2tzsSsiPjcW/WP
sHrrrkE/BX8EdTJJWdAv5thltu3sF5bmB1QBmbzATTQClY0EmRBiBOvUGGbVHGr8
776Vhd4r6tGJzqZSlsIjH4wrhtbfvYFfejBoNdDJJK8g2quOoWYL6TaN3qeiZIUN
KsF86kNFwkxinemVJe57/+wPo42reOccPmfHlwGPtLohrkccunVyntrbASzg1bjf
wHDKhzUP2RVxZhO+RXL/opcFAQD8zuUbstKaf1XWZeZol5whKRLtL7tu2WnlkTLe
guOaZX+kfPErSNEEhvZl1Rv9pltEhQ+gDch/VKFcQOXxZRUFuzQJQfjzblXIPlmO
A81bL4eTOGUMzTMzn7/H8c3bGRdekY3/4NOiUw51EkGWkK6rV0+osRHU2ajTFPw/
CNlcJZGdQRk81dnkh6QAILiwYZczvgx2QRetzHkZAzHzrWaoxRDuLNetgXQ82buR
FQLHoRLItTpBIkZYYceSlBLs2I8xoj+eWIkP45Xt+8oSjSl+VRpQgctQYMdKyp5z
2IZcdQrX04AbQVkkzEWiLHo/1NpbkjTGb37kvQ94OD3siUxPKGCMMijRHOjbprPZ
j9T8PZyasE/bLK2/uI7rzyg6qp400IgeKa2MblDYu70tSRoARNl5x9E88K2GbuoZ
XYFHSguVA7nZmxJ4Y/FelebW6myyb8bx10XP0AeD+U3hF0WSB1xw53HPqZ4frE/Z
2WAnHI0mSHfUNLLIgSgETYfYBg+5pRitq+2xzdqdjbh6XlSSVUUcp2yPUnVWODkX
BP0lOEjPFCcQw786MzFeLqiBUQx1j0EwWI32T2b0F/P/dxDX5mQ+uo/4kWF8YjSp
x41uM2BwP6zbZnPtJ7jb+44qoXd1l4oEccideLK012pcYX1YSWlDboZibRUL4Vhx
fMAckuSpiSw8PezSr4ATywdmP7vJGLKOy0nZe2R5+hXX+wxCkRaiEwqJ2S1QW5eL
Ai73QDAUorw2qQ2CNzcKzmhSEgkzjVuWIBYFd3lZWY28H4Q5nqP0Q8udbs8KQj7F
RzVlZ5N94yyvfHETODvBAdzd7TNArulyCQKMnq6QSKOHNmznPVbN4T8MFgc+wGLm
DUltKtSi7yCUbwrcXZSMosGnvGRAdFdEwu3/hPnm1G22xpv7D6ZAvL6mIsiyEgco
pjsRSUMMZOLvCa5BZkMfcaXUUfOmNjYIg+L5ODBP7Y6DHedLp+dVeQzfgwZm0042
JUEKZH76VXZcguoRAgxVx3OzIGd47s6ud9Cl7vZTP4T3Ta75JsxyDgNWLc1D2Mew
Oo9HDBxxH1znIjax6ZOsNvNsUkBscBYb/4HoUPRmqUgP3MSTFEm5RUCdzZtH31DD
tJUer3usanfH8nU7Qw0/ifQiNguNmfT0j5HZZPJ9Fje8HM/9Opb3eb9cyY8ZVlt9
WewbzMMFgMz94UJdL5Lk7rX9nz33T9/Yo2+VO+b6UpuYMwBqnknPbzdBlThmyKOS
FHucFHKBEXpqCdAVppqRug/1NgXSjSykz2BpxTdgRlbHgs0+Uyk9tnuP+oC6ROq8
6KUmoJNz9O06kjGf8Xl4DAzwYMB6nHMxbt5cRKliUZCRSfYWEAIAyW0KEd3u+akA
FeDBmY8EhpmEeFR59ZarKBfxHoo2Bjy1Ar9wBM8LeuaIspmsMbYHOhP6DlzWGnZd
4ait/f5vg637HvL+l0FA52+tEyuZL9jrZuyhuSz4u+YHhHrQ8lVIe2aRGCKRXDqp
R+LsQS+XUVWxpQXPkOhTK9QA5ib8Q92bRz/H6kVy18hM6o4ZGmKY03KjLd4mtNIu
FnrG+LsRF5UDS9Hb9STVxuctc5YagyiklxrajMca9o84Z3cuplhguptqTW6a2Itk
iaEkhFKQPgRtgSjitPt+lL7oNDQ1/Xo3qx0r0mHMb/6S2U9F7jxlUYxUhvKEvJjl
rRyI/U95mOdgxczDzj0iPaONbfF51/ZAHuRNMyuhzuga9S22N/4cEjcr49KUVEl5
mL5f1c5+6ZOhPk5i61g3B7IcQBST+t+W9KAo6jLUChargd8vyo/W4W4bGJFrP5Pz
l7MQvfXLMOFyr+PGRxJPDVPbNAABESwMi5WQ732GKwV8yHQ43wN/xBnuo9TIDf9w
eY5ezibmDgqGMTp19SZlinK7LtxoylYbL1iAF3cS73Dqq4AHz/5R9dy2TQEJqH6k
wdwoaFjkDrRO/+U9KWHMCJ9rg7+aPi1MnV7SOG37pi71Yk9ZlSyqFIbYUSIEqb6i
3sCWQssqAlc4az0F7YGYZnInqmL0w2ELUPFwvGQNFr/iYV5dWqn7+fFvumR0Iwl/
r1lf4jyw+d9yxpMgwQSl/MfDUpNz9nFJLArTg8Z8PX1NIPLbOHnr1quQzYFOrJ1n
8uWaQW3PqVASUBZWTkQtaBvRoyxrlx8nVdNZ+hyXFi50eY7H0yJkdJPCDV+Si4Uh
3Z15tzpaNCe4TP3qvKwqD9ZY88PMO/YW+5Dto8v8lILlF7SqDcqsItMHRg2+KDE+
J+CKU/AU3pGxFmCHOi9HOd5uZeGHWfQqVF6M5IPDfkM910ntaw2TxS+ue1s40QAc
RU879+Jk/lhiFsYzg75aXzHxkcXILDtvPjGoc83kB4eoyzZNVGIxvSqJqXy9yWzd
PqiDEHs1amNqUT7XRGqsvOeyQMloTbyoxSB280Esg08m4w/CbHFK9b5+ZWA6OQdZ
bkiSs6ljot1tTjercGfsbo3P3iAz65juS7nBs6md1FypV4K1+yb2pCGVnJYuffzF
kDFha2WKwA9DLUA4/Px2atOv8oqm9uS0vM4HblFhfvxL4Z7jzhgV7RTV/C7RkI12
/f1JO2qN14A8PbUTVZEZdklJ1ju+g+BfV98OR8xqJeovPXFAkGWtJl/UAiicRDiq
xev1tXzwIhPLOd6VhNsJA4OmVpXz86VRsg9CG/5DLp8Z6VkDlGUzCWlQIk2UcmwM
cE7+PGzvFA4hL0uWh8wATR5eQ5wLFjTeTphLx7GrE0MILg0/kLgo+/GeMyQS649t
GWMN/x0K+gl7tDxLiLd4s+SC9GuMfflRr3pZZE4Zhh3P4BWWZ5we64LW5sLhE8H7
8fuuSpdI2r/FV8wN5bZnh0yWxEQapxt0ELme5zc2TPB10HZJqO42cqsBvZ2hNaU5
Zpnfda3By3eZMCNOQ7sAxe5SIWJ5MyTNJvnfoolXGC3C6iGzqb1eriDPcaJngD11
I6KsU4HXzQC90llmY0BE/0hfof0ZcJLF/aRooHPg2psVurfzQHHFIjWCP56U3sqe
3sW+1vPSuS4LLf1Xi6TAhjPkvIlOF5flzv+XzmjYyIpKANKWUsMI7Gz2CvzVK8Kl
bZKh/DXbfbMFVqLoe6gBTfCQ9KHCxow5l5iJ1TVt23aIbL2BnVIe3WJJKs/mZxXh
UasYg7z0OixonNhb2sIqCVfB6BXiik+Twe+rLsiCy11+i+tjypaoT15gdj5a/811
ugLQr7si6l7VnL8rBmhk4qkzjCiXcTOzmlnER8a/z1xoQtAuLYu4GvVBKRSA9oae
b5y6RUwwBbSct8ThrtQsJDk430ahwL8LOyMxwg1l6A2/cIOHgWUJkP7liiN7Dwf0
74gsW+DwHhOWug+MLq8Rx7EokHilHcqQ52pSVG4QJXtBnMaZFGlKwm8xFKz/Fdg0
YIMhkccIKPHzNes4lF+Ucrr3E4/doSXMWMWcT9W0EZ+iruUCkyzlVXamRdHtLesy
MoixVeDaaTGKZJWx7U6edIqaYuc/gbsQ/0HTDTTAmtNo6V0r9QqgO2X6hGyGbepR
2/f1fOIHtPOSz+TJbOG6joMaereYsSWxSxn59jMGu7/rQDaMSWXrVaCpJqhrHMO7
gclnXLGD0pus+qIs2Q6amSN444HXYV1kq2GNnVd1XeZyOPT8gs2jj+mQRzYxfhcH
C+VXirciGXEkBnKF0ljU7qXL0MMxFvNVloBAmfsqAI2jhhy9A4UbNdg8pYQtkMdz
HiW9I+ZeBes2mBdh5ZoWnGt0zIExWLjH6DU61Cls1NqICjrk2qb4E1+coQD0Omha
BniKsSsdDPb9n6iDXmb3bQceBO1+0C/lxU37Ido0bWLXoGk+8q1vO0hGOBPBZLWv
BsANflv4z9pP7hm6L3aWfSUGM0fJm+baJ+b1Duiess23vDvbWQRmY57CDcFdEne4
iyXSvmoNrtW86mkrbZHTqfEpi2QP82pLtcQkBm3yj2PA6n1/ll3thSFXBEj0qWo/
oWaJfxZp1T1GWoORTSAtbcb2qqb8xoi2Xol+Nf1WA1j/ZCRaqAvi+4QeRJoNJC6+
cZw85yj1gA+To2yAmPPV6M1/1QtmwZVsxTz0X3FnJh1BdRMiH0elltdHPzo1blH5
0KLSxin576IFqdMk+AThHINrTqXrymwdtVphsvoSHc5YYoZUuw0YAyY714IEQeF6
rxGAEHm+l8dn6DfywweU0ViNFk0mCkPAeo6Vh3yegXeNlskzPI9CS0R49iUs+Spa
JTI00BkC0usY+NuaUE8esXhkMi04QHDq/y8Ax9rGMoETqopVuscPTmZGCRsflHGm
4Pm9bhC5ClAbMvjY2A7UnI6NFNc3y1t0yRXDsXc6baOz4lBXrqWKETxN903wjD5q
Ww94J9deBCzWQKdaLpPTgEruML6D6gBKjNuDr3pHJ9GDHMZYabWImaKbcs5RDLeU
J8T3ILTJsvy3sFr6CHXcDUiFpazxjtBbW2g312smsr6vwVybFk/MMYzY4ofxc9qS
CNLQocORwR3WKEh+D0Ku+vfhsrPyEqcNFvunTS8qdUpG5wEmXPMj0QuCrw5im1Df
GF36+QaPw1J6wdQK4EXtWpgg0X+toBNabj6PXtyTrhqzTct+hgbwEsb7rRyU1CDs
PF4/nOQ4ZfKhGqs/KO1kOZkEKf//Ux7XLt8/ILYRqdcxyc4ZA6er8TstGja1Zq9L
nEgMdJDEvmA5llDGuLIxNmMSvoQOHmId633LyFFMb3suHJghY5jggDYLEZeW7wln
mni+xNLZWZP0+9fJ71YxoGnVPNASEZqjDkON4kWj774gtnZ9yiC13tVXplZLLQem
XJbWusqlUngyzra9XYioY6rWxIQvFUqAhlmSMgpiprj2XGBglKGnxU2Z206KJp6N
ND68HQIJApzN0D4oBPJhtq146qzSsHmOLu4bGAU4Q+qA8ZG7dhJWh/tnZ7M0E3fA
CYWRVzPB3V754DhB9vtRV0MhBkFJq7neMdAb3+tQr3xwf+eBQuxOazClQLL1s7zJ
wljStp3DrdilUZ62N6HbQ74La72b5FnWgF28+2Lh2w4+7NSC+wYIIJK7DfOQXp+t
f0+gJ5JM8jovETtay57JREgRrinkz4T9dp92GmwXJb+7RdmUR4uKUld3mjRWAQvs
8O3H83iID6ntVJQgzY2JNJRyK0KX6ew878BGzhyKjuarSTsNVFz0ovhzds4BHCcs
8oOkIexb8J/Gniv6oRGE3wboXk3omg+ame+4AOjEvUePiDgwfD80AB+5FetAuLWb
n05dLxkTvhY2/5Pyy/w94RndCYKaVrxSG7L9uT7f6BGktoSfG77TtOhxbaSn+iCF
z+M/NVgV2YklBq5R/tO96k5iCZJfoee/AfuxzjajhVvWg5+vGTB8bhs+Q9OM6RFz
ahj6pIKCVQzNwF34zPzMlfyQgLSvN/WdNwva7p9dCTctgBNaW++tg/4yzOePjqzM
3/WAOiQh4ggHywLVrJKR9nEOIZi31J96v26RDe6E3ud62RmQS0dLyVFHs5ywx6tF
jYdMywnP/EXzBVdvyBfOX0c6isbYOShfX4ijSwhVGvnH6SwsPF+K3eI/Wxi2fIwj
5GIFmx9bcEUainSq7+l/EOKPo+LFbuboiibQweDCkZiKqjafugJkDC6jbC7bh/dN
QS4hbxo++wGa6Q0FFNcxm8i4SLkzplcdYwKalaIF6+ApcdWcrMid+2GAulrQnveN
MMDSBKuHtMxi9ho9CwvJLOQ8DA/kDYbra8r8zlXPZyeTUOOdgawoq+ywp564OzJS
m5pzHLWj9YfitPWjUpLnpixXNf3iyVT5crwJaDzwPc4JtabBAOXfUJGF25dnqNKO
Nk4Y4W8xPX2nYLZfZDwPloTS8JA8hMSQRElx4EMnFOz0tju7TSokns5TQt/UEHFw
MVNGHjR/74XRVL4tk5G5DMtdLuBi1F873MfyKUujHRSdK651vfsjor6/PaGDeEl7
PshIQitTDU7Sj3gaBZi2bgl7xDBRPFkMvpPk0oo2aD3Bx987pvCPRR3NBasTKMmB
LD6BTq70NAqo9Cg0oZZaZSCG+CSqRpCn0D8SR7/OMxZnDecQpvtV1OdjI1L/JO9N
u82ZQA1Q3xIqaiTCgtEzFTFRwduQ6+qkvbbrZ+FjUjKt88YbwesMwT9ZLshCHwGL
gpcYGtAU6AAE4UiLnRD9SxOINbjnB+hxir6i0zCeORSNbE9KlxS3Z2Da2tu7bPYp
UAHC8wFNWoVFuhSKVrF92ms2w5WzvAdsUGRr6e3x736UhqtZJebsnC8ZJ5vNX3d1
034Tbej14owNEfaPcLjClqUx/iis5u0uaJCmrOgpnZK9sPLKhccMwLaY91f7qd+b
6gw9TnIJPbGwXM01NZkNmCLqjtFpzUS0BbVj3KEViNjHMRBHt004l9xy8ZamICdi
kybPuAa89EeK6j6JPxxJc4d+qcW7m6rTbGjPfgXTWyuxsza0YYADiY2KxonjfCaE
Stivlh0Zyxsoglmm/UQ7zP6x3S5Om+14uOcdTruTyTrUJdb1M0566Rf/EjBcuSqJ
t3bPu56/uCd5m81N7H2rCC1jzzxEcTR0xaSmaISG9x1gypVtfZoe3X2cv3k9rEBz
mxnUfvj8pT6qk6X4YdkbzmKCOvW1qaU94dvNu7yPZ4rdIZP4sS4g73pk2vNRhfTp
Uf1l6rbwsmkV0bI93X2sBLKI5qycf7s0odTLVQvgrfwMbe1ckjK7kPP4hWey6Bde
T7FA39mk6+xnbwFphGrvai5Z/9AXwxxbBjsuMIa4FZ/rECli4z6VVn6uuip+fusz
HaPrmNEgVBL6B4MeYr0dBZ1aJ0ymtRjA+wnVQ0rHSsr19r9qtmbCemRCFTN4peNp
YuauxXB2DqMvGygGPe17uvx9k3O+c7Z1qpGpaQDMr5MLjPMciqpFJltMGf1I1WBn
hI/s2jT12lyM54N7ndxevuZgM7lj8mIAqnHbGqkqmzWSdv1L0byT3FzkTRBOolio
2b+S2dxGsv+bJdf7BEVGdqFqIhG2wlf/EL+Gk3h3fTu2aOkluS7G3M71nvJrgfaL
ujT75m9IQHvE3IIYp/NERmRM2MezQQZizFJGgAccWClD4tqgfUrIYbTCyHQ/TZkX
qBcWwQAmeDBUejN6d2jA7kkt6jDK18jGJj1RbosfxmNUtlCvfk76/+EuGOmnsw8W
JumsR3Osovn80etzxovTN8RjS4lmM1FkrVcf9I4XKjfXxAjRVics02+EqkamX0u7
+JxbV0Hesa3m/u4lF1iMFCYGBrbrYA1LFnk63cJp5RR7vrALtyqUQH7IcLjauBbN
NUpompRY8KFlih0N+6/PhwMUt3UyT4bFs+edB8K94hvJFcIIBTKTfbD8dcHgVe9C
+CBff23yzaCguaDGCwwZLkjL04/miti8QsvJ1haFBY5UNeOpH82zsa/3jbTxOdC/
AJB+PA8AGGkdCvinAdLZpSBAAGkcKhQKSqjaZ+9ti/uxkTTjSwwGw5dKNET8nYxG
bZEz7zY+z2Mh3Jm4Bj/oWass8k0Mea7tsaJ9yx3AZCQzhM8yx6TEHa0u3wjK9BVA
2d17h50dIabGkbLLA1lcUhNKlXozQxiKZzpMwUmn+iTZRO2Va5cDC0DlnNz9bC+b
PdMUrbtcgHdCDsDVxd1sm1UIAc78YIrhPVwnRguvkR7HapSU73n7L78aneecSY6U
OkS09B1bsE1inWv/RLZou/hpy8/i//+EceCLQ5VTmkD8DKxMvTZEOXUtjqPe+ckq
pJO0GmGld3xxJSOO8I74iYKOuGvDnNsB6xQOoidgNjBpl/uj+NlSRVQtu8Nq8TDR
X2hQSKHmODjvBlKHrcgkPYSaXP+WZQHiLDqhmQtxXgkj5PBS2mAWCjmWEpzX8m66
y94gZp3RDjhFrkQr3lc0yjkC0jhACFhUaJG0IAJvxSVDtM8WVTnFYabJmkm7PfAF
VcyK6bYnqS2LJsHCyjKfjXiVZRkhTKh5pzpN9qPxBU5SPGtbn3Juza73ZFvRhGw7
liukGI/JXGcnJbRGRLNiXHwywlcl/iJOgmAXc6qwL8Dp+yo/cpWGTkbyJ0uwdSMg
i+QfoKh66lx4S2AOuHowvSvBLkIBkR89oCZ5lzOMLQJ3+mK4v4e9m74oPljx3Pqb
FMSXtkhXfRzZyU8e0t3+/aWkPoVtLb576632TtIG8cVZJiUKBrzpQkAFsQo4miCA
aEhm+B6kK4R61jCM2GO//nWccI8esPd0jSRtu49c+lH/vc4iLnz5RNbLYFAR4ITs
qZFYcYHzN9mLtJToUeQxBkvzTiOZ5DkLkhAHc+XvnDifg4HXvUV95JX6ES46Twth
HeoXxtsVj0OBeIGEXYDNi1bGU/jcyKwnFutCMz3+CSSGLTsMcTpfljITiXShmsW8
WKRGf96b33K34bU36ctuLBMVfmoPNn4yK0XP7w7hgywxxMr5Voswfl6PVjvkrVdz
gSFVmoGLeDSTHUE7OI0eP6k1/5u8/GE4LJK3TYMB6iiqziZ6ppuftGDy11bEG8Xs
I0uS3HkHQZ838TFut3BaZy8jhLtjUpWZImxO35aPEwk2tyosrh6LuY30mxbyvpqP
ZxRQwma3adxtyKvySiB2GYJVhWY4Pm6a13P8k0iP+2vi9vD5WJPa6Le6hxHAgV47
Au4APEhHpm/eXqIs+RoSZybvIKfMfpz558Qmcf5yF69vKtbM0Ajyugk7VLP4UiGo
mPpRAzIHuIK+kFKHMzK2kMWGoD7blM/2g/iCPXWsthfkY+CD1NyD88CMMXKX3bq3
61Wfr/O/IF0He5MpfMPqurRArB72Y1tbKp+XPB37pl5HrSX3vZh/cf4lHdtnDkaz
2Cb4zIvYfbP3FFgZe2QHSI2qNWjNyZ7/a7RpbCet4vT9vdLkJ7YNgL7rekV5JiIn
Lths6p/SyT6Z5uB836p/DB8nMDjpptYpXIUT84Bm/kEBFdDbi/Gz4Xm9o5P7tOm8
016Zh+6PtECPKfAw9dYKofA3DM8kV4fFs/Z1TRCbgt6g0gEqAqUQRSBNDbsGgent
Q6JM/MZwPJhY0c/p9kTH2JiDYAnUbPIW+2W44YOBWsCyoc00GTpYWaXageka259v
gHQQ/R3/5p9TjHASbJOw35TawLhfpfazA8pSTXA1e94HfBfW4QXFWQCCEMnVBABA
YlVdXMfUGgNRj+ztvBpaamlnh4TUQVXnrOs5hFwshhRTvDhdWmHoJ4Je5JvndGID
mRB/heqgZ4Ki22vsqUXwy6/rZo/wuhZdVnFCk6f0676nzc3PZMCFxymL2u9Lout9
a/Efq92UbH0CX3esPEajpzGxe/UdZWuK526hGFUVwj/767SdjfhFiq8gYv+MEVT+
sOilk9rUm7x+GEAbQgyM4lAtemE+4xs3/iEvRZEpomW+cTN/7MnyuRlD7+heT26v
7WblLaK1tr6xp9aJTWLTneDP9d8rlEjEh79s7zR+HSvIY2622BCb1rry6aqQgImP
hmLCJleQDRr3d0QMpubfPeD6cCcb+mJg5LRIw9bD4mifdOiic6Wis5Ulma0grSSU
jePvF0bvWk4RqDhIcqbEtUvoEpILjrXffQ3d6RkiARm1vb/vwzg1CoyvcTSovrGE
1zzsFWUPIl9RVHkKYf3ahffipOgdB85AL9/jOW2s75151HzLuqbcwNyuGO2kGLo6
tJwEzctmBAiqD0usb1c6rIZkmJhtBMeX9N7em3p0Lazaei9vXoAsJwJH41nEWb6x
Uh/XEYljFf3sZOgq29jDVZ0kb0EBhdcYZJCdbCQysst4G1hhx1hHao/6vB9bvi3z
uWIFsbtwanH5DKYHAweuD3avJoaCT5JBXumIAtf1//k0GRbxs9TaWUBdYxd9sBM4
VYDrBM7nLM0PPcM6nfCDhmimYuwVGMPPanw273J5KGhi5iLsaAPvBQtxXSauPtNN
6RVkGVEOiFZPgYg1um37aiy3cIapKGA7wu+41HqYYEHIcP8xeArQuBy5mYbMTFel
Q6LtkGbBlgtrTn3YOQUrpXWih+3OXY43szmyPUJkGcDq2zcZqaVZQq0yXoHTnqDH
rgZNpeoBpM4sNVSs4ZS23kW9cG5zeuvtQLO8l62OydssPrDSaeGG+YeXCwz+I5Fn
SBXznLH4CwLfZXTghVSnCbSuc6vDU55Sl+4vZ+qKd3+QVxGEZUqb/RavdCJa82Rb
H+XkZCzAjIUeLWbu0CKIoa+AGvsZO1RKivCl0Tf52WkxmZWpgJ6pAyrg4Pvym7Tr
tNfE7rfPRqEWNIPc3NF+FIaDlaJl2VdOKAkPNXFwdADWsE+1BX8glmMMJncZoNYF
B3TbCrAZIZKiRZOIpy7QBZGjjBw9b3bmdYRv55ookY0KLNgbPCqZygewy+1uwTmR
e4C06UFR0AOkLv56u7NWjg==
`protect END_PROTECTED
