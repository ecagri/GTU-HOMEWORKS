`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
twMDXYCRROGgUtqvo79QTPMRMjKS5v5eEqhvM7BpNXAopIbjtFHM/FhoeXQfU1sJ
7nAzDMAgXxm3qhCQt5JxCgvFzeHH3JZhxOjQlwpmCt6LvNUYnjOgnOot1oN8MyBi
LxBApdi9Co54CCj3RwRKIcQ0kQD+Bh7kA7div/PoS7tx4R5B3smeNyDAmXLoolgP
nnpm6238Iaq8o54wjdVl+2f72dw8476g/NpwcoEO68ptpkFY4qR1QH/0gvgQ6qgE
sEx57QHsK2fmw1KWcWsfpkqsP/2qk9rW0o2rZuSbR3C6c4vNi/+y7wIYlQP1X4su
k1J5kQgQXukXO0nyt7W3+Ds+MpsEKRfydkF6deIoUM5J2/IdR21ECZ5yU7UsZ+A5
bZZftwpsdNVlsqpMT3SZ7DCZRIJQVJPVXbTvUGRHMoBDcIDGEIJ44oAMBqGDNuIm
gyFvHR3kmeEw7y1JyDS+ScCVCrU/F6jr24cYKqrODT4/MXO/fXBJgkPKlG0b0Lki
pEElcJg2ZBJG4ZMSJkVCtJOczlcQcRLjT+EIedKnQ/hoJNZCBq6sxU8ta+Yku/My
hkFcOSz2/MMqDfE9pacqXyFW993Aio3mdr/koPl40dBIJ8v1c3zafkoH5S4tSGPV
9JKpq9EzaZFCwoz7yNKoiMPP0rDpQGzK6nOZKWPP4wWNNM+3+W9IKbqq459zx4O1
Dbpf6MQ+XKRo4rsWIO3DfZ+j0ISn04PVgdfewK4jfH4L835KoY08xcAQ5n6qIzly
rnEhV21tJxPx+nYs5qQ3xYwMjfNWw9lEYoRtyrVqHnKUXhlXsidQkASmrucwPExz
HPAqrGQ6HHcyaYxlMrXaPAWNYRZ08UjRE8mfraxYOXpj16Mhf9dxJxROoZSjzdx6
/gGf4W1f+Idfi21drKGWjrVciO/8xTSu8/H5corqr22nuZehpq7Zk/h/A9fNysGZ
xk6w7S8ZWMIQ1ykDl2/AeRWwn++ketDv2sRkUVcDtwmimHU9EUPr96fKtKjM7nbF
hQEkkUqANGfLZi9N5k7OCcIf0T8cFVL5a5AxC+VsgHguuN9fQxRRvS5onPIVbyII
G0vOeFggYi6/fHMK7Lsuv0LePaHq27uwcijcMWOTewCFnP9wqZSYmQIMXHFqmDjz
EKlPhWDTRJr0O+8bOWpmFuZOPxqveaCb6IFzjcrlTUXvSHvCFtnW/rt3TgRS6e/E
HF94tmIRP/I2Ffzq1UcoGNPrZzFxdL6yIE/2XNfPV89T5G3xAoJxTvIwqO3R6rsL
eJ0ayzVx8317wJUr1kJkSt/RlWIVPFX1Q+cgjSlNuTnzGYqUNxiegPnQJ6cQ9U8K
zMXHvM7JSsfdek2JOQsta4vywMBidqgyS3BhDnjKbAyFi3jTgJ4AQ6WJLKWY1uIk
HCuxUikSTkGiHDwkQ1sSu4OI8U65ISq2dAvEgFhYbfAW/mzwkV/u+hMua8Wj9NW2
uH0S/gufJqKwZsZwgq0D/Mc+zWcBv27bGXklvC3BTWq08JRSM5WSDltzuVR5Bib4
j45dU3kWXn1ClMuzi0slK1TaqaHjPTjZvho5YShP50sjJEB1iyTTH41dTF2e6yte
0z36gMrvR4e/f6CzGlWMP8fxSD4oYv3aRaaT71QId6Pia+NYve5Lkn5s3irYlQVe
5//LqlS16UY/VA62c4FpXsgrV00mJIcaAQFxs857ZAtgHhyH2GK6F8ck1bhY7qbz
aP0DO0ZrkawoeYnU3t/sGc4+NWOkBdq2LYNcTZ9vA8C3fPgYb1T4GUxBSC4mma93
eAPYd36hg9Qp/jAHmYbXbgvSMweq9Wxr3yCvQsGfI4N2v4NeX/NLL9xHbk1L4nKm
BC5ed4K69yNNukuAwhTV9fN86gvFOUDO52KsEyGAkEXASAY9k7V4K9NiEcptc+tT
VcjnYnIitKeNk6snZl7okEhsYaqsHPF2LqjsKJw7Y9czLk3JKDnImurzy7omjuMn
+9p8/p3p0MoTfdopbRxwb/CjVbQ8lRNC++sWlPzTB9i4iMoH7jrP093oxslbc9oK
/AMEH3LafooHkxtSnvJNBHqjd5s+wus5VnQkZSlB4jHF9RLJYbPP2f4AOZ6BoCaf
ENm12hJUYmC6wTO+q0SNDiBaDLC2H2YhTyLGrGxj/Iv8qoZbQO4UNNtlOwh9WnNU
4BaQ/oqzYBChBnMkiJXSZ5jj7+9sRjQXoF9Ca5O0MQ/t2J8FwuO0Du3XXS+j0/oW
yQPeYRFUTkeqRNsVQUKt3A7juMzD2cMYNxWJXUjlC9avI/sdMS6ZoSd1cNy5sZFI
eDToGLb6ukd3cBmoJnAJnY7KOPbzApkl7TvtEZdWqYHvWOcsjTlpY9JVlQL+p8si
BtQNudIMPdOGBZEcz24aaYPR2EZGvMQ5AWRRPI2VwEg/hpM6YiA1vJ90ObI7Au7U
dgO+EM4by75i9nE6ujaW2XTQE4B12ngPnmODNaZDC0fWhV86g1q14BruU4EuYoNI
o4ERNmdd2fjhbYPoCn7BikgntdQF0QT4wJwfMymlvY255iqAgTdX2js5pHpMgSrx
Fq/oHwN1DE8qfMXssUNtIOiqpENtaWwGio+ySVFPnC9TG4fxT4TqDAg1cEyuxFUc
3oyEA8UheMwqR1/YPpN78SoABBN3xB55QoLj94gdwZfF8D1cVWdQ0qgCihhu/Yuw
oO2hvkTeFXstwkLmJeA9qWbFwMNK/WDv7ORKsUbJcyGBPaOnzB6hxh8m1+AIgAEI
ArZQn8uiztaMay/xLjzb9TcgCGb2AQjhEZROwNqtYTMcnca3q+IGjMeT9HDmUd6n
Wx8I1xMHwwwF5SRbHyxiGJIbG1IPScjoVRdJgBsUcZDB/TSELs1Xtes3AGx6M/c0
yR3GDxuv6UCDzdpLBwyu2JpgVGjlFX7LOpKeaKNSeobYKG9o+HVzVXl855KnlGVK
3PrRxq9FiEEWJve4+lxzBvH4wNPjR7PJtfllUEcpBlNe4gPQIfJz6FKZ9+V9pEgY
FSuFFSeawh5A8mhuGzHqxu9rN9PlHdYNUkgznnNqgxF2ZZr01hriiy4Y82C2k+z2
05sIIfND+B2j4EHXhjpFGJkbmM4Oh0K1763RQirucP6HyYr2vAPsSSYIW9pcwGF8
Os38N6+Fzq7HO02YUI2ld1lx1CgPSa5ScBLeEkK1PGhEvhJd93g73MA23sKpWH/9
G8CRjo/4nXAIvxvNhxQBd1U3yMukGvDh17QWPhf1RQ9tNNvRFU+mpPnynSyCSNg3
FUtUA0SG1h6JK+WktUHW0InnEBRwdbG+laEqoe9elsTEpnF9PKuNNEPxwFYq2Pd4
f4gK/fUWpzTge0rLN9EaAXgaHuX2ZGe5OmKGE+NbYZs3/Akaua46mSm+5cD6U0vv
uw+n2k9am/Ur2HtpQFFfx7PI2VW8vBd0zNYZT2158Gab/sfMPmRnI3WIH4hX4u5M
TRVBQRaJY+AVrK5uQ7rgoh7TP3HyKO4kCF9524ucMd6u2SBwhYoBiz4Cxn0SLDXy
5Ciosxe5XzVql5uMAqAyqWcenDDM7c/P7pm0bfGk5RkgpR6WpzpuRwp/A9uTK5e5
Eu50GDOrNIpHHArt8EEBCRMOg33Z8K8lPAwbEgIVxN1Bjr9uMqG+SYj7P5JJ//yI
zCLmrrXG39PA+Jle8mUcg4YJ3uwpJNe0ct74wtPlZwYr9f4C5SmT4CR3zmWVObM+
YwlxEET8/ONtbjz3WtZ8b1JZv1/c/Q+3pUbNlf+ClmN6BPJzgm/iClVEHVbd3Ifk
Et/69VDJxA8vaYEtiL8GcUf+ZGtz6AzX/7rXdloeBlaoZlO3M4NG6n+M0z0sh9/R
aLXgOlZPjx9/6kHalU3exbVghMaCfl+NW/JYEktwezFciQddsO1SjPnfuzm9Hnk2
iR2+NTCNqUaWRbsZp3HqLQJZHIOTD3lzAwEysTsojYHuGx663kPJ0NJ8VPLC/Smp
t8mLdHf2EWHfugyQzxAtYC8OdwQR5AnnISYCMdv5V0gSJH/nM9GDX9awsGcxuX9R
QsfvdGgiKfpDwbKdhl7BPcMd1re6KntVvL82tQOL5GT3+i9pM7R1dudZSWqyc3CP
RX/TXSdgs6c+6125qNpWq/yj635LPB/S1QhhuLiZi6K0E3Sbsasb7NuJG6WQcP9Z
JaIAOHv/1BiSIGGJIH3AtplAkbvybWr38ucibp2kG+cOAnQDDyXAZlT56FPdt8Wv
yf6KmiGfAV1Wr8KDbswRQ8BTJi8aASwReVoa+TezFsN5Lj7lu+aVAibb495haWpG
nK31VoHzyGT1U9dTHcRESfamsCstIHkIo2+bQMzBWvUCVbRFZfcYd1hUL6yI45ey
9z+QRU2+K6SPebR6qgUsrvL6upxzC5RzDP1XaI7s7oDSK8t4Vr26K88TfoGF4+Vt
33AIHt/iZ1Rpu+tT1s6DdbzYqYfjw3lDJImNGO8+OUHTAdEIf6TJl8sB1SFL1+7C
Q8dIpa9KrfUCRsm9Bh243GBhZ7oWqaWgoKDsS9IQouWBHL5qUQktZwiSNBzAgS5Y
IexA6ZfBlP2norydzaKVtKiwWCxUqSy3/z1x2gmflmsaJPBNBqezMNtPLlmYX4yD
EgbUYRWPAuB1FpicLtIUreBDqBnTpHKBgd4ZpAJMYWIDi3iSLY1LF5EGZTJ1Q/I8
iDsuuu/tUBJPWG6eByzr+JhoUOztiyMSMDGsh6pEhAZY2O6Oj/J5mbrxNUTTR0vl
npxkIBRv4MmqtsMBLYpxMOnMY01GBSbNqcbmbXlgWMW2wxqXyIaoHf8jPlicD++R
tK7ZAdwovM0N01uJljMAEkkTR7oue25JjZe2ZLHv0VQSDZcrpqhmYuAAdeipfrda
uJUMT8wv2WDSZsR5+Gioq3gRnJ7Tipouc9gENoSn3ZNY35uL+hMxOY4k+EXbTNLM
EVb0FBwkXmII5ddJ7dhEotweTCMd+6lAkG6DadCv9IX2yTXqeUzG8L3XzMknIx2I
NjJHCqGTWKX2WxrG/U15LlD8E6aKVRGC8cQ6rp74nEPx8EdQlDGCgAoBOx0Nqv7+
/qdJLmcD3F4aQA7SHBjQc/WftwN0UkCFnxZtC57wSVgwM0X76oEkaIpLY8+eJqQV
9dN+GCE8X6N7akkjVAzxuBeuXM/6RKiFusM0Kq5Ee1XHVaYkW3LGHUx0KEEpoG8d
NTL+Z6wadZ2/0ya2Uxft82KizZWx/JJ4RNTT7kHbN/CCJ/m1YyZf7W/AGm0THC1Y
Oskl0k8inyjLQJ439agPuO0mw6DYFEhMwN4/y6JJx5hshrtTNUuobRi6e6QQ/YrD
yDc5q9Mo7jXZCEYRte/kTaM8p0jUhPz6ffTaYPSlVYbjZhllPS0PB/fbsngkBkI2
hjXInwj54nfWK+dgfN8rkt2LHoGkoA2jvq2GtIiC5lqb5BOb6IYr13C3l6M6jnKy
yEMlnySm4k0vuiajyRDWyogjiZAW7r+jKz9dNFmZTltDfGaODg+6Gca8ZnLhgI8n
yItjczfim5QsN+RVU9rqPoOtEi06y8qWdt7JrN9KRwT6IAvgZKY7sn3VWt/7Y1tm
HpsbM5htJkXkJExIxbMK2RT7m3qbUe5zv1elLJw6Ry5dJBF22qbfaSVKs7UTa4/Y
IyVFh9hQHCp3E1RJXLb7UxuUBUeqWsjOqvKABXqBUje15lsXojuST6mBhUjPsUoq
WUM/D738GfYEvox7wt3ryT0xyzWGc/eiBM4TEMoN8hEPcoOAr0+gCghoxylIrK2N
60RCDGU+QVaPFr0TIkzGv9UYnny5fd2Nu/s9Cm+8SkD6VIjGCWMCNU+4omYix+XC
aEsuKy9nW3Hr3Q+uZeUllHm+Cg6FL/hn/SUpGr9LCu2ZCzMVSQ9YYq0+u0hSlU1s
cZiC8S1q6b5619kjm9yCHWA8HLadVDlxTTEjxqNttW77Y4gBdwXaXNrQU6zDeFQ3
Jiye/6Btujmp4xdIiChglV2vlHSmCoXhm/PK4rX5QcEpSpAAM0vy6G5U3bOpYZ0t
PrMHF0SV+Ub+T14wZDQwcSMTrxdNiUTPezkHfAzrtljSO7uJYYmIi5Xr8xezHJjr
yxlVU2bap76wQRP6gqoPUu2wcZ1lRPWo5nbt8wUdvbyZDasQn8Imr/fc/e6urAPc
1ymYIMUKI4Pdc5tyjcKmwAZDk5+27udCsyns8dA5G4cxykecc4mjTWAh0dTnISBi
JsiZMnS86C4wqs9R4KcRkeq0XjFoCJZm0c4vYZZcMuVnNXpgCgsPgS4ZmdzgmOO+
3IoM0Qfl/lKQ23J3Dt2t2VZ6iy/RMryhh/7aHgKJIjIBtFoedmdQv0qM158BbpBG
yuwkv0Nh5y/FDQ5g3Acb4SFf66s8o0IWzpJzAfQu/pyiTXzk8avs397GSc41c15c
8ofW36Yp2/yP4/RSVaytxB26TGT/IUcIsMCBy6jQ7ZaOXkbaPx7hZscS+o0epgmN
hvnKV5QnCKM0AG6IouPPSiIUeuy7pBjRT4xFx3F3YFL63uxv/SNq3hXMrbRkbNGz
fZWJkDPYtW7deQu/PqcMGOORxz+is095GINRobRZzsO1OtH1jPQX9UR9aMoCksVE
7SwPU/lNapOk4KUWMcOQkH7EDPiS+gZHEO7V3/paPBUFAPlHf1008cgzXMIOpq0z
XPEXKTvBunw3xZBNwMooO+gqW34YuVjXHiZ94SMqBF0+hcbV6TAWTLz85g4tVgy1
D3EYdZYAhtmVgLXSHtHfr41VjDzzKDGGozSsGykv2cUZWiMvEqg0Ba9DwO8DlWWR
SgjrlPL3aXc+CkuRyQRpQwARbFWrGBJt0ODkH+LnW50Lq09k2Dmmk74sj38MUiaB
bs/jmJCk62gDpuLZl2Ey5Tbdx8Yl9tEQGcJ02bjGPaV9NOi3P6UXXRMUL8jgzHay
Cli+JURk2lf1/4fDCVCkdOKZcsk3R482uq9UVz/5j4vGXqo0XTVkFSkIgbM3GgQX
rTvOQpZDOIBZYdq0y3SdFSyPq+zpXjs48mgaNMUXkciYNp/bpC2a5wvgw+jJZVAx
2PzrJ7j+Q+qbCD9RPy2io5gkVHGHqdNEpyWsz7MJQdCpd5y6/u0CEED0kPNmy3wY
9L/nz6tNtYErODUO8aQVGruKJ0JQSeTiz5p+1naekrSx96I4RfawrgH1+2nLpNGX
fP7ktLSLf3wFsrZEsZXTYEK0LzQb7/idzEoaOmLPVcZ16Vx2M/Swi4XvbowBiWqS
mEqq4qs00UoeUHW1vJss+DeaY9vgSPWSykRIvL5rnMaAJD921nDBaaTWJhzOGIG5
BEOl3h6muJ9xT4DwTF3Gc82nxmJCAKED4+NfrFKsAAKkRNlLfHIxwgmJaVT4WWoc
Y8kAKGYw16gUc8mR+SK9DBpW88bVjX/Z7Ezx2FUBkDUeh0SB2Si+BdkyXXrmb5T2
qvIBkBOXCkOlAPvH4ynEAfUh001yDC3B0jLkSx1DN4x42WjGxAzA5X652I45WxSK
LX2xp7jBRCKTkmfE6yR7+b7KGDeSbZN5Pn+R7OUzxIlUxE5YH6V1+5pM2N3BW9bQ
2c4kxAsMKe5qWK8Jr/hqQUYX5bVGnvbbSi+6QB2kyfk6zvKmVtvPDRMYA8aejy3i
LXxX92ftWVFIAYHanZZygxoi+XZLryLDTCU7VepQMDbPHbKFGj6YLLouYlT98HmT
nAkp7SsSpDxdRlW6zINTboB+0kX0IodiJOWhp5zZIdnMDhF9ILyOaGXOdJnVwSRl
CEqpNpzkhaj8O1xwIs1Djye6goazwWfzyf7p8fTeZsONYCXx69lgQLRjP23r4SXU
MNYTBBJKCSvDoQ9wRK98NkJYlnZuyJQNU6t/SMELdGq6CEYyrgmmdEZ3igqfyOp4
Rkh2KGqYsZYX0wMM8Zy+pIayWdicDjmCVYqRwzI/PgG+wk7R+IaV8svKRdCE1DKW
fuua/UU76u+IJ2BAVIgd6I0GMPQpheWMzDQsClGS+F+194B1iWc7uW5d9O6B2sBq
hwsSAYg53V30U/hWDxA3SHG5MD1uRbXzNZkc8kOOmJfBLiW6KTBcpNSoGqctlISK
FdBe/AV7QZQmlJb8ZK6HzFHomELwahQo7j7oxzbANuzL4TXV12lOWtUM5Vw3jVl1
zdV/pQbZj8oGkkehm+GQVW3xiqJDLCu5JSz68yER/lcpQVj2I4sVUK/Csd/2GcXZ
5iJnbpRGzElXUV5H5FSb7AfaRf55ta6G33FOEaok4Rjjx2dGiMFylVS0f0iK6CEX
K0IQfm9FLpeYFqlPJs4AM6uof7ENAHigXLmgy5S0eCekuxazrL+rKhNzt5dBIBff
uJMrk0wStHIvZp1mEIqaYLowzeVPuvjGf1CvTUG5kmXMhoIrOUqSBsOqkyLjXORj
7XKhfZzQv+8NrtjfLm+0EGpaikRnwIfE0AdDu9etyoYqixcVXsz7/OE/HQ2ZyLvF
ZqpkIe0QIkz3bEkHlNGnPyJUhHJLreYpfwR8E/3SRPpGKe/8iek6KuxzbRmNxDvd
D/NfFKDwY8biS6mYM7QqWbqO/cWeuVEtIN2qHf0GwSZF3ryBT/33pBGjbRb3PvhK
PYXFnYvFNAmLqbQgpIAujT+ZVHgGNTFPxw7CEH3XxYtr53JAHneIbObMOEM3b5vW
RjC7iQ+1nRClEe6G2mCYgGdDra69z6U89iEdK1tcLuT+xir5LMaZaLCze8H0kokb
D3JDpXxDrF5N7vCWxVInUcc//JlPizyvvQCcJOgtvDKcWs4U4eDLOapamlDycRHM
W2S8rXqg8/wwMJqK8QzciUxmWB1ndu+E4vFyKD9Vw89HIf4AKue2N5jwrwXrv65Z
oCNR4sXkk8fvchg3qaofpqDFcj1AtB9V4UmReVB2aStcC+UuF5Q7PpwbZ7yII7g+
2mFhWmT93f+MsZuWC/JJ4QacyhAeGTPHWU4N++D4frjFZEQxcOtrH4BMStUZnHCP
yG0jMM3UbcI5DdP9oLWMQmOtUMPMrd2tKbeWxJmdoEAdFgVF48Z8yRQ+YeOa2+Ai
kEown4dv5E8/Jz+nTqmpNAujr3nI1/W/6H9yKxVBzq08LgUmTbDux+gaKeIWRGu6
sDGzwYIKHwtnfXgbpqmb6v558kHc9BA8VhuO+IZfqtf2uF2ferSgX/BnTl6tRc2+
qJwnbxlL29y/TtKqJce+W4VdajXt816/MLI3CpIUd0RDbwY5HRcRrD7ss/AXXysu
ohhY5rCvGm3KwE9SAbQUDlUCMrg8eYTOHBA/x+95bBhHuAVH37TqZbG26uRLmREU
ZpDw5MhlTT1rE6PZoyFl90n0pDHdusR4QP6VSBfGrPAmR5XVXw8/rtO0legnQjpk
HSMlP/xFvp5Ei0+PVkGVkKXRDPRAmnRiY85L+AxK1v4GLYM0aBNhFSTPiCqwz9HU
`protect END_PROTECTED
