`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CC05+CCwLTF5S0xeUWEmdTGeGGONmXRwamlt/Hj3fyiN40+AhMbxaqOp1v3Aa7BH
3VRaoNkl/697PO7VWplLBiNeLjgFzfgdf88gDqVJvh8shStFpqxTinQp+f/tMBrr
hPWc/AVTctVPuawvN2/PRtZ7taEo/tZWZSewmHpp41BSKPbPDSpkU6VpM7e7bNbT
+8dVJ4pCbOMUlpsAui5XXVC72h/culylVsTpmUJvlk3DdorQxf3UJ+NLou3hOo/P
Yz6rV8nqf8uTgQ0W3B3RMTJrgSWgkFuacotd1dj0AQlbmpFBSGSRuWmHOYkEDTah
W8on+DFSnaQHot0uoqBkocxsF4b3e+lBoTHfltV/dNFrbo7daDTst0XtcwLGf1jh
Czla82vn4GWPv2pipVYN331WmiqAOiljTrQF2FtrVSPRc30pS7wimkODaJlaJkFD
cUh4fCz64sKB2wEKfDuovzlrYvxp6TmYtu694djVJ9R60te+cUy21XJRPYMSbFCq
MppUWdgeM1QAE1Z6MmTwRYUK9WOGngqwjoLAtiuvZvlBc5QOC2c0OBrJ4hRGour3
yNS9aWWFliao0Jn1BK53tyUXkZUVA+u2cKEfD6Uj6L7dv95g/0G38zI/1bAVqCs5
BaeGDoemeli1XDVjjS0hLuh3VtZQWucAR7QibjcEamqrSHHV1gvWX/TjZFJuH2AT
cKQqHnwn8x1pKx/FNBrMWmiJXa4x505SmRfOEPu0yvQYdi907LoajUzyn4lvZaCl
oKWNSjBch0iGRZhL0CV6vaqUOCXYStpBamddZp7nXg40cz0VKZ3j/bVgV6sj/cOd
sb+hVzBova9CHVs0OP0GkB/FfFhoNFUk4nuIdGvlI63norfMKsAIr4phx2S1uFVZ
Tf5Q4haFhviuxq147tWCAihk83tZgD5zSCQgu3l8QKG6o5zZkmm9wAmmc+SiDrlg
wkqwQhsluqxQaNyQA3J1wVMtn9f+dviTA20I7OF3jfZ/98tkz633/5h4OUMTAB4Z
BQpKkvBcD9mx4W6jXrhjKndM2ATzLoR5L46aakAngpONvd9G3McLSzrhUU9fcYYD
0ah622yxt0C7IVEgVvK+FgDmSoeeJ7UhcBqfHC+DYfJjJDvp622Ihpsf6tCU2Z3I
ZnNtTOOv2KoFS1ZoG3fsC8YoSIPJpSd1JkfkNI5baq6q1+nT7NtH6/blL6tCCHPq
+vO4XgrXuGICBCcotaaR2DY3Al5+NFuZuihwEjz3X9nm2gt8epPFCTfn5rWa1YNA
Cj4vrWrVkT6nvDX/ni70dTJlaSNvlJilDU1kzX9ospCG2TXplCeOTqnNJ7nAP4+s
nzt08klr43ey6peS6YfVXSH46f53i7rRgBIDEyReQjqzoBKLrNS5+W8eRiUmkMYf
Cqba92AzppPOF08X5LFaZEC/trBAX5HUIT5yo5POAHB2FbSoW8hsZUh/Awk5/YoY
o4v40EIgNSZo6PPvFA7fwh45F9Ck1/rvVt8WHc+Ygz66PswDLkwe1yVv2qTBvFvM
dNkEtsZtS1Paf7I1Fgo5DZhvwLH7hlqPMyJQTPDXAtQbc2kMz/BXPvSgH1huL7iB
+2vpvxk+JExZPiz6BvsuXjqeaGKhCT8vxpj8j4yq1OUkhIrkfBIAl6OPdv/3hG2W
1PCkvykuI9tuG/Bgz+BhJHB3IQd7GqpzFO+Iia1A/23pZqVShiVdjr3bhosOwnl7
wpRrOwrbJPljZTQskW2djiw2/UCrufjrcBbVhKWwhVMN3U6H4mt3qlCPsEgNFo8q
2sE3EmjXLX8zjreHHxn8ddc6AbshhqhFtiSqIQnVoPD10KTrgeQWhblATlqmRjuF
o4J+1Uy93m5JnFIWTImg1+bsBmTr1nsUi7c+6qxg2lVn4QAr9ip8aepNrgYjr9lF
I2NF3SfEQlZWjFp08sXBpZk0U+3tOPAV7/kRVK9ckILY1rh/A3kXER5dbsYZd0JV
Hp7gyEtYMmBXJBfxI9blgCfW0MRY1aSk4lmvN72sWLezD2Q0ILTFtQs7WFw2WTFk
GNQlgdNqQxYrHxRrajbWxjtedcl8TNrdJKs7MG+B9k7sh3iratxVeAa33vjQCDkh
KIUKdgquZQg8OtZ7Rcl33RpA2tIy7CWTIA4ymgnTGK6twNWLZ7TCu2LYA49MfgOH
CAimgToYpbNONWcQLBGPun13DyU+FQC1oJ1QgeHJnQSuyx0d504vft6LcMKl3EWb
Z+mGICI65nMrpArQzGVww2oChDE3EwcWhSvZWto+9B0Kke4xBy/hb9vCMgCeqQ92
4t71JDFtyo6tyz0fp0TtW388I6jbPei7PdrBYcBcJQpKgDipsueA6846Xxntu0tL
xy2wwg0G0UkbJ6xYU1tnFKKn1kCzSZbv2/6wghD391oUS82HjBh1R4qv3+hsFBKd
n/jV7KpCE4NOAJYJfGifbPM3bF9etMwSqHvGSb813TfhlxMSxM/7Uq+C64ID79XN
B3+6UlwPvhh7S6C5HECAZr03e/mWDD8nAoB1NeGNi9IZnZXCWac8epQp81USAxgY
OvS8aoV1eNC3pRBa38UIpg6GUbB8SV8ANXqkpqfYfG9eh99bdr9RWnUIGfpAcOQr
tD8sbo8yevo1W8KbPZnwUnE9xOlqmsWBzI1pKWdM+fAStPSc5NeedObEefSN0Cfe
vBUgpNHiwPeqgPJ+8JrLAx8mhaPpDQay+Ks+ke/hk8hEDSie4Q+t5YiaoW2x11ja
jT2E5PQGvgf/ih5X6dIK8meWhR8oIy5j/Mu6WdKyH24iHHbD1r97Cjf1hnfRpuzw
4H+hKYiybL0xhJb0GAIFkYopbVk+faSdC6ExFjfFrRdtvo6435yTWa+1vhQLVdXt
54YUZw63qOWK248O0GjQWpkgH7KqigK5dHYClZGnduz3CcFcsIjafG17xpezD/8r
ECEJlIK+yW/kO+mBFTXzL+0zb74wTj/ZYoyGe5Cy6vzhTIHwtppHCeyr+VQphURK
YdJsTd0xRjWl3RlfKUw3TGf7nmoz+bvAzjiUxa8Y3kJ8OCYCQ55ZivOg9vvnZHK7
wM4x4UQ+tU7+Ife/LOzyQ8bDZa3+wUtqNKoyH4/n+LsZEpassgcdRstXaRpB2Qta
u2ny1PFpn6cBLbP8T1+qhEUVrYDnetoI3aiOcnBFNoVaEOExGwPHt5KbYKKHBhDr
Ca/xpa5CH848DBdcrQ7Pwxfvjrl2d8Mtzug8pOY89ABHuWMVR11REKaLZRqCJUNz
R3R1ig4haWXwIsduLEpc+2dNKXH5KT4MCNSNPMc1WwO7rdkcIJmKGyX6AGpy254t
SyHfLW3Cj2G3bsnlGx1nyXZOqNws75WwtvKoJHR+T/0qKuS5AtgbP2jfufPcc7NC
eSXZ1He5jvYgHf2uB9gsaF4Dh+RVrLcbKerqVauiImmPsZVQyhLZd5CXpKw7WZ3k
0SBLt804Go7s/h98pW+HvCbS0C/bkjjNQ4tYlLqU9mCBoEGo4Pt2G6a9y6+WtVF3
tLigfJ7hRjoR1gxQMm5R4qCTMYWWRJ5D+UwKoHFl6QVjVrWDSbK6l1va9lXHloEg
cCU2/50jdvpwGAgyz5zHhOG7MTpr/VzIQoXtM9FW3qOlu9KU5n5kClc8Pi63S11B
wy6uT2YaWZ0a9Bui37P85i06mekt1R8ACYAYngWiG7ftR9l4IzEDTwoHIal8sBW/
IianvuHZTqIFekgDoEZIJz25YFSrWBf+6XoD0cpTbSi/D899ONgsHSgYcC4PJlV1
zkm808mb3V17/duTi49OneuSkhS0METfEWp9/QYslzqqdgnjdMJuA/gm6TVYE6Cf
S1ohBgIxPh/+u2Eoy8AvkHNPWar+QZUrsmdfDxsfIXhG4Rg//D7ogdl+ldJWjvlH
ricloCN3v6dHMwAMf0ZyYWUi8vjChlddrzLjkGzmMTS0f+LekML7bmHbCsrZGkGW
34w3mSiLXzERi7Ujt7HrxTVDGsB0ylEPpu3pxi97ujp28QdPb4wU0i4oTK3iOQZf
oOr5qU8aYRItAgxEDLjNVp9i+iUk5YfFYSHPFiUT93E7NzhdlU6BxxXjIx3WGTHJ
rYRW8wODsPHI2F0mF1cs3+/inDwZKHVuz4KTx/q8VnUkv4vkwl75ShcF0mLrUXw5
DV8e/4FulQ+bM3nq2vU3ZbURSn8pgNzFbNKmnMJYPT5zDoFaD6XJQkTmUmshLsxO
bs6+/JxGsm1b65mPNXj2ykrEEXlniKIQ7yAAx7kws0rXTeks2/L4auP+sT8+RFUy
HgNE5pt17RddznzVz2o4M5BA5x3J9cv8DpMKnby49YLO1DyUfimgj0gWRGItWQ+T
Cv78KNZeA/rUdDOURvPjDdR3AmIUvnzjnCrlSOrFi+YfAGA+lI7dlLCpXD1XwvNy
hPo7w1wSuha/JJU8yhr+w2zlW66VUwRiqHvLhEUOgsIoCNPKFZHOp20B0KaJJfnM
TLPpxarbpAusqaoAERyZTVCEV8Y2wZwgQnMYq8W9OQHlocxgCQ9GZeHcR82mcIHS
Ui8OUgwyCBYvEDuAZWPdWHnGeY9HjVIhAJYgqv3ER0TS38OOLjn4AREUNJE/F1vT
YkkUvBBVu4QfdNCL9Uk5O9kQGyesBrMa5V2MZHJAtOYK7pKxVXXptsqacVqsqR//
REImQ6W12qEwwSqc+v53BO7szBHL6QASCRYVO5EXzi3pcYbZnpKjDPhanFn68Fvc
3+fsUZWW8+VAieuiLNBRtSMXs/c/cWnQQ1ruCkdeqSk3Dc111g/EDjPER+PbH+mg
5XhxvzYWjwSWszR6ilsWI2ncySrCn+5JqT4fyKUYt2VlGrw2ibz13Cv8C2+z4huz
GakzaHrmJQ9lMipJ0kj1Y3pcHp+swjVv7aEoWVXrxnlG4jAC0RnnTTkEaqPyDGyL
N6JVPFRx6ARA1+0Ne3JI5SxjuIqLQSNrxrVZEf11wIsrK9xYM4IFCaU9T9Nd6qrm
Qa7tUE92ak/5jFq4EX3FUOdKhoWndgkXPx/3eV9dbR9zRI5hg7f6Ny8tA3h97Qa4
JpSFHg3nvBFptNl7wX9/80VFEewZxJLcN/cL5gQwiHYq8geEwWRcN9LWUyOYtZe3
J9v0QQnmn0PBIJADOpCjDSnGHOksHtK0HYmIi3oySqsq2qYSX1XerpbcPJu9wCpA
rHBwjry+Bazk+nDwQQZ1tWUeSgsovr0AbjDEycNQVkwuJl2CPFJWdtsoqjR8sP2F
kCxHZP00QaCZhTCxcYKn0f7ibXt7smGqpboa/c/Fw39NYz5xCXw/NPRr6r6/kfEw
9TcdTvKlfEdLuWc2PHhS1N24D4V0zaG2oQD2JhG/BP2Ca3vGq61jiT9oor+tSjsS
RxnOs4GvoGVMBpG8VCrYqd48TqLzmq/TELpQgG8b0b6VAn0v6KVPSn52NWAouL+3
mHDUzyInlmvt9kolxdaWFweaELL6qK2+HI1T9AYYF91hJ57HfF7uIWqUpjds2tdM
LVclIIb0DWbbaxSFUChnEXAc+y6eyccoovgYsZgqjlyXUWaXSqr2tJyH3GdzlLcg
NvXUgeyyz2tSWOH6xzDg+ocG4dg2dkoGUtHMvYtqqMum2GvgHsHcItv9PNkd2q0Q
o9ZF5Yw1eaNA6ZnESo1pR1nJwjt11yIyv5wmE69YwY1EQaIX2cOLTOUuC+iqRUFH
+kePAeJ+oRO6PZFCNv/qGl4P6d3tdpcQIHmSdNanunC4ToCZ9REaf6hvTkmQgtwD
IiEpKAQ6+Fl7xGvmT8BoQwi2xqkZXTEpDAKolEkYv88MUH8DxoPrX1t1SSu0crIf
4BA9LEQFAHM7nF7dVCcSande4P0wtoIK2cRjDrAFyD8NlAK5XK2g2W4uSQMSgifl
fHln+LQKKzcZDz2AT0xasQV9Asez2I7rUVW2SJFOL2sb3xaFPDUYdRwnjXVRdIzQ
yoY87bpG1KjW4KzMxFzjEvX5y4WkuNzubiMOkBF51JKXbc7NGffJrfaOr4kR3BLm
JoTfmophx8qy00YtwA2VNEYXOrxwphGfxQ+nJAQkmvOIvKGMd4GELFZjC2tNiRKI
IGRs5rLVWboO495bLg5U985lbH/Ztv7odk+9N4Us634x4iVBK3Kte4FGAY8dTSmx
IB3BGsSIn/8geqVif1ao6w9cuXLmRZ07ipQ0htmqHT3RA4+39Y/7aAf4eedE8/qx
PYEPR4sA3jWCPG487tX15Bu8cUMTlM6+rkQ0y2zSFGHaJ54GURLnfVzXPjBYPngO
QWXCzR6j1+UQ/qKpilftcbYNM338XHbH7Om+7QWcm37zul79Plr/Jd34Dd1AtuBv
V5ZaIAhELO1fQu2HfaDHh62RMZZ818QWi91NtoeFoi1rRuuyai+Nq4KG91762nCn
5Xfzm7+auFhcikBXM67ZZ6N6cWEcMiYEjNlnzjQbDjVzksWxS8wNULeQNNvYP8Yn
8OKTHE0U5UnVUC142W/Pepi95YV+QsM6scllOZPFbW3ZOErtr75YXR9rPQNSJYw0
bKlib+TRKUDH2lynLItS79d2b1cZdygHhhHdpW9RnRlx/InlcwLkyqC82XmyIaRx
f0la0gmMaKG/JjF9m51kKC8njJ9djRiC3P3QxKFzRImHbjPT3T6JC+cr2u4OGTNH
UEtc42HrKKfe9q5FjeLAhLKj6mtE/AnvjMf6sMmXyudhw8dnl5BcAdLTFlk8bOAk
VQqCpIddKLFBP4lAhIj85DMy8N6SEz2CDH5M90nTUEYcv3NQkA8g2oIRudPD7TWo
8OVysxAOSGqeS6CEExhkYn0VApyl0X9+sCwxCWh2y+XvaJNaitj4X0dmRzzfvwsH
KIu+U8Pf3wJl8IwbPrex6Y6dw5fWSQPbEJXnoNgy8X0iWUgbW0t0p2hBDy+PN9ak
5XR3n2sWyVkkx60B5fwRrAEFaX/hEYgDeOQ5Gqp6+nOirnCFdmvbMNCx9m0OvpG6
5UiUkNTkWjVEjUazrmz0Jcmnykv2C7jc1s48gakGsbHCrb3Tkg5sKo214eXr7j+8
kPLoXTt3dA7GWhWcsFbzyVMxBQFoD5UdHN9/288khI4Plx7LADcjS7w4aJBgb8pq
9V1MyA4qRdub8lkDcZ7ldFDPz+5eRNC5eJerrYB0Eejadert8mKB+ilog/ToL0+i
A8Uh6eqIKkLryXE87hicY1BIgdgpnpHa1NG97sn/LPkhXrsZ5d9ZbYrEfzfr0X0O
p8TeCmOys2Co54UR4IAskOSIypWa/SIUWxN1zuohk7jCq4nduipQnik20zGD2EjJ
7FAkb4jIq0FwBw+GEh7YCU+uZmNYitBmTAYaNXJrcffc8r20P9y+wVy/Lce+RBXx
fndr4txxX8GKCGRwZ6rYfjtZYm/SfEvfY+XcqsCVQRZ9CNr77Ezg85mKVlEv0XAE
FZ/dM2aN1x450gEF8giWTIdoIHBfmMAW7gizOtjcAH1HPi5PjVrt759U3gCIH9oT
j3QBOjHOYME4aF639FCm6LXcew46VpnMwkml3c+PUu3JJ/x9Nvn7QGiBSrdnZgeC
p3y/IxZucxvzfVOkSPqBgXuEMC4Mo9MUoNR88XoEiePRilAqo/32MeeXLDkSNjYD
4SC3ZARUxWbD44BLYEgsf0ctVOnDbb5AsurLHK1W5mEya5JKjF/Jh9h78R7NSgKv
VCLGIBGfHgrOJDLxuMF1UWEWGlR8ks63RFgEmqVVUQh8bJbKNf5xdKASQ4mMvr/G
J3SBCuB1ox9PNEpGE5AplU5xHs2xalQQfhOjbR0PMrM1UO7dEeeNU5uITMQbqwgy
ctk1BO+5BtXKJkjwUd6blkbTdr3dweZYzP8yfcIswPbuWdSND422Wbj+DWrZpd28
N3pYCdmohmisoabnXcm3oUgfUOXcb0rav2oMYbHv2vN6s9D4jbzodfdKAhV+DHkW
IsgQXUqU3arlxyCR3Sfvy6osJSF+yeAShfZ7lRQL0lBOvaek8LSXUlbBjDtQgiFO
roMGw2/sCmRvbHRRJ17st5YWi5Bl2l9IkofqcqMEAlSseTqxJZFPX+tzKIqjqaSU
W7jJiHfzMn6OJWUMcVcph2O2BSfCr9Es3sDTqnusLwtSY59wuPK961gl2g+MsSLH
UNP+93KaW9fiLrXtvpP/+6ISf8juhBf3R156ntlK5mCDe/YSh1xhyXF5VKqIvVY8
ixaE4WKfNkcEV+hAYTki29FVJiXuPQ7Pg7r1uvRE+V16bZ/RbuivojEpZ7ZAaNLc
4TjFf7teQhT3i2cVjhUTqB3aoA4Itc0LmBUlyDYfo95MgWX9jmoqzAzu2YDE1fYO
x/6XtbdBj3BDOnDbq739gRJAO4LI0OtjDPRg9tPu6lquwj21cu3joOpzpE4qf3Po
OQmfwoVgfh8Q5JgGIfZiuzkfREBhdp2oefr24TCQXmHp/tQd0993dTPoOsdnhdHP
qagQeFvtYzC8qEobcKL+OWs1Hiu/X+ZgPnFO07Bi7FBO1OHppduyXACBBvK/R0X3
AbQfjvYwtIzAwNdig7J4Ugq3rjhqMfQAeUs9GELZwfZaOxbb9ucS3rvQoE8fMNKQ
nQrrxEvLjJJO8sXyoHvkX8CbMxONzIaTZiuaMK/fbdBCS+6doY3AY6C6rWKJTcY6
nTv1XvggjKVv4PYFV6KxbPZvt/rwnd6CLH5oln8gfZ/OHkQfHjsgZREhMZF9xAde
Qzy8yuY/w26lmQP5kcPSzofKJuCR0EXlIGG6ubRkq8r5s8qvIPZE1OCM3mq7ON7u
3+2OOhDM/uF5MT6rhaKPemF+3ZkHY+AVrfjeJlzJzMQxj7juqdk657eINO+IM+pb
dIfUrvjpbExBrG/HQvWGe/YU/nHXRHXwt1vz+ev6xmDIHCV2uOKOZFDYOkoAOFW4
jA1Cm3JBX/UWMWjMfYORtaYxzqbQuCTxfnDcD+VZfq0r0T+jzAdf6y4cGst1xQ+8
AMIfQzZTDjuIB/AbsiIRaKmugFmA1VRU4hxKVOd7e12r+XtV/MrjcncHVMGqxfjL
yfVUkBdH0ZDpVIoVydQVa3qnQpp29yz3gQR8xFyemO6++gAzHJMNDzLSt/PkvZFg
31AM5PD65qfTcS/Cs+EEDZXFZmaH8Bl/rekbItIaDdvHXfLQEa823pCj9yngXgpK
xkx7EPD7fOWGcpaJxDMbfltQIJRYxruAk24hRzgZY8iOM8e85qBmRWP65ZvRcKtq
xDNuxZebZbIUnxjXMdkKB0euSCTG5Snr/9hVKrYFjq7fLqngxE+PSvEgMSfXBFcA
NPzapdoUG73Ag9zWFdgrxMZJKTtjDBdA9KMFEpWWG3NHZwHMTSksqh2+YHlv/kbD
OZtimCliDaOJzvQW7Ewv2W5WIUUnTuJcX6YrmpsCjFeeF9ikBL7pFXpahyV88L+Z
Rh3Al36ScJhZF8QmR8+BBXkkuZDZ+B8V3z/ffauLnHlt7iF8lzd+ZjZvwMnnlkix
tH1C+PqmSB1aw3NxLao4w0IMVck2vdgOwX15HhKTrvZt3uVZDcsrdzWV7LrM5BsT
USPNEs22nr+OLK4nmGdoxD/n0WIdZlIH2fq6JSc0dEd44J64G3J21MBHL6E3ufNc
xQesXdx9hLnBcVzpSFc4DMxs+XWq81K0UoZxsRncKdTmMVytfYQcrFDlB5J4Y0RS
UHA64gEEPSk4r5bvzR0WLBJm9plU62lqmcZS5LQYAoOnvgsVfRmqxV6HAGxgwjuD
WCtQDm4tqSDktOBPFNvRbx8aosEgKp5mX6f0uiRMMXpI2dnv6/NX/B9GJFaqY+q4
ieCrG7oMqPmPoncxuC/OFCM0Sx8l6AWaL9ma21TuuLbkq2UCgRTjHXa6WA81s4SD
9otwIesG1EXLc19ngsUvQ3HVWH9x5/K+Y+Tm5W4Ww+xa36qa3cVZBXdga+6PDI1B
qti0thXSVC5iZfrGk6GG1B1HtGhTnYs5TcyzKn5D/IjHlgUrSSGLDQOAECHMRccX
rloS7D1ZtZ+u6XAoDiuS6s+hOWkruKsSuxvywoKKBnBjPmAtt8PTm42OpMWSO2vw
g15acmRbxA9ppmsoVLjqg3vUixbYng1gyDBlDMLWUljaX1gDruymy6mF++SQzKpc
jTIIhYcfXwqhY6tE/kRJmSic11GqD4lDyjg9dWxoEAOvghVEg/Hyb4oF0X17l2kL
2oB8MKo+N+RSeJiVwJ6rAuhq/6U34b3GnvrPbj3csZvwfxdETCxqsSKeiwPM2S6t
Wvta/w1KPVOCQmJNPM7OeCaJWbFZVEYTii77/WBQd6LJG7WRtlKE7upig7TLh4mA
2hznlPZ3D2NtIIs93FbIpEI+KdlL8NpMlkEUYTzA+4qW0Vfm+R/IZXQ9jhHBN+9D
GXLqDVLEVUM0uGxRuPMjV1xGJSkSgHuVvmHV1ouAVhBawqx5NJ0zIh3YkAatjvyc
SwjvL0+5kqRzmB5RBVzBMZAXpQ3YppCDH8tRzAH+1HvXW2FgAdBbEjUhGKXUB58W
06LutK10tH0u+5Dx0EWyV2YpDDfVf2prGe87OasrQkXrR0W3wAZncUUuUhKB7AOB
vir+tQVnNpOku8XY6DLciLb49YOgG69BcGqGpNieb8TWO8y+KnCGRv0nMzVKepjK
oOWYUg9y2ESUonRpIEza5Lu3A1hv6KlCknwJkiUdsKSPAln1bAPhYtfg4O5IIYjt
HcrfZsVrgneAXjl7gPb+8ehqnOUsWlaO+FpTwzlViTgcyNMz31JRQSjM1kAiaaX6
EWSxFyekfZ+T71vkvpk37sB8LhfanxiffchzCIU9Tpw1kmtTmvMB6miyoqm8SVTR
q+no49n0fdPu25IMqeQZBXMBEHjpTCQ6/rCdreKn+VkWVsM5Mkg3I4M4sragmuT8
ofxHQJPNs3iRXDFTlMI7TAggy0Yns+yYCZKSiIsjB3Cf2HeE5OdJfyKKLbiCQu0q
GRWL5U0ZY3949ZsgXrJwcGUNrdBChmpHx3CPNOVtfwZny2cMUGBwaIzvlxIBwQaD
q2tONMkoJbVH7sGvw9e4PIDEx+l+BVY4EuU7vUP2wkDX4NqQB4I6U1Z4nOtAIAPY
DunsxMEfB0pMh7IT6CG8wiv/uNjJMPG9/hknwetEoXIdYXDowixQ51qNK4RQ2z9t
vV9nkXbR+kdQj+XkFrK6SGqU09N6osftralbNHm2HGEAAPUEcg1RRPjpPW3itexM
RX71wjjdEOeMjak+de/W/M+R72JRp3te44r5jtVuJhNxcSUlUY4n54MUzspoU9Ej
TRFTM4H4fwi53ljxiYbc5Ay5/HWOWrHZ3SrxyO1SAKNcfCEAHQR4JelFK1XLUccD
vPFPKPuqwwc8QBnn3m1mnFgW6bb/DCtNiWFvNiVf1Ii5ARBPTHmzMCBR39S9EX8r
6gFcX14oSrDSnW4isD1G4tscT1+tCPdfX1vDEsehcKI16hWyB50xYfl0Gzo48/ML
UujpQsT9hT2sVLWiDMfHgVygcZscJvilHP1oKEEhd071zeHe1g4VZBMS73j00fhW
1Xwu3DO8bVjhCq4jtrggC41dRKz98Qy1CjYEpFitpynClvkBlOhGsJRKjDPY2mVR
+PLb2eVawiw8+K4PEXEuEnSlkKIxgQyCzvfAUFUEayUTGJIx7fbrZw8e9DAAaI23
oLiACaY/H1XDZzl6U5tlShSOKV6miiMGTlZxMGlOmKpq+j/9b9Pg3pBpCj0gGWDu
Gmu54lUsXfxUE9oLnyQNC/LUHWjvHXnOOPbZSf+VMcoIyxi6shYM+yidzbCAupis
OZkmbELYKD+TWbNP5bk60DYK26wUQPppomhzXJ640Uo6EmVvLUIqQfRjpcBR4hJB
ITRrFnzICw319sbLJQQbUhfpV3h5qN/jNl6cc1jSwR/oRLNtDivxGwtqk13S0fD5
GMC7peklkMdCiCyqPKF1TY9TrJ7EIj3yQU62J0/e92CeVSz3sm1mR/L7Gnr8WJEt
lJlA6kDza3fxQxr8366LkFT/Z+wZJ2KUrMr/z2NRo9EtJrVRLWjums+IixiR1k0x
f0dLpobO2eysxY8RFcdmipLowdO65k4R5dHv1vcsZIzkQ0IVygnsaDtexFst6wWy
8YBFsVMAuH49rqMg3ELDYPpueNsHJYcQwVvSrf77TWaXwWyegFa4UD1M+MkZ0uhD
H00zi7jF2lLGlW7+Ilc54jFdULuxQNmUg1TVGpvxdV2r7XT6i27zXxQq4imqJB2i
m4V+3IcT0H+wd+tlJAo8sLoY8v9biTxbGwdDtbVhbm0g0NQnQevk/1eHvVn3OHTM
B6rkx9RgOaZwvvIyWocBB5msTinm4fT3bO3+ZOZaTG3PKaWw0qMm6OInQkKaEfKA
o5U+SyQdq66BYupQ+5x1FAR6q0WvMA1BYjeLhXf6BtePmwQ1mByXWo6FJGHEHd+1
5hQ6LvuuasJLaimpnRi4unO6f+nqzJ99ZnhEbQTN7HqAAGkxCzghtOfZ3dM0rC7Q
iNwiu5F410H5+c7zDUol4SKjZHG7jMtVRWoZF2L0O23N2djkfsZAnE3G71wVMT5G
7QXET4BuP+YExduCJO6DIawdMnQ1MPwwdReK5zsBH12xpEZlUs1Bo7iYhooW7tG6
JAc1ZhBqOyZMnFaI2P30l02ed4g9+g+R2UAR7DroyYYNp7QMQstQPjpcj5ewG1k1
AckR9SZbdCI7RfgJxO2U5CdmHghvXlUmavbedJ+v9bFKM1g7vQh4rq1P0hmT+tht
WokmRO59z/G0EtQfg0EF++mWgZcZ1Fmx1+seFOOJVy7LJZnHSlLYGwh+CXcY+F5T
HmkBvSKdlxOt2dQNMUzAzMJBFDcdzODPLRNk4OKUZZ0cX5c518mNwbOfGXNZp87t
9bnMHlDl69HbljQZOburVi9jzpxNSgLwdQQnuC+3q0eCdw4S4w+sVh+KQjAMRvqs
Tzu/0niEcyyQ0OkEusvgQH8LFTR69Xr5paj8ptyzR8tA1zCDNgujdSPJth90zZtf
Ayt/LKPCVlJ++B6hG0J2VwA9+Mn9qCGpDgo7CimTMI3e3R4XsLeCQ+kDz3QNjeJu
/VlqN7CJtUvLYHq7m12n9ZL5lUWY65GmdyuaxXWCUj11aBrmuKeBHy+uDEFP8izf
/yXn3DCSsCxbIZHIUAzmOQ+eJtkuhJeotWQh889yCsJDiUJsYpCPhy0rPvjLWu7o
Eb3nHGfmhO4ioqIIERnb2725Q4tnWb4aeJiS5RGheqW+EKwH4uzAmRyOiP0YjQUl
rFqvgjexkO33Zx4z7SxwiYlRdUml8vkcbljaoZ9IAyuzuvRKE/mT/4HsxkJ3tmtV
4dWYWegwkoiyT6vKtWEpQBoPemTFt3kaT4wfoH/h2sqiJGZcs8E+t2j25e0CpkTk
DRgKSb7Dvl/u2i4XD+oYBDARMEbvtFoteX9cnh6rX2Cv/bprRYgdl4vAH3AAOAF+
kF3rPrMYSE9+4dsc7ta87LVpbIpqG2D9XyeWU8wmB2RImbHbfoGyAMLE7AIZi/9j
DcwrocZ/IzJA1Veq46Z/IqkZ8eqHE7yoI1m4veE5RPVhXbC5idBhLc1v1ynUuF2n
yVxut20gaeGA1GhKWtCoVuUUYolL8h/5NcK8gjcoHqOeONeH+KSAt9frRzgYyBUL
jjfGwsWdogmB8zRbP74zFewswxT1n3PaL2qPAfeCnhz0qrcQQbhPDXEw4alOlMCK
7eofx9TjwPoqpZDpnqogceNM5j9K1kYVW29z1HrlH+PSJ9G2nF0WHf0l24lTxexW
iXna8mU/fnssMknG5b2QTa6kRLiW7b/QM7KGwxnW1YLZgWZcQnjHfoHzQH7H+eUf
dOJEkegiasPNYewXNn320ivNrykhhq5qbR+NKxxog4TgR9uOivXHobd/XkAsUzaK
R5+0JXghCcrW7sMxvDJSB+5gl9zto3Ip5nPF/LVkxAcRa329wd2Xq4xj+BzA24FD
P1OxEouj7+xNEQI9Chm+XxFFFalVPZKgcsYTaS4vXObKoPTsT5YEe/ZyM4c+6IIv
m5itUf1fmYN+3dX48L7Fz0UlPF46iOsQA+0fLZkq+g7PkEpU0XqgwBs48Z0ROl64
zFDaiP2THaWlNOXAvxCzluqTOhADFTGVhBGTO5brOiXfXUKpFCQgvEHBI24FqQOF
+kZeU4+Bd/lbttrcDE3eoAEtGmp390nj0BlhzBOjaPCWmwwFYluG9MRTNWZ6JmAh
bvx4DT3kWXW7mrE0/HAIDl/ERRVUHXq9f1BJzT1ymy+p+nTs0li+JnSAVs68inm6
6DMWn290FOvNK5ZmGGl6N75vR2SRGRpbYpFF64RZF+cjmlbcqeje3JriFgXhlexn
J/uyukaCRL8pYkYwp9QtK5mh/jDh6HXZlhc1jE9dXEjn+s3DC9npegAYAWSlO6Ru
Nq9Ra3CmDyCJ5AEJa2npRYOrZyalBuv79DURq8+/KhEN+2DzPYpwawkHQlgdo+SG
dd4tXztnvm8GRbbeW7i5yiT2dWk8lz3/TUQYZEiwICy6RwdHwWkS4Z1WLTvwb7N6
V3mD/phx7dayUuz35BrU1FM2Nux2sRLv8mwetgpTD8oQaMLNSZSdq3SLoI15TJak
bWasRlWsPVWVG/xxB3SYng8+aIJjrThSJcut8lYCwFd833SxgrwuMXn3Ivrz3Dud
QMjcDUxN7KBu/S+G3d4oINAAqbGs9UcvAjzPx2f5MKoaxEDOkz7/5iunKuTuoI9Y
Pd2aSeLw7eV8ONGtI51/LpSpiu0UBAml/JffmdxP2BOHA34I+QjZqW4ZA49RH2An
1wC9KfQnSbNQHg4f5YEWzqwam4a9bKkbWj4iOHr3Pd3qPjwcKh34BR4Li1MnTYY4
o6ccKJsnvoVVhuJu/XN9kXQSo4xV11/Isi0CMokmHbFS7Pgwt/SOxPm42vbd811z
DQq0hcesL8C5g4JCexuK6cEfNnxsRoEQvpkAFKjZVr8Lkl58hjdqEhbLuq/I3TWh
mq/M+GPM4yMUu0Lef4+TKsHtHtp3owtIjJM7SQyhOlo5Z8Qya78ngIEEuvpg7My1
k4sVbZVUnD133XdpDOwR5rSzcLAzgK8zhAWNXSSS2kVkLYxbG1dQ6fbKBIOVCKgN
95lGaFjnjTiEAVYKmUXR0G+CtL7EgWckCJKqckkIyvUX6PiTxbtc5VUa5xB2rUvz
RUqKuedKf3KlCODpuzxL1vdNIeDmPMtBu5IxL0xKzO1aQX59JOPBtNS65FALd+NL
T3F0KVvLoOLUdUSQhuuM0Howe2XaDEqkp2vkZkCKN0nZZDhWwjFiCYIwBUuCs7+8
x98huC8upeqqPVo0zYVlevs2Z1VI/LMrj+AorUnsfoLUy6DcceilUI2lk/5VW4zZ
CQiJCMbJwGpZQrcEdnESOmopsU5buI8WZzfiuTwEFEsvBazsG+Fx7j6h7LUAT2eN
bndFR8+lPuJbiLbwryisf5hHeJkpccibr2YVOKVVNAvDnGRs+jT/mH3Hp4bFC1+2
pqFAWGTGD/ofESblNBMPgpYvMvACoe8zQ0NBaeNOicb/pnrTITdLgFuf0FgdKM1y
ocvpwyMiw5lpTwnJleZ45p7EY2ywBcLqgIG7VK+vdUl9QKXhmo2fWyJ1c5COTleX
iqe1OvL/qL/krgi7Q+hP/aYM4FGRZ+xgFZy/Psd/tr7AFhGbTJ5S4eK5goUPYBIK
KDZzWXGG23EKDCfdDwjIbRYJr8026LHNPVf6BnNkOYSeSnWZbYSwa+iBz91Gz2Mn
VM2t34BVvpSvtGCDi0zemGoFZ+ITO5beSFa1SrXvDYnEwd9G2MV89aaNu42PWZAI
YhCNqmy5/GO1B049f6mxuspxWacHFiy7QZUc0q2ckyKP+jP4ixaXl77BrAoF1Eyy
XdvlvVVTgKJ5TMq2Trfb+ZoXv1rOj3iIWl0koBvYFojrufdzGH7yfjF+p23cHxek
KwvALE2H0Ytjz+Bucc2TtFsXVafla2yzPCJm36Z+k9LwqPFuxxRSRd6YTwKUDf6B
rY3Pw7e/9QwMY4L3I0tY/SmslXy0fBvY+BpOBxF59Z5DlxSFT7xS0m2FkF9IPAxF
USEts2YSThGe0sag3FpEtoUed+7tKxgJM/Lk+2Ie6aHa2OJ0VyI/udDWZFJnCwHs
T/PzXTVcsVRJEmQtIUfxkFJole+ALGmIeXmnk4PDvpagexvdjNTXT2KZqwjwxuRQ
GeexQzst0KVSglUKpa38PjVjV5l4WapXGNttR7VJOzXee7YLmsTXuW8BOl/2gpHM
II5BqNrLa4jKDetF/DZVPx4i8sufKDqze8sib0ctSqywy2n84IEZ5VtKuMrUkpYy
jLu0cT9UXXQwk3YHYNLNljNzIR0ndNk3Nc+SPTRuYevX2aXwN12UYNzX2+crtdaB
9Ul6GkeNlPYyALMEGIBVAD+gSYWw/OBTBZO1/IcWJspKv5h+k71PQb4lC8Wwgnu4
GsznEExnSGiQOvecyh0N0L0d9Orn9M9Slx+Fml3QQeqetBWUcYdnSLjI94eh1jJo
r5FCbzB5TnLqaSEsnN/RwxdDOxGORMYMvOtHbL/47SfWNgpnmQPf8N84GVZclxQO
JslPsZrYrQ73/xNub4Vg/OwcbAavg3p7mEp4Y0r6G+JqVUuDT4vOFLrfKtfk5JZ5
4oeV+Dg+sqjppuOuS0TrhbphEizuPqb4TbmsywrlF2SzxYITBicEaSSH0qX1ltZK
U6zTPHvkXDyQAM/Gof1+XryZ+i/8ZWSO+KzIkPu2RSt1pi3WiYQYQBRVdEdZcBza
R664G2NBjXwwxM+2zg1nFgrWtiq9qh/wYNLJKAT1vMSy29ANXRkAUWhoKlOrx7fg
YGY+4G7V8rw5gtknO8qdx6SBEemLc8NSsgxdes1fSoTTzhlXO3DIZWm2xIyk5kUV
AznpB3Oag8De3h15x+yD3BqFSbVGisjGnb6qWq+HamJBdqVN/ki6mQBdUbC3u7Fq
8TmHZXqxwRDmccxycOQw9iwcD+nQAws+fxWmw/Po8V3HK2IXfUf2qP5BE5w6Y0na
st3up342HhOXqpznEzDDSD+EGoxPdDpHh5kNj2l2niK4Wa/tc+/F+7oh5yNF2JsA
kJ6PVAIVgXpLaTNFr6SUjnZdM8Coo3FhlZsk764AvTjzj2+cPL1JK/1gpQSPIqwc
07BPNFYDFR2e6itswwgbzrkg95JLUbAKEOOey6vH1T7Nc1ElgVHGE6Jn5ZWiKxAm
DdaDA7Xt/0O6r5FEFV3+1gj3bshh9iPqAvvwjBmFlsgYtTIijx+zOcK/nVoyGXFe
uRsP5orq94zGCh4UM3PdUxA/PzRJllldFRLNXUB+4qiwCYiLT5LtUFoN3wEk4s1A
1FU/2fafC5gSg0EGR+qV/XADt3rLaDSy7xpY3uYAr6K3lfs77VtQdTvV73/tsu0I
GUQmDb+Nk8Qjgqpr4Aba9raGhLlXIgEddkWhHOChK3znSqqCzEOq0kmyznoblV5Z
EhQ9s1z514qB5k+3iO6XoWl8yyMn8ovMs2c9jPlNAZ/1TaqdjAeEeelPKA7Qibfs
Ua8vMvVlVAb0nuoudH8hWPvScBBc8eR5z8NXhrYw1CK381nr+cRZQaoaJoJSOvBv
LCzD61m8tUJyLIxmFBEtT83sTklGlzOueovywiuIo66XifEul3i70lk2iHLyejxI
Ta1mjFgD/FU92yT+9Sv2BqEzC/Zhvk6XIU5DpdeQD9ysHbvhfkSwxx1d+jcysioz
P56H1lMbqcWVo/Qtl3AXJRE6SmxSjLGZSQI1e57rAI9ot8o4lwoTcs6Sk1GCv7MD
q97IkQnkTVrFfBRbzUgc/eqhPSd/C51Nlix3Vhe7/WtDJE+ul/SjIOnflXcCnir8
KGTKz52q8sK+5ysjZDujFHrvY3Zfk5yhWfqlk7ZHCW+hbfLq0ZHJXxVtizwDC8+j
YvNqRhl6QnKNs8myAQk1so3Z0u/Uk+JO9ke1XoitCtZD7+zLjqqWML6uYp8GSnqn
S70BghyKF3eI4+89DuFX8iegm1vj96UoZNQO3EoAUsMss60Pa9DgUKUzAdMBJsat
/HjUVhQnQRFWDTl+jiMn6q19PsdZA7GuU7wCdatUEg1uuwesO+1Eqer1UvSPp30e
aQp0gclBeNdf85WM0beBaf15d/iDKUuAuNepZGc3PVDKHoGhA8Zn6Xli7wmOEPNF
x1e0ZfRPb17GJWX3xUdh7JqVYEXW+qu7OYEuFw5M2x3kAtVws99DLL/9hJuAd+Ow
efg+cwlLgkF/vBBgNmx+ZlZpPiGAmqt3g0Kt8OkPLuKzRnbSS4+HuyhlPiRQWX71
68lbSh4fZx3Vc/kr/3RG0/oV27cZaHCWDvbjpQ8Ty+AWOWqa1dTrDaHJWJfhj9dT
aEMk2eagvzLiJfbCQKGIam+yYBSXfD6+J15WGQ/aKdu/e/MGnSn7opN1B8WgGNaD
xJ0ar+c6f3M/47p5w+H/wcfbOopUX1WCaEH2VSZttlAjHWqAjoed6K9G4vSVnOkx
lMpcUwW+vYkq2v9cwSJz/yftFB/GDNIfKMfZuZh3gflpjFVsfbO3+v8dzRRHk4aC
kNoqAmK5np/paz6Ej+BqSHVxn2EAfDcL/foOEo0mkgFWRB38gpUDFzby7/S9QoWv
KfoqaX5Ikp6zUcNx55zg36pG0MTR0bwbyHlAxCMgP1FNsdca8rxDI9tuGJD8qY6R
n7n1iEtlw6Cnl+sL94gEH1SKQqxKkkT5czN9o7fQXulMedliIjBihTCndXEhJxPC
D0fXu/lRZza0UR/LkqPfproE3+bBwdlJTwnGPZQMA5i1JGUgvlaRff+SLxzUySRx
Se8hxN+gs0z3AKOg/AA8SZs65aCRzxlLTzstD4NEv3rzIAyknn7kOIL83ea3W/Ul
zQ4VREmKRMZXV/aO8IqFr38hrMNW9jfVtwt5uZEVfU8KJUeLSbQdFXtwpNpK5DXB
D49AjLL4P3VUnpHUi2iFgVoEhrDnQl4LsrxPSqT9xvyWYfX2rymxwSfho1dvEpPA
Up21bJgR9mUAtDA9xd+9ZcQjOMM9P7AIUQzN2Ftg65O/fkZuKtrYeJUYDaMnUXlI
TLyJwGgMLYwMyzLlnCOZ7Eq/DVTx++VTGZ5xO7LuudLRkpqSspn6CnURNq6V0Lgb
dT3+1MrqH+rNSNruMX65kqoZBrj/cosmXDYlOPsVE9dPd/O0t1nc/SQctwrJ5auP
360Zc6U3ineF/7B2hE43Nx06yiHe/sDMBBI+tDy/Su/VdshASWbSfdwFSdHFsdnx
xzKujUZMl+xMg4d+ePwtPvq+E9YwauAbOax2p3rNIs8vZEspT6NQxIbBEVsFQ+yu
LHvA2LBD+GgsGMZuWj1B+Ox7Cbjlx0KvHZPkd07bNmTbnIxUJovuIxzI46xHqtWF
1oqerZYz9sT/49tM0SWBF90qJHgYZrgv1v5dcBPkjKTKrMZ5Ep00b30zIyTyWwOP
PdoURlNNQLxVygsKefBMPR6HcCre7l2i4s4ABIHlojkvAFQmbmY7F6XvJRjX76Pk
zTIG51ygi48o4+2ZQuTgkt3lBIElbEuxPL5CmZjUYcJyQ3b8uPWdw1CpYUfXtXt8
O3ZmT7UY9PJPp/Zw8phR2cMMgwWFmL/WdxGWs8NgioeUDZVEj8Ddg1lgpye+X7uA
gjrQuVCfn5vHlbUWbyvA3f54BmT73w5FZdUCp9V6eApdCW5ar3ZWm1GMPpTtMk4L
yGp20PxpdsxX+OfD9V5GQTrBq6Jhgyp9k/cxqcGn7LaYIJxcJ6quyH1GTvENn0j5
LoLJCZRzNBBWc5A9n/+XEu04aa7OxDclZstW7qVx5vBO15RywvxuzxJ08RUUTt3H
7OCQvSqfg9YpxlIf2vwEO2AAeSNKSlAk6y8NkWooLh+vNqj4/e031r0TcWFVYSjv
FEeBzlEgAsZgQujWGfMuxepIrg6+GmksdPo0RQ9eOh7fwXwjq6Wj7gBwSJ1/9iJE
rvPRBbfGBU9M/3YG5xOsCtfno9W3g2en7gD3jSYsT4VedwdDUf+Ac6ffe6j2LczO
Tf8vVJPy9nfzjmrKEKfHGspX1s4/RZjjztqw1feX4ANBdNgC56EE8M0fNMT0z6eH
lJlSxTYBAYeBDl1qOxJONWkFlsrT9s6xINxL3dDl7G8BI9Aa3bB5kVmDwbZyVCR6
6J7lcbXKDzgLSwqB2KPjrcb1dIi8rWECMWbbEXxGDYUVpudH/yzKFqTcoKSwmCfi
fqhrrygRxgbuT50SjuYE1O3UMVtk2YaArj4u5gNpChsr+ftHJkaluw3NEtX7SHaN
4mJvhvyOyVPCCIwLwekNNzBxEeROMmVonCKFN4xQCLXou2aDhjwLveIEjQQczcYZ
lsLu+6qikaTipdM/HOuE+oDvHepbMuFA+J7E5wkJrmHuV+oAOjxzpkcfxg3qcmCw
G+xV+hRblKUfofQXnQieYCjigCHYKosXWr4HbBvdfgkXdJVB8snwrzcZxpN0BWte
57faD86NzJhg0bw8hqLS2Hlrhg/IOAPaOREcgVYYH1WZOAfJ0iceqn6fwzCWBy2Z
UtQ79jM2aYfk6vVULV7Xkik6Wi08/u5eCF+XUlTcsU20+5pHTR7IsxgIFoFnUTFg
fB7xpzIkahTUQtkN9LhTA+Lx6x/TKkGIW/p53nWwkp7JRAlEQF2kMWzyyHVAugBQ
d+d0jAHHOyl5gxo/bTgnK8bcmwvl9FuCZgPvhRdaYsgkczwQI65+peobats8pnLT
NFh1qAX2hDX/lb8ERpOZcPZ0f68j1uMY3ddoyaN4fh2Vayt2dag2iXe7gvgz+Fl7
9HHQJjEv62/N9rtWpXcB6FmvSHnfWi56FEYlIPmKzXOR5OYVg6T+eKpycqLfB6QM
/5VHhAnuw09XNI5i8dXiVf/ZrCxwVEBHTKU6LxyxYZB0lWjlo+/8NGt0zGM0JPia
3NT23KScxC8X1JjELgtIPGYELOmGc3p6qk84iOuuHV/bdsL3r5dZHPOUu/YAn2wU
UNxzlFI1Oy0T0Hhtfc9ir8k2FCA4EuJWH8ylL8IioWHZNd55+E4a3hjASEdXH0Bz
HZIXYnfGAeLcbriw7MR0t4ZQMFoXCEGVdtH1yhJiHmaEa04bRzmQidhYUIO4hCn0
MdJToP9u3vSeV9s2RlWKQH9OTY4LFrtFozR5eEe+kvVNgGc3xGV+2qUVxq9h91n8
P60/jA3SGa7++oZSkWxsIkkOr0DvyDMSlQ9CMGZftci/MSFSaeFpwKjJFhgPXTrv
PepGhhuPhVoqKZnp50lvxyJHfbLHGTPfxE81PWlNK2UazdR/6wj5QuCg9PhMT87r
7768JcLEM0dLBqzkswtsNED3wOnwOgv3WA3LUerwHZ9EJdhgYY5rqihu6Ti5M2E4
o2+2bqOK0uORxN2umIeCxnG1EaOaQt3v1AjU2x46H/Ho2VfatiCZHt66V8Ckmmd/
pJxZ1OWETUjN6mnYiNXnT69Iol9JXTngxJu57XJn0C9z/iS0tXlw8uAjo0Mqr/5F
wQyJRDKxId4nMUpV5RnXEykQC/MpuUdSKUcTgEnPbZYljMZjT5TRs9uSHJPC8+EO
FRMdZOT85HkPcHcaEDttiqQME44lTs6W8R+JMao7DWgkQNMkHqw4yYtJNSL9iYHn
XuCz1UCaTWPODd908B1zDW4+UVx8oVMj0fluCBu6Es2CLn/P4QM9T5ksAd/gsXqU
aV/bHx+GRIkD4s99aoAW5zQVdHxkJbaTKeVYToTSjDcw+5OWXLA1lj18BTHzvscf
+xdpuKuMFZOHK2aoS1s/t33cKRBrXy7XXxIjiMlCh0Q64PZGbOEhdUCSHpze4uTN
JEqdjuJph02NVTSCeErek2VC+5sqKbJy//9lDeBOQlFQ4u3Cq1mDUnbPZLHFCPn/
PX+R5fDGj7YY2skuGUQrDrfPjpbuaU1pszrcVp2ux/Y17xLtzApiiNiT8k3/MBrd
PgdsRkq57rf8rK90CuUCI5gUXD2+6shbt8mYaoIi3rL8rXYOQjB9CpASjiNjx4U6
R1KOXvXy7E5I+5yHsNyxnmFtTrWd3QnMLx+0y4XW79lNBHptmaCUn8NtQcSnP9iX
woS9112cjUUJApQyNixOxsGhtCfPSIWmRnHFOkRAkWvS24PrIkwQ42HxBG+57vlK
IdVdGw18Bgiyn3CkYRGrVxGSgqCLDprZawh0S0iuYH/Mm5KRTWtZxSumJi88eJ1J
AFVp+vK9UCm9nyR31f3wuXkue4uSuKjhEITjJ0rrTZKRl9zcDXZGcI1QBifjtjCs
UThWj5idkEIBmYLhMflyvLuTlQK8QAKrZ7lYUlE+YjHhcMa2owVd9BALUYIFlzeb
ZD+g6OVrnshY2QFJ5cZkqq7i8plUjrEKuFwEYDew+ugCmDBeGIzxX4GlobeV8qLU
AyYAhTJnAITaPwPtoOHev5QueHb54ovfiepUdBXg8ALn5J9BgNTWYsBlPWQSsLXn
c5b72MOhYzauD24kLcZmAY49St7IashbE0/FvKzPmQPV3xozNY/i8XdJTJZgBZCl
AEZvDTc8c3S+S7Zechz7l4UXGxtrDNND6f5eQGnmTgoinDzvp3Wti/x3ZBdb9KsI
s9IeMbriAFQV3ZxZCfMSktwLxNWmeRMrgvjs6NgYVMyVwT1CIHW04TqmaCq23WsH
9j00fq3kqmO7c/l7C8/W5qGzr5KrfO/wX5QZG3xfeRfnA5zdaZ9cAWRRMqnZeonV
8Ww1Z3+z/N/Rny1yjKGKoJKDI9dR7NW/8oE0gidntils1huQlrQSrzfpn9Ighvl3
xxTGl7a2KRCZV1c3ouDqjqwZZVakWWXc0DUgwE7R+c+b+V/yjsHY6lDGqZXOLzw8
1rQbP9QOr/FvSb243fbw1ehHnuBglrYVVNMwXusYdsBQDXh1HSeWwBVlf9L7+eWU
L8zlYaJTyU6lSCYU/mXxpNwXeVy7ID8lcoIhoLq8IlNmyYSnxdAuF26iHl2N7ufC
w71upPcBtujcSmqbBf/ocMj1Ljbu36itDOQHPALVDpgbl05KXR8PH18InFM0yLZg
jF4AHLZGMY/mgOvYv7Aqbe3D6KoR359EmyfN3cXcs++3PX3NRFLAw5oJ9+juDa0r
/lbmc6iWoxfDKOoLUqn/kLrdY7LgYkV0qBcu2Le+dUpC1y7x4wMTGvavs66CR/Xv
j7UNdRMcOIEkg1xO9cZ7DWqXd4RYnz1Rot5NWjf3KGLnXfLuiBSeBwp55SODUZ+o
6jzi4j2LVz/bW+t/OKOlFQHalFUYfNLfXx5M9o/wFltMEEblOtozMiCJZ/Eln7di
sVcOF9oAX/nr5iKhdy3G3vmt237bEeJ/Mi2NwMC75+wzyfrhJ8TzJUoWg4/upd/Q
a4O/g7Oyl6lf6XZgRwWq7OrfclQ1K4C4xGbOJAfMs1JkfL7IGrdh0PE4xqT7J9YY
7IaoV5JhixbsYKEMp91Uvi7yF21YLKvZUK/KRuu9efbG6U51qw76EBiEJ8eDiTm2
lYlqqHf6G4xB0oULBVXRC7WfCtR00jfvJcrabAYdzQbP96Hsf2EndaAZPcsON5Fm
vav9zqcPvcyN1irxE2eKNq+Hw0/K2ZaG7GgRCvG3SSk7YkR1ZVV6DdpiF1iVSsds
VZc6brhs+mKwwXRJfRkoTgCdkl0iJ81GfHDokxbw84TJYtvGFXkjCiWAKyRcsDHb
dMgLP3X+lbYafyBDgsP4sFtQClWjcTNRcKdEKTzxaNuzjEX0F8j789IcdpQPQsEp
BLhYOAy+DVKCoL/N8FcyDtlwJzawgFcl3T31iYXnk5mc3noxchNEqt04HsxLw26b
IQOes7j2cnE7/PGLBGs90dwECBKXF9yUQJL+bWMmCeNF9cnZZvtVQ8J18J/2q4bP
3KCAYXkBj+Bf7NSbtl3bNcc1kaukhgyNnCMHncYboJhgS9RWl9sFtraHVhMbqFAK
Fxs/QOP94Fcy6KKTZ5LYVavh1rn7kL2+hIFIbnuRZ+2TUeq8IJY3j7HhfiFiDMBP
szMgGk2oNhsFwx0hvoDLG3a0ZZWpUST2ehW3GR5UPktJrS219eLKAEJJJhTpmAIW
Z6hr/MVVuYyg+4LZx9cpGd5iUYEJ8Quv4QHgP5KJNd7oQ4kog54fnFBXskm27cv6
pIicS6kNYO70Oi8l9kG/usZucoe5b2Jl+4lnUrGzPrVNWO1uztX6/cJGcTKvBvmp
3wQkviYLuSCqGcEBL8HtnoTUvV03BJLSgMo0EZzsa0pmbEb9oIuvRcpRs7ogssuN
LVvNy4tBu9RtEuvNPIUVo5JXbMgUWQEaR9lWzX1ozszV+GfraP6+mKWc5fFBZ3TF
GGNKbNV8CbaIFO10TENBeybk6x6xd7KEaweENH6GISYR1eM8BO5x7Ml+cv0+MISu
vhQsbUlCYT87JBd9PAmSFgovKisoR/YpGSgiNJw71ag+f1GSOO7fln7tRCnTak0U
sgwisD3YIJBVX0M2SJDTaEWGULl5iIBwnVQ8wTuBp0arxPFeMBWSqFIlwNc1XfEE
7/tp+E+2PLSJEmL3cy9+AcsRARqTC2m4kJwe8RS1hWM6199BsyLE20XFr8xlo+We
ohqVNXs3ZfIf2w61bcnHxzZjii+IXxlsmsMJzqRyHNhmHhTBdvxJ7VPpmon1Y2oL
p2hnHX1cyTTvPL9lNHFDtP0zVD1WiMrLI18bvPB6ayz7Yg+1cmz57sJjVbSB/rcr
Ywv0url1JXVfrJmoJUEelKXfjj3mUlBTEVviQ+8pdxDk2UyrvQ3E7uk1Tov6qBXH
mjqWKMtQAa5sNwRt6Zef1nG//xR43ItKMLLlIE6Vtaba1JgyGQ5RqBnMYKer/D4F
FCQqaqE4x9Vrwrt26doqANGAhHMUX0ZBPUdPdlKL0y534rfGYOzfZ82kAwgZjxzP
y/YpALCTQxYQD2UKN2YFff70C/eY63VQvFCdW/MKQlqEuksYZGjYQJHJyUOcIf9m
7/Ha3ZU3Qj2kO0xADrgitd3MyZXFUiiY0ArwA3QluuNTRIMOFIljqmA2PODxGiuS
mNrCqVghhp5kLzzXqs+W/+u8gb0FYywTr/cTX0Oye3wrxwJe+JqFZU9Ba8tZiod0
O2YYhc4rbHN+UYPdreUWnspMNADELAsafANkeJ4YA6knHIvCWv7deToYbArjeH3o
opXnzHBKnm6f31YcKn+94sEChiLX3HgO1vujIHjOBqg9GiWdxw49r2WmvdK8i8ZM
e17Zvp2qTmGI35zAZGbwqQOSyw84dXbom5ae9Aak3sajEFTpOzPBty5hnCNlg2dm
8dvPwrnRIIvcY4LdzwEAzY5dvjbOJgEyC2lVURS7qjCytIRHY+Pf2ZvTgoNkLI8o
G5DJfUJOTdWvSi/enw/+gsl6775IJmu0XGKcLiZm/8nVCMqIt3tr9KLoV2AnQaHx
+UlTJJ9CP7YI/U+YbpBAMLBW7VWLKvPkuJ5v/5YU1W/Jnf5n5yMd6Q7wQeSjq/rj
tpQiqOvTiW1vPDcbv25QmhEDCc22E7/fBCKGbEmdhS1b1CiRNVpKZfPdbWyQ8r6q
7TjN/AB1ZuZjgpxm9Yht7cSI74LGDznDycupfj75VFvOWtDgyQ+EcribaZOZG+ri
8xxBGVZieYBlYB+/SyqpyfoEJE6+OZDDriVUhBrxBrAIJNyVzY2R2vKUFgUK6u5x
F+sPDI6b/OV85NCOx8iOpwSmXLXgE7m3TqHSZc+QN87Y72GdnCCPS/a6wU7sexSf
9ZopwmJLHdDTr8ZoDJGH+FWLmOXAMTVs1EXiA/FM9wR49So8zv0D9z9ZYCbQZ9DJ
yNgFyQVLsjfPFVmP8rVWI234+5ccRBU8OpF1n3R8uKiaAQUWVyFm4McOu8TYZptc
KTLC8AAz73ptA3j+KRtlRMVUDPcD51TeWa4A91tgIYWLGM9Lr0GPDYEtulEDFEtf
vbKEPcmJtXqOOoWQbfz66rzg5ZfJGPsOPRjcT8y9Z6IwA6QGYBRXUuxwWUOomJ9a
eZa5R+E2iYjDiy+8Xw2+dntNiqtHgOCpDb8JngqkD+E3C9o8KFdomWFfiBOu63zi
wrnb728B0olgbCOey07HEouqAOw1RAYKjzlgG+EXRXfN27fcNPA0ueyVDeh9ws2Z
SN5mOLJXwPty7LBTxuSaa2mxEczGU5Pe1bZsOHzmngpkVEdwSrBhXI10by++kYAz
q+zCHXaTlvxhsxBzqSA1XZxmITMqtlaM36uE9GOtoW/t8biEr4HuxqlLkwio5i7G
Od80ItV1BobQ8p8CMZNRc7EpWIuldKYsGKkjlx2exxdSUAs/aNwuAT4SjiHbIEIW
+kEeP/r4+p1pWAlZS/02b9wfjC0jyVoPMWbK+jdWMB5RgLVnoZOsofRl4VLymqFT
tYS/LU7hSj1GpgDTmeYXxeZEFSkysCt9XUDAgbz8n3vVk4AIifingeVktrf1kWng
M7Y+EArNLUY7RITe39FsYuRGsyj8P/74bveQ+V/kloFwTp7PneaAJdKaoHe+BWl4
aCdvt+Mqw298EDjMLO1OcKc54k0khyt0v4U6CMp7OeYSBb5DoCLB9D3tCJutRhHf
mHfPBnjElHcLooPZlxkcdDDv6qS+KlSo6+0c3+v3msC2m1nFiowqEjc9bUvJOHjP
FHWp5IC7U6D6dUMgDR1VlhyjmSkjNPE1WO/tTCS5Z50dQlKO5YPliJJolUdOWT2S
X9PizHr8UcsW2lWjkdDf8/kb22jkrB688W1Hp3VCgYpZlrZ/Byg5WvvlRHm/tltz
Q85GclOVqBBsTXesTIQKJN4ynuvLJV1+SQ2BdEkvgdOYF5cDMlx53xKdwYI14yxp
vISG9ZSJAFK5hzx5bIsHDEFcR3kFlMKJahFXNqVFG6FM1DwS0FRe5jk3yOIJ9edM
FqgvKs23ZK+SwLe2sboR2ntK07OIXI8+yanXaIMN73a5RcP+BG+nDliv+2Af8job
6/YmBQwUNnh6i5R22Vm/57GiVYXunXRBOu7iDQ5gZ/AUJMx/qAUHucXftAoO48di
aI0K0xjJlrkjfB6t07ERZMbmIcCkLCtIkYFjbUHk0rWV+47nYqgNUaePkobHA1Vm
CpzVvILNyskzyve4EGVVPapBKcBudmAYoQLPlfTaGKLnfja3a/ui/Y5cd+SkweHe
Tu/WwjaKgEX4sjxDQzEkQQkFX5ljiu5SBLidlCqmYsm+7YmZH161Zb0Z+nRe1Lya
1S/NO7W/eEk9IGPSFOnX+KBFpQoCJmsHIJVgkIRwTe0cimAJ5WIwDVAow1aPmMtl
U+Xxu3lQORuBdZrgsT+r71OzJ4PbWfrEPht5FcJ0pninvKpZipJucCYjBQNkDmds
Eka+JhUQRWg+v7L5TEaNjurb9GgcrKjckrfksRBRHBAKqAU76Q8lFfH4+wSHisn5
4cF8kH2b9h9zd/2Ue2J/ESaqsYKG0d7yY36SflzlI8GLQvrSDJd17lhKdZBZe5dI
0inWhfmOnOJYNbcykpS6+w9je7NJvg5UxU1pD7epPlgPpAsp7aa5Gevq8gln40IZ
Y0Hb7kwgB/NtEMXHY9630U3VLyH4Q4QwrVeRzWsq0C+1wE78vCAYMR3PAu8go8VP
dxHHbn0DewsbkT1pmQrWG/7GKQow3UOvM4tlMzufAt1rNhpBg0XQmihw6/2e+9vc
PKQwC58CrfBZJ0oU5ty0295dpzfqLBgtOwt1IC1RFZ8nf8NcolBtr/+O46Fg7ozy
P7r9W02tljDD7BxEzI7fZALI4JIK6hXogDCW+y7lxzKdI9gugCGB6UY3BQy/XlIt
qtsPs25Hzq5q1sL/JvZtFHDavPkHJrySoj4Dh874nYA9kw9HtL9unLVr4OvkJ6xc
oQVEtnG5EOwPoERSZZ95PCfdVCOXzLvMjUCp4BgO1cKPGzkBjKUvVinw4NTKpM+j
G3MvVb7CKEhD2BewL+a3Vi6SCGXUShBgJElFCvIk9Zb4YmahLv+hmOkrwQEncSxp
riedkYZSJowB/RxG8uSSZTATKEcdS0jAg9dDHq8i6O5fzaJEL0eA/CxKFPyXRr4R
8R66Qxa5DeHiOetzXUG1RJd4sOeXmVZG1RV62Dz2XM/hrYjYMX6p+uFPlL37RUrg
X6yxO/s2gXxjg8JDr368Mtvjon1ZycsEyqMsv0bjeW6c6UczbsLulLC9GUsl5u9W
AA5ual6K6xAVaz1l0T/tOpkh3gX7nKBYRsREYzfDWijm0uj7qG5I0XQZBIFydU1x
ttLSEFw+SB23GdkrVcaJaKsI/oz7zWH+87vLXddTWtLLCBXCrqncmvnPM2olkcu3
adNEQWWthWCOda7W2cdfo/gQTwWRxo1qHheMpppj6LF6Qi4HCbYpoMM0ztQnaGmc
e/Qfmv6X+XqVy9QsVtgeF+YKT6a5yZ7AYaJdj5U4La0jaS14uYBlGhZMhPZHpmtz
aeMNfp4RHvFV8kb3GT4o/uFlqMW/+xu7CyYyknFFf5ouZNdv4eiXwcTl4sq/1O/D
NP34JfoaCgInvcQmNWrSfTAvYY196PtLRSxWFePUy5cwFTQ/mPttyiT7e569967T
DOUPNia4ZteM/chB4J+WN8mPnkGz6uHZuGlyIAvKfHF5gRTqgZ8griBIsFQEM/yt
R46+L4JLjRzj6DvtXDcFoGiqQUcQ0X5N5CWevHuherPTe/MYyFn2GLnUFAAUpPqs
hKEpNiIqh8GmQjA/xIBa7Vpqww+yEKLmW+rVBOVFB5DOfBNhycE195iVS1A8lj8B
YWINAUXZuvmg7jTUcoCOW+ZSStZ3EH/1Rqu6ccggE+BOg9OsXHzXMdHsp/J5amQt
AC/SQRPNpNd1P97P8PVJ6Ldhu5gI4im1e9qAqIyY8oWNV7w5rtlLEUvdWBiXNDJp
Dik0RE5Cc9CKnT/GG6Zmc2npzcw3kIuMlkOeiG9EJDFUFgX0FmtPPdvLBUNfxAJ1
vRjRPzdu3IH8rRHYIAXKaPyseZ3eHRREgemcwzvqCplQwLYAHvOPx819RhtVaYqN
a0eBacdj3s3gskJ2MwSJTEJT3p3vpXniUm6DCLgOAE7Zmy8L2Pq1BOAhWnitf15v
/nt1sJDjhvUnaJhYbnvkHJB93JbjjDgO/oa/r65hCa+C6aSq6Q1n9AFjXPS5tJGN
EGJkE+y6Aa/RFYMy7EuzNyYryBif4Rqxv4U4rEwRyzkRZ055uJIZp5BBRn5s678N
eoTduzziV85R5cG5vTDQqop1/E9NA3YxgTIa0izJqzEKEjNa/x8R6fhADugF6GTN
YaxvSOsHZogmBaHCPTxF4QN3bxa6juU9LN30ye3oeypRyK3l3vU6wnJalQUHGVXE
VKigLv7VdxRWr2/uqkUXs4TboChtkM9PNVCt0zm5BOJNSzmrQSX30Yh5Z81ox4Mi
1FcYqTW5ISQ4DIqV4M+EExAvJRN6eY6Bpkmf1OF1ukgn0pkmbLJQIxSSGOxFuSq7
pFbZXuMf+qmVcu7D1zydca6/h+M9xz1palaBjdkiBJXsqUCCbEZg1xFJXGULgucu
qb4O6/IS441xvVO2ZSRj74HUarAXHRokksYg+A9uZ+qGbOVyhkImCJoxIu9EBVlr
x5TMJ57ZkMSDr0NTlzMNCsDvuhbCfQOW7OwXNqReT99084HmhcYc9pDXZWlqKzi+
JxNuVjW1kYl+DPYbdkOtH/gx19fdykuNfwh6tVcvHK4VqyGuBJkvP176hC0Aao87
xAV7cafnIuusFZsiWGmwsWtZ1ZT7Zb6sMpidF43yRQtDKbBRyoCdVPToiPUwJwul
1JOl4L95jV395tu/58WuWxRjx8akQERTMPGm6iwQEOLrL9Cts5/IdkibCDHxpHGy
Zar5PyQqo5qWzAgXim3WIcwI5u2Cl7ZdP7+F8S2XiJQKejaBQU1D8rLuQ7nUXXHc
0eVkDUJEqjaJpCzMKrgYiwPPUeUDjSWrB/51obu8xZFJR6vqxrYMSaSPuP3YAY4W
4HQB6LAXrScaVHdJvvrrVIIacE8drzvPCnzTptSOGvvqwovfEbdOnaatYhpANDJK
7Xra6HSb0D2LAD5R8brUX5iI0d1VGoJxPgDX4H9XUhGOHmyvYC1k46TwZvFLIVsp
xhhmfzsupCVFAc76L2hG93bF4uvWsmnxHNHosm7+Na0m+p+hHYmNq47pFlibgzqr
ueGu6YR7cs17P410De6wEP4dMPTE9BGTu3WyF0hMZKYhX0XbgQKycFhiQEIoNUtn
h0d3LRcMrahz54by7l8a1ZZvimRL/nZ9VfeOhBp999xY4dBzLevoGwptPGpemVx7
WE4VdU9vupIXRR3s4iKzwRf7c9SKV+Sj0PfqwQDSo2nIuMpopBMuTUWBTnkx6w49
F/yRASfGCnWAYZ22Yug1Rqd47Qoubhv9OCqgPGhE/SlSxU/+A6QmtHsVU7ukUJxt
WeBpJe40NEyoamRl7y4DqgbSL6FRAm4F2Z+Ix1z9YXdz2XnxpDI+h9YN3uCJ7cGa
toyxpw4aQh0/O+i7uTKOJhBL+XWLqcAKTW5liFP760bj2BHoOEYOtRazIZREjxeN
FZ+AeddbaqRfIUM+c1zJD97BqhzDQvxqcDHpFdZcYdJiHcz5wRkDEuljM5gAojNL
lWJlq6PN9FrDVGIN3SgT+U3mplOu4lmvsDTqQqJM6PLsYbkhXCxmZd5xJlmbc+ac
Mc5OdMQ4A3I8+z78TL/xYlTNAh9h2G9VWJA3zSUrQG4xtxCy0D1kbboZcWpZcovz
E/gqBl3rtcWepPQ0A9oSifb4gzD3l68CocytE7z8JSLWFBvrI6TC8yxSnE7GQpw/
jOxpdcRpeMq4+MnyRoMORvj+BFO0QX1NIYsIepOZX2B4AHxQ6Bz1/w+M3EPfkpM0
kTqmQE1Sz4YO8PBc16I6t3YdNa382OA5jvNCuI77Y2FXPtDuamq/CdZpGtmIaBs6
2rqSPhVUYwBgLEOCHuJt1Nh/dXSABrTFJuxtHUiD0WpYqKCZoICfxZzAwpqRBqwh
YQpScuyjXDkOw3VXnafXHDPQb6KfZpPEWOoJh0dN5PlJos+vWshtC0n/0ycvbf9Q
1fvqeffYHWestDKM0b99a6QP9UI+TO4IGBFrAGwXUg5w6EcR9p/OqX/ywl7gdHpj
0LfpSd0qYGeowXhs5Z3uvzMFZDvkgv5kTNBjX14bBP+tydrCgGDtluh9VS1SBivr
diDsScd2TystAI0Xbz5IR/F2GAAaZH6UoD7o/AN4XYyDmjM0qSqI5zBq1tHis6e6
TvrYglVbgcwCKL3eqn1rKhYKsuOEy5dHrCU/UE4ux+u875HxBOmYx5PJc1+5hL9P
koRG749TbsWmcVqZs5BISf4oMWItUH2wH+7W2iP8PXwwX5RSS8tzpSSiHcQCqgPU
K+/C6nnGkEHOCzYhS02v8zjsQDc3S3vA+sjgwhzEEceN8mIoK22+minQJ3rVyEfL
Abjk0Cf4Afv3yJswB6k1DNjIbtmJjWB40RobGqsSpxDUEGDmovXp2BGsfxsY1IFh
F6LZ9pEyQJ34SI5gXOjvgV5qgOTa05V1xIjY5G2llaxIXK3C0i/qllnYsniVpoVY
mQ+8hHNMRPjVmz2peLcnJkdgFntCySClwTCZLY8QiKexh/Trj7MCg0yn/w7xSKiV
S6OARYCdUgxpgjIauf7l0XeUkb6Bsj2Ktfhppq0s2uOIykyOF1T5J2wZzcUUeiTN
YuGkIwJK4s9z/4kjle1YRMO7Fp5J2yTLVyNScOofd3I2QfqKW8aWmFU0AaiX/x90
es4BFKLBgXiLemrQcaEh3e2ozXOwB7wRHc/SQR+FIng3RMY2G2jyZF5329fgDwcY
xWWJTYIqT8Us6+97e40CUDv7SQqaZKZGHfWumPJA7OO4z6LLBh5mSSAS0KJ/Gulq
BWzKaFpum2b966iEUT2EamxBvpwIVaQ3xI22lqFXL1ZLxtIb1AWa+zPLbplaS73L
nuD2DC5A0CqbPnyDq/MpHiHZX9FBQmE50SNdH03KZeZw5YHuF2BYT26gwRz1xTTC
tHoOSgMcKMP+Oe0g/FtK+GydPdQd568ia3RllT5F49QJMSVznO43GRFeGcAmihMr
vzH/LAYv7ZDJKOsGeITlDCdhL5NfsLh5bqGSp1Ex5ChlkwDYgfGC+mN7E8EkpkSn
6hfQJajUzUdX8Z1KXhyLtASbWfbVvHKpsoKBVyzGsEaFK+SmwZ4m0Nlw+s+Ko1+3
pd5rLOGrUnpNvThlcFdBsBAIjEZVHzCRyEokOrOVaPbD8V4ju/hptxCHdkzhpy7j
uOUeHiYpxI7ECYipFIvvKFiqQ1LaOV0EQDGQ+uIiuVXlSPc4K8i4+j4X8YTpMfED
7uDy2vV+Hmys+MsomiBgdwhMoRESpNo2lrtuUraDTPeXHxZvNHlgEjsXMmSFn21+
oz5NmlGuGWlq3ZKpnD1bS0Un5X6yhQR8NZdquIZN+jA5JHviwN9U0qgmQEK/5mdE
AP/ea3ijZLIqq3SNGP+FDcdtNAtRbpwomMTlfnrCbdhc7PGMPCKZ4YB0SI0nmyZt
4K0BZKo/UIcoBxO6iqCcb/v36oq3FEqZ2juf+qUuSwnq/pSI2XUN3W+g8mrGAxZj
h0X7VF5Abe3evS7Seac8pilfytHRODwe/dOcyeK4oUnxowl30PYd58bblDe9FhLc
7DcKQNd+MrPVdLfPJ5iwKjA3FZEjT4Mbcy+M0iMw7HTlxYTvPJdM6/hHFje4KhB4
9kbuvgQ3KEewSaLnTqXesL2YR6YLfjP1ql8GTC4K5SXyWOjg9OB4I5OEp2NFSvGL
TwL6SBEO1MVY9PDkxwUQs6UIf3TP296ZYm19OZtG7yD3jbYGzVaLS/4nvlnI8GxR
wqhgtieS3A1Kg6Kirb30Q+iKl0Akn4F8rAjmK8LxZghcNNd2/yYiYiif36J4XtOJ
CS0G+Khdns+ufxy2LNZ10t5ZDxIIW6McM9dlVG4dIddRmMUUEHT9cRCyAZ48bKGf
1XNdKzUHEn5lnuCtmFkKIt66E1JNSdjVxHYMaU3reXzE0Ck3aIV4E/NhR+c4AI5U
TlT5Q5ykLvCLFnmSCZq6IYyRKghCAV0hbBGz8K2TcyiZ+Zyco1uqme7oZ+ikS1Fv
5j3kuUz3g16Q5rvPmChjWpV4Q/GIPnE8g/Iye4P+6plaRWvLskDoPBl1e0YdMfmf
zOlgdF9qCUoMBf0JFx8YK1ddjEIPuzLMLsFO55nOFropEZGb+23DneRJ1RDawjt6
mHvLSEbiiKv4IJKTjXXNLydJ7wFf6YgngLQP8Bv9PRmvnehMAmUiqa90iVhvZDJI
yqJJNzKGVXY2hOeZosJu8RfZX7uc18x9lGUxb/ddybczJkCq1f3ecs5RQJNF12hE
l50cuK7Lo7n1y39N/CIIQ8Ihy3NJ+4ZZ5ggnGbl5npE7RxXolMc5pgH5PTMwquaX
uf0tJV99ij2cGSYbMIUJJpU5q7K1P9MtMHfB5lgS6Zgx9peyZ78AreIr6hoOfHum
GKdUmpmLMGohWLT/0tN7edoZY0agUrMIe7W6TNbBUizoO8O+5NxKQKXTa3ptrsmH
anJvib47OGvZG6oIxqP/jNgpK+0TH4bwrleK7F+nCtsutHDzQGLEKP9YuUp8zM63
HgTu2k34w2qiFYNO5hBMjuMQol6nWQb76xX1iODHh4yoECNLaFEM6wcqG8zrrj/B
Ty9wXklshnC8B4YdZfI4se7lAkADyVTKOdcrVxRlozyDGhlrTpbmhvIDUfmMnK95
b2ev1vu9w3VUZoooNGv8ZnMzz+H63ifwXM6Zi1sy2oqQiOoOadPt8LTPTcfmKr7D
r9nUTuyWcwUB/IoYVPhCpHncthGywSdWmpK+ymcDiiyvmRZENqN8DPgR1O9vjCFB
f+/6BcMtsXhLeIRnRC1t4nGTYqYfa7wyHkDFbH5JOsAAnbCSc6D1WgMjRmXQ2gqr
kgRyLz3WqPali6si3MTU6T0aVLdkxYZFBri7rTCtoOTVwkBxobg83EK0b+DilTSq
uKUjEfYeZEWX+/lJ+6s9jmfv7KCyotEGe+AhJooFnd6AjKEl8wRzDEJ86IhWFxgz
fZctsDkpTKDLSzcME4E+cBK0jg15S3KRZU3YlOMINIxYGuOOSNSv0+B/H+SKKe4l
JqelT2AI4S7sq/gLU423/o526LTo5u4mG/IAW3hbg5TgTof6A1j71HWuZZMnwCs+
/rv4eweDF1Ts2kRR0G6zCzBEnE5DLiuTNj5MUkuy2qT/vgvG8sYJGwVl+Dj8mxkD
wdp549dpl7ic89b+9HraD/jUPJZCLFn6RARbitXv/jmJvlKDrihwbSA9KkiZJ4zh
iSgnKvHrEo2La4tD+MTPBVD+yXvsXc1BThxyrgP3nBEzhmLo+JcJNnqUaOzwdWiQ
KEVkMBC7o4ANGaLng8BolPP8s2lqVv6k2p/RgMrBQmtBsnT+R/YotdSgJd9A1psH
D91YHrWM1mMkYJMBzGcDOHkKYbW7r0b5VBeL8ZOx/PdJh6A1m1G408mVzor0YWPy
QYkY/ggclA5nqc/2RCIn6yzKyS6qckzNA9G/2NDQuw+Sa9hbLkeI68tJk18H8sss
lyyJ3d55Rl6fHEm4lyVBcGFR6vNjyLd9RPY3iO1/MzlsnzRAIYXkiBNuhvmxq6yH
WnGCG4KaOVHVrieUSZ0BlSZCBFn5XBHqDzyLglWuhxO79ysVR13jKeRQHX1O/iXn
KAzfzWWRflU+ECNH9sJs3PsiC4OtStmZ59jfDCcPn6t+mN1VfMrUga57M+H2Wgcz
M7/17W5DL/bRJAPbN/fWgEncNhwIeP/B8vHOqmKFtubfYoYFFn/Qlceuy1fe4E7S
ShrbHfKrfD1OrbDcDhDlDb+nWPnSMLoAbKMxwH9jMWn0+XlCZijsJgMEzNKDxAGW
i3W459VkkVKRNUdjAdOaiq+Sd+2jizbRWqrXaDy5Wwft2mQBg8V/OLfrecKaKdDb
JlaTDkiR8y4AcpU5nv5rEqE4n7jgjem2WhQC9sUCKxdDUvhTZf4yoj+pjJWrzjj3
dNI/6Ri5BGjY6VundbDG3NG9YcZ6F354hMelMZPJVyTHcLwtIi8cVzq2gRHDtHNZ
youG2DF+X/8aQ3sDH9uS/HVWZ7RLcGCrCbAQOxaeCIX5EKjfjsQEFBlTxzXKi/oR
6jqnJwk4lXcXu6Rsg/JRw3RuqBE8O14oOezJTNYDlHzEFE6ywGOBR9Xq1a/Oo1dG
e6XpxAUHjPjrN5Igs0ynbXDxPB+y/GgzwEoxrUxhJbhqxuT546xhNuq11LNef2Fn
V1wc0LyvFS3m5Hw7KGPx/h0uVqeiXM/RDhjolDoWHg3McB11XlOaq25AmnBs8tNP
rjiYYt3YXLV5JYjNkwaoR037p6Y6xrrx/wcpQukh8M5tliZeNspE1ttck/xRpTMS
JZqLaJgbBFAlo8uqo1dpQYNbDqDrfxPFCJJRlJhIxNBbaiEFEGCCRT4y8g4mDN0G
/nq+GarApI1Hgsp3o+Y6Ih4s2kXx7XVoC7awlxFs5VHXVseDcHKsW4TrxVh+umC/
PHh1RPvgvkmC9fV6hAoscTWdrVElwe3BRHOdvaRvMSxDq1DB80yEW4A8lWeUtJl6
hRlVo7Ym6sXw8WpTYRqybfeW78cxN038xreoU+Hb190CQ8F7abSRjgSvaAXKC38R
MS/woIVxTGdYsncC2ki4LXHYgrqINCKkknPUQ6ZYaJ8wKqw5KyILR2ASXqKBm7cL
stawt0LfsL8pbpdJbm39ef3pqiLIYDi+cX9HNx01t1WRTyCAvWGEoxxaluJ2UtFQ
i630pxq6PKmJECttYU84aKDtj6pxvL5ujMMQ+DnirCVC6rigt+lmmH4NOKmM4qR7
KRp/+GyUcPBExsj5IyaUf4OBaweYEOzFgkhi2mUeDViP+JWEhOk/+uqvp4wdtNMT
ch8Q5GwXzOAy2duK9dkrk7qUriXCQQmEorT/oecH3DrcSDeIs/lvSEYnVarx/GlW
XhhtggBrj4/KNpsbn9ZjCaYq2xKe/jNqdpZ4vGQ0KeX7xEwtxZmrWUAfV+9p9Axd
b0Y3CQPYh87yReEHibefj64zHO2aHB2eS6EWXaNdyk1ebhFQcBrgM8llxCKbu21B
Rei4WGSeK1kr/ivb6+v5zBGARv+4zrBYUOdX3GscCgiKRFaF+3C+ltzf5mnnxrQT
KBA5iSCdvAElHKlPTEKQ1ou2VWfQWpA3MR2/OIBrWXZBVc3P0emNDeRPg9fUc8PP
DnukWs9hwlxDlCvI7d4+lXBBbvp/RV6UsCbMOFUrL96dfubU7aFU3X1gKOw0XjH7
O0W1DHjDktEDYtQgoo5Dn24sGklf8pHjdeUtjHCJsudz3pvZeG6qo7iMDl6w8PaF
oPmKCK0bBNxsDOXlZrrxSyTDx0Gvt4moYT5CFknRpu4Z3zDBSQL+P9s4VcaPs4Go
98ZguEHx3GMUjlvHFYB0wQbgErjb8GtNnHOXKMadikN5sE2MNnULr5CMb20cmOHb
ORj+nuO6kIuIyD1cgIMvBWmuRUqNxI14pPqkZo9UMOu01fQIOUkMNp5lCTf1nPUP
cQEcNpl+fj3BP/Yi5mK8FgcXRxKjlQ5ec6eLSo4R1ifUVb3GqGo/9A7Dv4AhxagT
IlhMnH4dUAQX4TUOAuedWx6k+tKdQwQcYYGBsxK5XFIqLtfX6FxMxq75D6AECJxy
Vfr7VYDUEIiedaZn89Vke19rCJ59G2CsbhCAQtgXk14twCKYFvW5vwbzfPFaEZoU
S7QIpNOqy0grR6UQ1+MMZuEvmGOIGB1yjA6ItQLfjQbspMPcdC1PtSsNNR7M4Hpt
TGnpG4rg+0YYEu5wa9as+rRfUCfmDD08l2gBXVfrMXNbhsHTqb0vj2sTnVSD+jW2
Xp0WDNIx0kQepiIul14zriTeaHUmWeCFNJv/h3AOUOSCmch+g4S5dPi8/KKEtikz
VKtvweZhWxosG6JIhxWgXqiR1p2AKGF/gGCMGtNSalPjHadA3RT0bxKupDAgXbHQ
TLiQMQX4z3dx365sxb0lorEFLGi4bnzO9H7wrKDIBDgYSbiHA0eYPCUOPkVjtBxP
7zGh8OayixQ3Z/S0Sm1rryBZduUmj5psWQRxfDjNk7hVXXokE/Ia/vRPWHIxph+3
N6Cqo5RuNvTgQlfALVyvCWm4FzH9WD8s1RfiT3I65Aoss6eqQ/jlw6Du5RK+QPT/
UGYQ7WcEeihOXTygGTfC4GGMqqKj2e/FfiRhUAMkGsRtdTpQjD4sRBpwUy30yxDy
cgLsNoRQnwta6VUc4xpkp/JX/AIEnEeyZ22xtX8FW9kX5sUqsNxcnnR1EgxvKJjY
P+dM7aXoH9EIUefC9WqDowfHPK+/jFdfMgol/JsQy7IoCfkprrJbt6VOyets7SO1
Ua16Md+yxum/2j7IpDa3IF9XzH8oZPVSHzv/OL+f+o9XDKIa5NahsJA5CAYyfdjg
0iwcT/9lVJntLmxHBkQcVVoDQmduJaoWYjlyq+Otspq3p4ASnJ9VDjxq2zGFLB8g
yeBma9A+XMAEO4Eu05YEAqTfPPUD210s4Q2sP22mTQpJq8tlZdl4psLkT69yR8SK
80g/0aK4tfcLWE+VZ3u6EsF7mGOAPkI5GB7Su8MINS7FRteEpCLgiYF/m+6g+Ac3
GY6bmXMA3vxFK/fLyGsOdG3yi0tpO03mcMq3lIIER7mWgGOsXIPvoBDgnhNRvGOe
qPM8i/YPqObriDfkfCqaU8T2jCbyCh0let3IQ8lTr+zigr8S8Ijc36OfDV4CADkf
TIBpk42nhkYDGcc73Q5Qzhd+1Fux9eya89AqHPM2rKvtSdM4o8Gjlvh8LzfuBFHt
BMfkL7C3VzTv8S6+dnJ6ZA11grj3vZKND+KNt93lshnyeZh0deQtyujWQA6PFKs7
Bfifyy5BJRtI2XLmWB1nIxsLVi40sL4O+iOylDFhgX3BJg8i0d5bLooR66V0nc/M
ajxSCGP0kj8V1ieN6/cJVgDVWmFPFfDtxOG6bJ8+NlfgLo+NPYYAbJ7NvzfojvaO
JxpfF/ycqD6jnKG7B5lKzxHrC4JYMfVQhhzjk+PhBigrPDPkJ89rMoEIu1OQEEz2
fcLWyeWv0xosQUvxaaeEqFn4N0FgPlaZK2oVv4nv7aU4bG1TPbeMxbqM0xjABciM
z7XGyl+CI0nKlahDTNt9v8YAsJbJm1uHXZQShwVi+7OJrvD7oYNwTIyLf1ty2ijO
Ng1LjAt8DijEosNi8WiT2D9PPS1R/vO+X2E8Rhwv6kK2jXs97x0eeSVUtfYhHZSI
oo8VtbBIdxqfmNvp18QQyWupxm/F5/8c5FAMcHo2LBC2+ywPEJ6SG23cEeRFF42L
sOH4HksqJJlXiwBAFasYaKcZnfCOuuK7YvDo3GyJYF2jm8AZnBzDnDJK3PSDu6+k
8fSFB3BTr7U9i6yCk/Z51W7nCSQvO1GXlA9BFyT0NmxJooRO27YYnDRu0qjrk25m
lhnMnLhD3yoZQgmrg05t8WXANBuzk3s0JD3eZlNMl27tgVy7wNjcQvZxtePLuMYd
vMqiMA+ByHb9JKgnt+VSHCQvAqcTSmJ5M5HYa9EqWSfpY1/mANH/pYvtcBa5mFMY
pAqfD7nVhqUiadfIhFAmpi4GpwBfz9076P6mZaoAz/HW6eAK2CcGcN7AFE1g5IWL
Nz0X4DwE8RveLRvnAS+G3Nb2zAiJkWapOHRz3/H1rDMGpxQvwEsL3fb+17I6H2uv
gr7nEsILEKGidNfsXIq58Au1AvJKFhFwBq6bcyClRzbpT1LD5TJ02KhWVMiWldo3
0QERLuBRT9JVaTL+9jh9yV7uP5YWFJL3OOE3C2g5/RnFbFp3dcAmK31Vqi3xB39w
19qQFJm5ThbZuPQN6W0EDZwPhi/jEsZehv4M+uGezHuj0kf9xWn2b9Akd1v8hKbj
eBzsjNmwgTe2E4miJqy9yx9ncXghVb1XdwVP2dKgU1aJXXbo3QuICvKsfiXUY2hp
ob4pgjaZmCprJObYLR9aY17ety+7eTlv13p2si5vIFwS8jJZiMIfIZcVlY+U2x+g
xng8LgoM9ZWuA7UTqePYPkn6+HCSnzeMb3fuDHNaMVMenokZ0rLfIijB18PM1Ft0
t9/Tp9bhleTWb/y/4h3y43ddaj26vnf4334pbLNb7QOSqRAa8Q0KVogPvQvQMoF+
POp0mv4n6LWVXT2ARHZEuJ7mhq4rurGzCMgHo0eUKu308my2BoIxdQ74yCJbgMdM
gnJvUMSKnHj1A7kRzsip6HrNcgFG1liLAPGagtD/1A7Y56qUD9WkPQBa3+NRllvu
wi6+Gta+S4CQEkeshvTJWyORKJklobgB8wtytdRDFZ5bU6pDam3ktQk5HwGaQxF0
f+Bvzv/DkB88vC8uD02ZjU5pxv9w6dXoGowMpGT6PiD9IG4f+UMaPIXIz5NEFUAf
jvxUJo2pfYIBeaO1ahWBEf7Iu8MrgBHuIGnHSWmFVMZC+FTcNbXAmD8+X4rfeUXY
xDtwBxZcq75DLHWuD2rAhDklLXQXg+rQrrJ3B6NyafLO+mS7k2VDhGR7c4wsiGkT
78OJ1rdqqfAxjFYBsC7BmUkwYsKb+tAuiz+vIU4So221McXeFwGDkU5tJUtge6tH
WKC+u2uBfjRQX/v9kNj1F0JRdKpyVgqUJAMQ2kUkHUENhO8kSL0YwNFe7NMKd0ft
F7dQQtu4XDK7i1ng78BY2E4mSC+oxW96YsreSuRHQzLhGrZnx8bj0QOAXZACEtjk
HcuP7XjZCgmTyixQ7tC4J1W2jj9RPCAtMOnqZtbmT9muzea0VOGplzXqlH+C2mQf
EmaSlKVmzPkF5YZ3Aag5Lt2YzZSvCHUeJhzsXsbThqP6vCU9aEFx9vsnMXpVdRGK
jtLEdIkEEkXGhuvD7hwaSXPrhtg6wNn2ArIfSORPFSSYYTDnGySsSQ47Len7ukV/
3BA5ko4vt0k5dJhpBSj/Ed3wQ7lJinJN2/+B1s22s/7WszAs1hQcy/ICvQiVBqBo
R7QrcMoFTdqHbVq5FuZrYNkt+2h9nyfnjTR+GfS0FNEmy/x38w/aJnjQv4jFI7XL
Jx1Q3VrtmFWcysqXbc7ZidUIsDAp2Vuu5HyH0f0aKwBL+9PCKh6RCIvkPtnd5IT6
TpTDoE/j7m/lRRf0c3YtyWsC4VLx18KIDY5cUev739OEdaIr6j6knWWY2kvyEIH9
wUdwr0aZUs2NclhWzcwIIVYIqmtjTV6UngOP2PvDzrHJ6cMyiP5T+XwbkTWp24p6
jRQlXioxHIa1yEhesHI7drPPX8ePvASEDnGHqk3g7kJ7IFZpi/RX1TFNRFXYI5P/
uKVMAD9atXgby+NyVEskC4bSxfPhpwKQK8ahCt6lM8fNsnRrxkG4hWWk3K1Y7WII
1bxGn1LvIZijTuwrWQ5Qpr+CiI1GrgZTSW/ji5THIqt9lwCljGB0kX6mNbz91hct
7IyUqT2QHf260XN729cq5AeAbUjhKel2ADBxaEdAUUVQy9A1ZlVQlwHMb0ewssuA
xQTYERUWPxeGJMLUOiuk4n5Yn25H4W5wrL3we20NdL8ts0ggo5VKyxrtslbGbdHy
dsG9YLr6nS4lxzD9KC3vH0d4M4VthZAL9Wj7eZgaHOT+6KUmowALUDGzx8QrM6VG
9NhNISrgFT5Xm2/MBNhRq04QBRqEPI8xRI/izXhClsP/r7ZdvA4bWoU3ddJjT4fZ
cPfmYDljB2Il4JEs0l6MMqajK323PynlKU9uW7HMBL5tYYzIBfidjv1S6FTAQqBV
aSGJ3p0/eT+X64QbluHAwjfTLM3XgM8lxpT3V8zfYG3FP1jPQQiO5fS5AMJxGVan
l8bV/XiRUIh8STrdYit3zVIUekllUO4s2HlTw/kvGBaQEOU/4/gAb4F4QZpo5Ysr
TYQ/TVtPVcL37AdltdQ+mS5ODCt+mWwjjP+iFlxG7Ks9krKFFBi/70SNpMClnF+C
P6Cd1GdFE48+ouQRNw5tWzgHXqHEuD+OtvW27tK9bC4dHIkwIK2yPIkx8I8UiBFz
jTjDttNToFWC2oDAbThHT9C5sevw0ErEzE4yptuSVkKKMOwd5+2NEAzczWJh/0wV
+pwH3tdPKUjAgYQFdAPWFCFBASXRUE02X1YRbh4goy9oKiUweT8ZGoP0XsgJcD5B
eNecSlrSAp3REYYdJK1d2hyjvvo4o+Cbdf1sy8d/zGvoQ/1KKPIvxb6qDgrnvtoY
hd2pLf1P2UihafEHZeSk09kE/F78GOg5u52KHYZT9fc5rDpOYACVq/21deW4TXRe
NN27L8qF6b2WmgnT38QLz/xB/aBDAtnCksyMfnI+ImG2zM9//CQVJA4IfWB2aUbC
/NFDDtwmGMxOikQgjlEBYKkCy8/1jgNYr3Tl9gJBUUNSy2lw2DDcdlvWx3RFMz/m
RvhzT8nEceA8iUSS/8JkptqoQiOARTQJyti4OFAqNFupmgXCXRqf2o1NENuvOfnX
teavtGDozddeOFD8YtR5xMz56IPaqlr/bDatSWcsaJTppUGM5Na4FyE+ioys0NOf
xxjOtDEsImuBgKgIJogCdBlDBnV784628oDa8G/d8TBKb0Uu1zHZWdrCexWLlSa1
cwbZnvgZiMlmBnVDkx7+6OclliebcfJf1mbqYrqXGBghRzll1YPLFOR2KrsZmGVe
dOF0nvuw6CsXs88DbOVAp6pmH40PPWpTkCQsrP+AUNdori6wxOjjx0aOl+z2dktv
UIAJrmJM5AMLbuYH38C6DJXi+6zaFPVsJAgW42moaWpVbURGzX7Fn9Kf5ArEMGYL
kVgRYt8DrdRmQphCPjkKMJTPH+Zvttmh8uqrco0ucePZ8SqiUeKLtjVrA/7oLDyY
UoR9I7vTUtc4iZQdiH7RNmgtiIv7c09jNnZ9l9UNynhRUsHrlAZvn+LNNBimjA8N
fL1NeQE6Ao3B06Eom1vQ2LTXRgcA/C75SjMgdJeOlPEjoGUaAIgI+UPthwwGvlPN
HADasYXHNd5CQxVHZY28b0lWOrqJb1yQxcwZz8LIOXczBDQKCv2zpWTtERxTsJ8L
R93vKvNcVgbabfBuSe3HLT+5qRO27Y3CurT+FQFynCyi0dSYguL71bnYu2s0Qokl
U/U8pjwj4rCv0wQuj7w3Z434mh+2YN2ESEADsZrwgfUgWi3AnYomKWy6QWMXe5Y/
MWMm+6GYes3sLgWKHV5qRf6XSSUdNsAirGZVdxDi9rqxW+ALy8VAVFq3EwACo+66
veKlis1beFu3utz6QuZ3zQSHrOi77+lzAFkx2MiUmQZeQcO1uuTtX/MBArLqP5Lt
txuu91FjQvFLLF160FSH9inYQ7/MmXuFDi/7D1fmp8/ns7hTQk/9iiiQd4u298sq
FteDfI2qsMqsCxG63gLLWSaIln3VtJTl8fbakO4EHpjaGrhFS4ipPeRe0cGilBB5
id1llqKKVgRt31tEf1/Oom5OOYMYDz+TusR9KU5lZbarYfOgSc2P6uQxDK/rzQW7
TWCCZ5gdfhfDg59OaEg9Q4QL02kFTFP6G1h4o87zgQPcgKkJkiR1ch1O3P2/fgSw
0hO5Dk96J/32Gthlq0KdBDtB4KHd/juDgB7tvzxbiJrBA3bqacXLw94DcAr3W38T
YoAMfn0Lpa96/htDG8uXk8AqbXTRN6YCVX2t0ZtgPQuRGpFqk1hZXTJTf/J9ybEO
5OTQV8pHN00I7rWYQIOrL7QLvHk0AXTx/DrQues3rBnxCs2QRwG9Km/8NlLeRMW0
AnQNdUyw4UczxFDj3+d7iZbS06TS2Qmz6eb6OhrckER4ToBrJf/AWWHoNb6fjEKp
qmWgQjHNCdQCBP2NudaWP6VrJzz3oUwc/a6xyzK+58vkWbKEVJeA+YMaxNrqN4rx
8Q+RoHpPUDiNg8swTPDmPA+dFxs6IjCwh0Ws2kB71ocARoYYxV9tPqqgiL5/kSmA
bphqL/AgZHg9iE5vg96Wo39ddRhNuRSMDaGc+X3gDThosEqcyngpZ3TJ15L28z6k
S/VM6BHCFEiTodv8wWzAUrXhAICNeSL8hhF3blR79bYfcj9/ulJBSNdN9uayQnZA
Qgh630GVBwxfIVwqJwvr6UfJga6YgQYsewHqB4thNxUpGXZKZx4shTaMJzxfhIUl
7Ff1l8Kg8XmMgwdfHaWOi2+9uWctAUZ/lRS04jdSDOuHfirLbDAbIgKt8CzG+60A
EmwmqWUeSKImRHYQgcOQOENrPefxsYM1ewFQkzT9U9Mp2ZuMVAFf4GwiQS2Xz4wT
gRvN/AmnEjWrppffeVCXEXwKqNcuAxoTv154grZdcmHkdg1/CRQX6lo8N0m47I9D
8AZolzLNxmXtO68oqIkr+UT5N2LTXv5/nBBUG9aQ1oE+wLmCkzuGL47D9oEufYx4
Z86qcPvZp9KAlr80+fMZxE2ugOH8xCIF9IGTv/o0PMc3rjGccX4tNdQWAZJnVkMF
8YbWIcn5HPLhNjfuS+32mgkY/UjEUZpo8Ki8zYWtqrCHKOudVCHbxXHFfkJvOVgk
37IdvLfd9JpaBpF5KOknKkBLt8PedqB/OKu6YVS2HVpB2H3Xot/FaiLmMVPJUTeE
OzypGh+k6GARqHtn0c86jvN9kyHzclts0EextG8ny0YLYkBVm3CCLaYUX4o6VvQk
bG2DYXmbBLEjR9GQN+X7FeinTZ4TD3tCZdDQAh+FdmtODgR7VNBPF8Zdh46u2Vk7
dxWoRaVoRpTfHfAkfE5aIeYDGMBMVemz07UnB/ti/mXCqUUvmAv1oWkA69TVQQxE
SYssmDPVw6VlwXHNkFSG/ZRqNfqfUMVVrBewW+VdVu18Db4DZU8DhgSt+X7/azS0
782H7UqLbqY7K69pcWHvR6Avl5EqyjTZ8oGO5CXeSWSmWGpJjDlVfu4Y4WBbVTtc
eSab3cTkiXBMCMKxvXJ9FlgFsAKY2pexHh0/9VS/UWN7VTOOKNyLTiRQ/P4HIy09
kwdFR+At2HfRe6cpTtbArJrnrLytnLGbMNWtkjAWG1me3kF7djEw+2dpctDD4WBl
NQfCv4Gw1a8b2t11rVKmbfYfkLzziv6q+qgOzP+HXfktygPtLa0VwlyZiefh1kOk
/6rrTv61Y6c13ubybmxtZLta5+6ksGwuhfmPBPl26c4V/AjQY1RecSmEgK2vhCXu
39IwaPHaSDDBsH36gTTuymxZZ+H1vivG79HdtvHVo7VgM86z61EUerjhGT2ToaTe
M0Kf5ZXuYBzqMfUk73iVCsbaBSUcJMDyBSUso6RulJ8i9MDEZPZHkfMaueGe0ZPn
8xgWHCs83T5kMWz6nmcyd+b7futGEDU9CSwrzMg0Baq3sqvScjGIS3j0rafV3yaS
W3lzZWQ4hJTZc+8eDvysfVjUafQ8BmFQjA4OisF2sSVjGEXtTTPdgsiOSlhJG0q3
8/A4OgL6X20ZtuYiEXALzyD+zs1Grwd4C6gIId7ClXfZFdSigfUaTCCHizm3GS/W
BvbCMpL0XHHFYo3w/bF/aRXXl5RGFB2VOwsHJcL7RZppy2pYHF1LOHokn1gE/k+w
7xZhFhQzmRDSwBal/3cRzFtLYlfVCRn4oInJ8hoODFfSTU3WXdR1kizNE5KB/4Qj
MutEgXq6bg8jA6ytjzshYYjqmUWhDbMZ6o5pYB7xYJau3FjhqTQj/S/lhUxwVbha
PfAKBLpA0Oou3rd7sX1Pqav1qviNX87um8K3SEV5SIbBrDdcybxtzjSL2z50fCj/
qwpFAv5hh3vvv9+s1x517scs4dD4ye0PGmA/PqsNRt3ixW2x97L9qQLzLnL2M0FU
F3yesFTya6HDI8BDNT4/uZCqBdSZxynJ4WxtUBn4/maV4+ZOwjs/u09w71Gs1c9L
M7Kvy5OSnlOhex5sVPKiwjxoufsrLv/Oa3JTaao40+BdnTZMZdm0Kp9+Onfd3ys/
3hLTw+CDxZnztENUpKlVr7YJHdw87gb3qeLDzTfiQjG03QZL25kwoJiZC14Yu4bD
KrYVuqf3uIBEl37Q8C1Yur6e2lEAOXQWN/u/VFHCI94xHg5AssrEh0v/rxSrKzT5
elRUP2C6z+mfmmqKRcp92FlUfVwRI+FVrfVl1F9BnWiCMpEGyGamEbca6TCrwAQ7
34LAMv8LkT5H6iN3q9+SFegXDBlZcG+fZyK23VSW1gJpysC6SiLRh0tQ/7FEC0PN
36LUg2JeIMgMikrD3iXHv5sRUWzJaL1TeY1ylBWszca0SEDW3WNT8vg/Bu9ZVgpq
Ev0mmvjV2iwsOYHffQquZ9l8vSNlwmbvTiDbIdMfhvg9RsrhjyNyw3QFhgw3igRN
MssmDiIJFiaA7kxeddaD5FYhoFeh6tkeGgcbF18eJIL/5+0EEEuqdrkXlwxt+V6z
vW/nRQ9NjFJ7BDSGGU7ReGrClNBRdWqta16cPsWgcH7F8V1QqkuluZzPbXSweqXi
akeRa5RuBrh0qlUAgwbPr5fYHjaHe13/u8WixE2vEN1WbomNmVdDL2HIx/lzWmua
2WlfRc9bPIue+chO+NlVePOnP+N39U5IEIBa7hdssO6vvU148VRyTSWDTyGW7U3X
VWujQkcraj8T3HvfdsgvUecloUWrWYROmURJ9jBOG6DSCyGbVbgZkUDFdaAc7ufP
dvKFCI6PTx977FSTXK5J/hl7DKAtJMZQJj8GgTDhXWVxnX7UXK2gxBfu7sHGjcJ8
2dDjO07iUUBLKLx1XJBBkJx7oEX1syOPyXY/RYHf6sg9mqFEngO/4FJfJF4DLlwC
oNliZUfJxd7Cam+Zi3Db7QMhC79OZbeK3URihtYy5MGWURVBoPC1LEhVZLvmVE/n
uSWKvvGxY9x8v0bC5OdY8oD4mwRwOrZ4/fkPdwXo13BPwf86WIrcHMQFi//nTB+Z
d36ZRfQ0kjUk9a6sBnXwAJVdtRukMEfUqQaYJhY6UqoLv/SqwBVfJ+fqDCsRC17x
4GcV6jhuq5vhBuaew9RtQNDpcuxSMIX8AxGbNQXRhy0raX/QVvHNH+czaWcpvt8d
P0To1pZoIAL75C3dQ8jdl2gSpre6pg/iU9w3AJAg1RgEkOBJyHc9vJ12evhgmSoV
UgHEaGtbPvWdZCWdv4rYn6tE0sRIw49Ql76RaA0gZ939LUJCyLeQlcql+jKcn2vs
VMdbR/5Mv5pWrb9qVbQduM0kvl2xWlB7c+a3yZI4XvW/hq/BZDJo6FBq7iArbOGm
K5V+ppe65NL42/ROh2Ldr7zRy6k/X83uBUvBK4M86SmR3os/M/s0ujrru+o9LDJj
0V6k5gLkWCBTZ5TD+pP0M/AA7FmPKnhEWIqvS4lFmcXxoZSl07Xhi3Q9kPB2hRCB
FTkHSM8XHfUboiCO+n3eGGtxpyaE8ymJK9qKaOlmePI=
`protect END_PROTECTED
