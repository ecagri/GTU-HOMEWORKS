`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1L4cG87UV1pcxjqFVMyVcTNrhDvjcPMyYkTddKObOGC4OEt1bH8V/q7Fw0bmxxb0
3kLQafQYso7ya2cUcRubMTpoS1uoVz+EKAb1wkRe+ABiJMjSfOya8WMwamZc0Zv1
wwJJI3RfAsqJDqet8DzZnG1PVd4VTGkAa8fROZ2MDipZYig+mvNT3D5AmRqlJ0+j
r4Xee6iRynv3RvEydCU3leqhmKpolOxcPYwG+GMYp+Q1VUWKYlni5crsPwVQ2sb9
xgq6QSjtFaG+ltC1I6ufd5MvD0Leeg0pkLapx8w0P7+OAa8H2gpAZJzh/QIJfHWB
BwxZ8iuniVl/YFegerVWqrN6gWu6CB7bUjgXFqtl1kCVUG6WtY5FV7UfqPFlgk3t
Y0mDcp6mBJpPuYBbiScuyN93ugcAgpanT7VvxqYQ0qIfvnu3JiBi1STBAcLIpERf
+d2Kw+fcEQ+BFAneRfYD4IdGKACzvHH/jZkMKOrtYCHzoPNlvhueMQkcFfv74Yri
pG1Skmq0BQurvluzxt37ByFWcbkRbhKl6Mm5fFOy11AUGbImVCawRiea4lWb/Iom
8oS2JCcdmPr7XwbvXlba/Bq3yOasg/EDHt3LGVs+dYYuWkXPkki9zuc4NbTRezX8
qiQQDCH/e0Pom0t9enMdZSWv2tW9+RkgK1Gexw0619FdkAgky9GGNl9unuPtLw2Y
kpqXHNtsQ5qopZEO15nYksH0vnJQj+FoB32zwpUa5jvDPZv/bMC5orpPqIWQRmaz
QJYxCfjCuuM8+N73N6OoNYbUi4ZejFxKPCsD3qbV3jQrLS+SeILln2ED3gAXM2+N
F/Ftd9LS0azf9cvmXCxu9Fzo55W+mXxQcyuGm/mLv3ZdLGevbEPERegMXBsGm2VP
fYcedKJXJGnxGnHi1d8vmFZdPcficFnebyI9UkEtj+zpmKl5irPc9H0iMm7SLbG4
rYjaZiGqTwL74MwiIN6/lmmIeYBUQlzlb9/tZGkLlLsJ6zvEp1ZG0eL70jgGcyD3
fNimNmI0aXs3pOL0Amgy30tKD1sGNRl4HFa+412n3r27vWiBZKbl6Lgmth5afnbA
CQQwefuhDOdrMu+3ZYW+2jWqIATC9deW819o7QDw9/iSg6BHlaTRVrfQKLJM3M/9
cFzIp2VwfUg9CWOXRwMh4LmY4oE593I93mGUIJvB1yrAOCj28wSFelYo5YZgOSmy
NEhLLfdp3YYgoytmvrGf7mAa+7wUNlzfU7cQpqgTpqRiY+GVp2uYoSoZBV38m0tL
1Luke30/D0NAEJdZyOp3iknLdkiuue0/1x0T7VSZiUlMpWk72ByJnPamSIjPISZa
LxFEOJcL9XTQdtvorp1hFER7M0TomsSw94W+oPyt36KrRHO141DKI97zSmv/0UbL
H3YaWW2eVnszvAoTMfYE8T7f+tIfzEThdgmB72I69J7sQPE1odhKxJYC9t5A26Sf
5LdgEKryCHjhEdpi2kpIGR8Q34X0eNVVUrTFLwyUAuCLscO9bCcrqsNKMBK3+MnI
rchgJvk8RsLuu4X0wrdoSSDsxrtQxVbRUtf7Lcg72EzOPIADOkC3/sioWIZExjbc
4LCWMQvL5sJTUX3tqtJlZDo1/M17lF7Oa5mqclHiil2i9g3sGe0z9gnbUOBdNYnw
J6crEu2haWYY4hfqrDVial1hCJJqbI8FLppt4hEVtUQpstE0WwxGgGu3V4ACj1uL
damIYJE8bs2ucAY6XpIG+7a+Sh2vdwYw6/4zq+7SBTts26DPrg1PIqCnMsiOZut0
wut3H57GCSKyD2b0iQ9eLB1tkh/SlwCLw8MqOmtTnGc01ifHyD+Dfiui6LSOe692
UX9JoIT91/m3/mVmeXbIJ+DDsA+4NTXsTG6/2o55lUmY+Kj67+Y+I/xQp4exgA6N
TWhPBVedFgYcQtMWnWTzWH9LTxNWEhD0kR+/0w4RCIPRP81+9YlG7nXm0WN4TF8G
qvRybH3Ac3lXdm00icPgt+j6ioPmGUtbIjxkgMiqIhk4/z8Y35oHlwclF9vWU0fC
OhZ35GxQ9bDJzaVRiTvjA3IWYL4ubFL/WkHXepWHUL/8+Iqnbvv6COlwJ3jx7ZCO
X5NFSvdXJ7XS6YkilIPYXU9/LOTxBdyqXTQxPgOpSi+v03JcH9h8M8gJ5bB4a9hN
KCAXTAehVP75rwaYuh/SP74AGrVd/dpbeusBAew+bbbh46zvSGA+3wWW4ny/p9tW
4IqZQFwm+TIsmnE0eyTr2e8cFe5IxzQ7mj5TwcSJCFgWaGikgzCoSbF+wkAIk8+O
gKseadWcLwYnKwryjfhgs9Sb5Zb+EngGP4ffb5k09C+/+blxUheUA8mJts4nj3EG
8ZKWu3kozCo0jzZsykwReeBXs4vtN7LYgDvrxz6A75RTEukCMjgwsQlsKJsDFdaj
sAbl8FC9/W3Ii23f0LrRfMzAJCOXVdNuI7CvwOfssz1m4TSs3fRshECG58cvD2em
iA2BlOHWRw6eWp+PbgOJgDKjdtKIzvdrJR4pD1EMEEFAQftJzMdxsr3C9fiYoBcG
A0MqqC0ieW+bS6zwrg2LRAevpaSQ5J21PqWGGksp5mM1+yhTkdfuJc4ZnQ+opIsR
NRYeMWRHk3Jxb5S62noDPWqFlkTJb3jn055XQQqFZYp+Mq17a5zW/2MWciqE4o4y
wceGswcF3G4zXShztvpk3hHV6Csilm4qNvjqQX+XPlaZ/o0xPhorvX2MshgDtWC3
hsp7etE0p4RPPzVBFo8Wb+n74Fm1qi9CmYvSEQiz6WZnqC1cHQkFQY33N8eNMo0h
Hxc4Hm6ok8NmDTH11OaceY3+TvIdn45pfl5JMzaGs+1mewXNwp6XTxgn5AsMUM2y
VBA7hYBYv3Ljf4jqqfhMBYuaGWj1UNV8rmxIvCiz3+T3QkuXamDvIohWjUr8rcik
GS+ulBTVKlRO4rmjJI5yQdptEZISlxnVdZRbWZpoZw/TvW5MPXeCFCCuFUWs5SXC
Or7xp3llmK4MoGBa5DweqedSBQCDrD2NZYcIkdiiq2aoxyUk1aNAUlCranSi+YSD
RDwbojCn12VU4LtD1wivJt0KPK52IHrZni01UZoYnrPElYfROWeeu1Ol53CJP+tg
F7wkBvviPesPS3eNhbC9MSDEHoMLTwoqOn9DcvdpBFhdrHP/JtFUdrJDX0gv+2sI
sgQb3anDA4Ixe7RejDTgYFnrHNUGRRZxizSukNurSaKu/p9ihEbqTCG3KDCIWiKE
Rr259uh4hiTxVU/QAyA8oULTtfUhkhpFq1SwWcSkFYFKM7aOL/hfGuXzIsWO/bBU
vC8PKbN5PdX2C8+Ble9mI016iwIjFARjQiw5pzEfl9kkKKm88OgUdE9invQ5frCP
DFzEoQNAHks4GsubwK73yMLa+FctjRM9uJ12xF7khyYdwKDoXFPYi1s+r7dq/Oye
PHGkP9Yh8uw7+fL/Y0m7m1trp39oxm3KiHEfXJai/I4OiyHv4sYw/iz/MgC0HtJq
jxoT7sGvpcHKsLSML5mikeJfsGH9R+ZCg+Rs/uf90tQhD7LAwvp9VbbvNSxE0u7F
75EkI3dRzjUsQ7NwYCGngIEoUd/Y7sW/b3IWLYmIHbZfSvih/199U0iFPI1k6O24
ZLK/9qMtatzdgv1GZcSIJZzFa+QeAgq6h7EpWTTx0REtquX0tyqi3ZRA0xe3U72B
kc2ZqdRfnKzCMjDVsuuaAyCbHW4UvnSTnIx2XLEhR9bPSopzNRf9oleQc/aM4W2k
RAkYZGuK/Ql7gFrkh4aXuvre7SU6JSMbG6FCVhlVDYDZgjKFFHmc0UlzOy8FMvn7
y2glbv/3od0URbr0ntRrqcESPXocabWkeFS5ldqi3bWqkDKA1X7/iEmoLcCfxHW0
3fZid9HlD3IXTYtsdr3lcpL0e1PGlnvy5ExZP/RYc2zrlFuFzXPAsns31Ra83XoW
5Hf4u/citK3+pnZ9TwByMdkwlqNg4HsGTZgPEvkeEzGIPRXvGipckmfzU0zq5YbF
aufw8J/Bqjmgj1mIdNZJGT4BzpjnYkykJ2OcgjfSvNUNOmMT+Alt3uWZgY+Fen6X
DzPklLsf+02UsgQBGzIKCacB7PBzJoHSOlZke9vli36OVD/ywm6DvuCzvSuR4vvS
CX3aLuVfemgli2BjQLmeWnZ5a+pKn6kx1Ufg1cQUdv3kBcyNYr//2X7QqeW3JGKB
wjLOZKrRoxqTfI97rtY22MFTeiPcdsNoBJnoGEBT+KzxOyh5CPFrycOnV5yW3T2F
rF7atvWygs+mYYjRMg4AAY5g5u92bo1aJ1U8rNhERmpT5gx1dWUpKNyzd0KNYoTa
pR/KKqHhqVTRRtIGSkCEXUmX73anKQeiCVKz2eoBRn0NqpeUCoay6oyKXsbkPRWL
zk6LXQe5kELxtqypYu/XKWEu9cqj3FecNdFlGUzp0UWHRsAaJEhNBfUJhnUS6yY2
67UTKQ94Q/Q+4CWD3ZBxCAtSvnwJMyB7kEy7cXuAYSLh5gwzM7jJmq7pJn+4LIpk
cCngX8ZoS4/XPMxOo5tNVX4cWXzIUCFHPZkTYF8iJEvCc1cZ15YnYW62TM9CJMY3
sNEUgaoQFYcucDJG/FUCHSZtUxyO678HmHF6Nx6tfqmZWn6flX2KWhl2FjvpsAhk
Imowk0TtOklxUYYi6hY8fRVFi5gBTmGzyQ12gh3FFLyWxQoyiJHbTDmt+zkajGgd
jTcVY6eor5je1TxT7pGu4U9m1rXDY1XBoRQSuG9oqrzhl2zy9ns8JK+cToiLK5jT
WQmvRrcZRKGghqiZVTho9v7rrdRZxSPYExRnP+dfGrjdf5vJn66gJ7HJ5b4j6hoZ
atzkXAu4wH9JZzg76j1NtRo/phOeDPNn0qdlwQA4qWESOJy4V972Du9z5cRd1T0z
yIvjk0aJ02USQpDhcuU/kj79x9BZzuzIZBaAa06DH53gLDNTkGGIqEpBuxrZkHHX
Vx3+QXZvaliisYUY2A0oNvvnqnfh/rJ1zr48xVphVCamYM0SYVsFbRBnhzCR6Oad
5kiv2ugfvf5v6hc2Rz5fFgrjVvIUdHaIK90PGxmHBXQ8A6mYYc0ndHFEt8miUL1c
gLB5gBl4RmT6yEU7ylJg5If1UXhLX5aQVfMTr8TlB1+8kfjApEIggP53WgP1lM4C
qo0psmoR4JK7OJ/4Ijc6KhQXbYiSA4pB2Yfe+T0ND7AZjtLrD16ld8g3d4bWG00m
FSqvQ8fqP9fUO8+nsSmG7OdxKp5vbi8noPYPh8y6muyz3kRJiDi9/Rmr2tUNsMET
Ih7n0nrMAuMmWja7fWAPoWilUUWPjUu2LsBC1ycvS3viH0484IvGTQPRPLbINMBj
Y5HUM0wymtUV02MQrtZ8LnKugytIfh2yLeLUqm7/KuUnw7ijpkKyRkWKqxXT7e7D
R16TmIyu09yBegcbm/sGvIHnXliKgN50C/2CQMiuD/2VLcOPg8yOPRCkARs7GUok
bpQHqcG0+oZHwfka9Dq6CpQBaN/CpeR4ts15o9keXsXMMyqkGXDkG+46wOeWM36n
QBNL/VU2IGkgF8Y7lC5QmsfDrIRaVIL8gUmAQNgjDs2GF+kW3UzaHAB4G/o/PcdP
wqlgs0He7XfbNsQBnOtebZdHd0YaR7HhtXRQXaQQi3S7Ka2INus3Sd0sLWda58t8
bWP5u78C6sroQGPGnNYrdSZJg7x1mGWs/o9V4t9PRLwyhTAbWw0ulJMSNcaeu5eV
Tu7YzWaC9uMR+6+If2rhrHJZq5eGEbTkq6SwtdLbp1E8xKORJ/7wr94QZkiakfLW
OMX8V8ylZgbCOYo7YtTZJyLUyk/rT3UWg75ukxJubQb/8HYm02G1ks7jNF3jg+W/
+Tp3U5N76HtWKMenuekFsJ0ZeeSjjSRsrsF9B84Eql/Bitz8dkeWfjZ+TLgBBdyV
GoJr44yTaIcATo5NZkYdCSiCLYKFEmmG9lxahT62lIo3k/l/xgiBu5XsEDWSVCy5
frTrfuw802E7ZFLDnBv4LjXQ9EfH/37rXnEpC7DqYw9MQiTtvunve+JNQNlKqvCT
kpLJcti7DEV6Hu7NCQGGGPydUZATM0fRWoPmds/o1M70+L+5Zt7UGJb5B7Q92sgZ
d8Is40OkdFax1Dr4fkpeyR5xgrdjLtL5Qhrwjp5lXKtgJFFRbJyZtnxJPBO76DPe
IpcYSs1Yiav1XbbZoSWj6VTja2xOZc0J43P7lbij1NPhK2YFsFPE2dO6V59GD+iI
B1zaVyczWs0hOwCbu+bhH28waxB4OAtHuQA003/MFPCbvM3ia3yR5QrtvHhL8M7j
lHwqnC5wq4jQW/Mrq2g7lmD+50bEhO2gAGcJULUWmiYga0y8DU/I36F1wDzjA5j7
SXlqyXXkGvjALleAtiu30Y9JHSa7Wjo4FvQNdHSmKdn4PpHLLk4OcFEzV3qZQtaM
52hqWQ3eD5UTyX0ufJ6QK7iX46y9M6kd89KXhP/zGhlHVcPThzOMsJi1Q/qkl7Ii
N4XJfID6Dg/7+dNBhMya4GHtESIHtvI2X6qzN0ok69tHngLcK1ZETd6/kP0M2Q95
5yDJWNDRnMmv3Bcc0vu5RTn0vms2K3Ib4Ga8/mhvsX3FYpCFJWJMWL4as9tGta2e
AyPAmS7ogjGGLzobNBmreA7aeuxf6+mrkCUJXusg6ggEtX+mF6zt8gYbfi7MwaNa
gQ1yno3HJ3FNPkrKO3Hm4AEFGR7S2Y6Ot3dF78OBjiSRrTWfscN1umIBKlqceBpT
8M0cfdbLqgfwgZju/4SlW9sgVEjQEtZTTiM8tIWumImGLSy4rxdxQZGVbbvrHXIj
7+mwVX1VD41oa7kh+YYs66VIMLZueCtdUjw3+C7jQjjyY450PuWZYX02WCOPGgzA
R1C265GOE9rU6IGldKDO3q5Z0t8smZypbi2LwtyIBZ/xdTuaUuNFGjZgZ2rRJePL
F+6wjA4UtrnxnaHADBoP5nhDnIoK1Tb0BR0UUMujjQ1/KdKV9jHFxhDeY+f50X1T
UGYCM6MBa/6YvPZw2SI1o3Ri/JhaneY52BPZj/+vidhGw0ceRsbrrNKVSKZL/CHS
4mkdZe3TxoV5lAY62eoqt8lzZJoaJX35GN8VKc0yCiTn1H+O1xDcxtLjCdTQ0qt4
Eu1yF8OrkSlRxUASoAdSSorowc3q04FTqMWF0CrP8sLnLXTKcFdpxhsFbjmi7XUb
H2KDPBlc+YAS/3dCEbf+X0N+gBoXD9k2B2PBQHvJq5qL+h7nyHbMCdhHMyhmeu9Q
VinsbG50vkgVk8lcdBHtBrwpOxPAQAIb2o5GXRIUy32M2p7wo0UsEV/p0hB0PLWl
K4ovpIvwvC8jVvmugwOpMaY2luZb6EpLvKhYMDm5sPgUJHnTiQuGGSgwb9p9UGVI
BXkfmY1fu/+bmCF4pUv1+NpeycewEoeA5Uj3wUMJAcHhMbo4qg/sGJNn+/SvKa6N
iaoVKeAjHiDpTAKkqbH6G8vUsFrRqZvAfxSPBuUa7nwG6r4VMxrRYJ4xmyhiA9ht
RwYdML2YecFMCCrM1CrFyQ00sD8A3pmZV7wbVuZZCXiePx468Fdvv4AWkuB9yaUu
oKJK8Y7aV4DHjaH0vKl/UFoaFCYORNo3Mmk5fQ3Eyp/L2c+c0bz0aJINDpMf7jnb
vNXJ1zfYrfoqJq/X3P4dP/RFH/53J83ky/snTBJN6VYAAdyrCowgC2JFiUTT7qsu
D/Vs6w5t7wNopFktkDly1A1OIAk19b0bkAhXe9Ti3pOMoXnS074YLpEhVPAarH+j
zfKXv3W8nH4loWjmha80YzZGJ7WPOO8EsM6pD+gzYHOxG5lKJNtXw4iR68jIspQs
31bDFviOjp1zXbSWjhsNggMgrrWzYUnqJW+hMAO8l1bzenZDXOzfWj1HGJpXit9N
CNGWbumBZmO2KF66WMBUcmyoRHqTg4MV7CxOOy/eyoLPhqlIhKWRT6ifUl42fxY6
5aV88KOEK0JYUMmb6dOD+d1qbttgJkNqv65q2klvDnekeJRozpzbo7BDjJ9Nej5r
jyCKOjNFYPYkyLonwx65Y5G6Qrh3EqQ7DmqXu4rc2KyNiHwTLEVvR/8XSY8mRbBI
fB9pVJNwj0eYkBYtBI3yZK7RzTFfhFIQcdHFIwdC+0a6ez2IuBv9R3vdZm4ThhAS
jtNs5A+3yB+1d5KYq5FdxHgfDo1YTnEFdCxTOOJoFXaQCsSD1ujO39CiS6kIt3FV
n9Uhe7tPQhxiunldpPBYvU1c4biTQ53imsVGggvdYz/PutZk1D9aSAvwxVJf1a1K
eXur/co63T7C9jLUz2TuS06h23jl5mzu1EsvhfprtVgILHSgmdpffpitIzeoB+N8
7h7gqjfQIh101eYQ2TTizE3pfKDZAaxlHaCDeiHJFoQrdwLdPpq0uZm3NAxXKu6G
yQOfntbRsiVwpkpbvd6dKUNJLAmluMmsIajFSnme1ulUS5R5L8EFD6PpOpHCP85e
/Gxinu4oX1R4QcyJrII0gLtj8AxZAmd8VrqSWY5OtI279On8mGjvSxOvmDiECcD1
mfPZfvTis7JpRfPpwNu8sUCvtXOi887NLcgKGXOPQ9Du61bLhsFPma1gZTsbk6aS
EFgq57YMmaANE5ja4wXqO1l6HExs+UElo6jn5naP/SVXlIN7IobPINW1FRtF5wq2
CyYHjehAl3BY7k8I+oB7e10c9GRdrVj8a5HbSb2YWuzvDwI8yt6rYifiiBtWSIf7
p7p1ydjIqT/BSrjlT5x34AYISrt3LTWKn5zI2lj0yb2dIXXeAvoVhenP50wAGT9b
pdBoPFdaM4FnGeke3lrhntT/f2A+IQwD7HAdtFXKVx/GJ25YhEi7JkEZMbEmEHjU
Cb51YxXXLo27zYHEjAvbPM291QJP+waj5ihPY/Yn73pH5dm6fTtZAJljsNSKUjpf
WRDnClsriT6n7Ig3MXR/bsrSswQ3yZS1TwaVuPxjGUTXcc4mqPCT3wSi41vgdhEg
ADLujl/55r2v8QloAN2KRelpqtoLgqQtXe/an0AumHql9R2J7TE0GInrnt5SAR7i
rXRcBUbzDIMMx4gUqI8xPjxiSsadD0yDDO5kIeO8fy1LXg2mylfVLh/FDMniky85
lJqy52hzA3UVA75FdC3JtK9PXWmtpe+/ZIdaYRyYqAi+Yfs76LP6WAxoy7qzIz/k
DVc03J9Lu5Hkpwg/dpCI1mOoRMaujDVQc09jAcMEpPiPPJt8puBb+nR5KV8zhdCk
bUrFAqTonpDHqpwsHlwL9REwKDXKSbcrTSXlmBXKTVhRpysGL+QIxP5mY6VeT60D
0m+hV9fEJRJWY6TiEm5jeH6feMJgYBZ3c1n7+iwpSgMCOaxL4RfxN2cfLNScrVvZ
wefGAX7grdOmcAuZIrIY7IuYmzD1jSGBU9kf1IYAAsstode9X5YKWQ7t61egXVjl
5GTp0sAPqt7d1WqSJjFDlHFW5hqQ+zYCG1eiJkT70l9TOrZ/7vuJeg+4fxOELar8
x6H1JNNxFfNm6xHruikUuEdQsFOoOwakJXhmNBG83kfh+hfNTNstomOTGH06qVTM
lfV+OZmLkNFrIL2miDl2xX7igdoLNMmwzqMi9KK/Wee7kpXkw76+Le6OBcNqTjwl
KThNIDgqMSFlhV22PY3let9XuX5Ru3lKhqR5vDeWo3OrR4EXfjdT2SIOtC/dJvcT
oRueQTYXPpXay6sxPBEX/gTBCiXcIrKaB4OsieUbmZoFXeJwDFx++PrtTth/sNy3
+ChGVUL2WwPtHFfCmmoyvCCUwizCAQojUYFs3FD92egDC9yrbj8CKt85Bvmbj48p
OeY87a2E2z7cQHfMJq1aeOoPFAdLTFRrJAMwwmE+O8b/CGL6IMrq/o/HGvIYO9jK
64kba+/9ZWp33Uc7rVs81UisETwQ5DJxxYTlkO2nEjqco6u2xJ3dOWgjlkHrbEyR
vk1sd0Q8TTMFf/Q9WQ7KHMOBC6MOhl2j8qQIrDrRNNz/XY6hVohHqjtf0eNMalSi
BVc3f+EEx9mL/WdI4tsjPB1FCwQOrTf7pVUba+7JnhiamXKcPM54Rqbx8cUCJ5RJ
LzuFiJKDhLkXo87kcS4w3AJUwz+JzI0MIAytQEZByOMgUZ2TBmGHg9tWo46FQlSI
hKKNF/YrqOxct0WNTEpfsfLBiLT010IrPsqTK4zay20eMYwAN/TExm0bdYCLHtbR
pdVQD5qdiYNqwVakpU3U3VLEDbKmhstLjxdJEaSbq1pRFSYGt0d2RMeCEvNBePk/
rwQHpH+BeLqMagyaQyHPh1hbkr73EZ4LLTtpMHg2fQwrtZfVEj38jmW2SxKvDXWv
6uJrnyHZmBMwFjS3vzB4A5i9XiqflMHT2xRX5DQRvDzoNWWy74IPtfNIftn/KXsa
WuJ4EiU/V5JzTLfMedNjj4+pF/GRJ5CEVKZ4SqriLYl1E24YJEkQYWl+fASGdSNm
tnvZIeb/oA3/19GecTAoWEryRM1A3J2vziUIcKsnCzkGMB+VDCb1IrPruEWQnRNN
cFjKMHshx+7+2L0tVqxev2n5naC6eMXlTnjWq8UO5tP6VWgje/cfxPqq/3MR6kzb
0YSajr/c/3PwIjb2lSwLDgoGWXonmECHAHaRTssuEr9akGdvBY62QAR93MSSopPt
tYuP5bYveLsVpe+HjoZW9wbmA4AK6Jm1HpMOqdRhZqq41NThi0sC1prsH4/2Mz/T
fyY60/RhTVf3PYToBgeJ+mhrPhdaRnzuJJvtq43vluheJbphKWfZaxGLDSuJvwm3
BiET7oZ0/4HutBnVJe4R+oXscp6IGUlCQesBDiCSJcHbKLL58VCMREhbdRzAuxXU
klk1OV89rY+j/Xqbc4WZ0/OT087r6Zb3TIBcCHXKJjHJitp/tnBy9ttpz67NYRHy
hCUPlMx/2qEENTo2AIoL7i4fwbOtgqOZs4J3lkvxlzn/RF4ZzFHH9sL/hKfa94Tx
E5YHR6wux60GJy4rVX3GtEtR72lVPaWYmxGKqTlzsta9DFdB8Ak2XIkGJEjlTsgs
QX/LBDOEbXyJDLyE72r3/BnX3r8y7nl4P8Uw/kWr2LxTqQDdvpTK+kokL150hYBI
nncoskweAwHSsYXltLlI6YL4StxjmLxAo48Q/FKvwf6Jim2YYKayY02kplX3S+WH
s2XxvMOpyuUIqtnv3TQ+TnCmOgiGR/zLNBmbGW7Gj00QQG3/pe6RIAXuxXMuFAhU
sSFpPVBwv0+sKDDzuJ78r13QW9IDTYnJrwYhJXokrtoAU8xkYDBXpe/9xYWtVr4p
6tN5hUD6g8PsX6BZPb8nkLGKpt5bSBUgd7p1JplkKt6pqx4qKEYlAD3QYh8CPEIn
IIVVbaNSeXu89Jwn7KJcUIBLtDSkKxIIzqYcvy5XDA829CWO7mZbDaTihN7fgXky
/iFutM0KMgJcmTbVVCc8OgN4OWA/COnLU5uTS9pDvF1YFHzHljqe6U1bGD00Fai3
b8AeVLPKCTZPp4mu+ntae2iCBPscACwe9GR9GA5FXXzbOMgyPcftmU+S1PO8HbLM
R5zJdlLxMfL4tKgHG3/JrWXmPdjUbWYZWfirr5V9zcg5/pbiBOjnhkXL+yYNIKSB
jOcl+Hg0zTV92P+cRI0E3p1ohKZbRd98O/xti5uEF326yACz+RXoSj9cI1B7zK2K
OKljn5Ve9PJL48Hcu0u8d6jHHZ4HQpxLGGnxidTmv9XV7UCYHeoc/nQWRQeepEqx
KfdaN5C2uKpFQGyeyN42fR1HHV0v362L1JpgkntSqb1BSFEJ2LRtGORjFmNGTnG0
fOyRJuLC1Tk6E1zkyGAEBUhAiUpfJ7/Jcu2AGlcvJzx25Fl91K9SRQze5kh/xVej
YiGiJic4qKr60XsMHB2aBLB0n61wkBe6xBvtAdSMdLeTAcUOzAUP0tkiYnavnuxd
RbvHX0fyozhXI/jLcz4E40twVniqjNS/Rc5V3xKDMoKShZwTr8/Oh53on9+AycTD
mSjrgE9WlXIm6J69Cxk91remNuAPKIN6+YdKkI62VqRxpcMOiVzVS9tfnPfiE6mo
Dev33xFrUH+Bs4kJnYDf9MQoZOYgT5oO2AYhLvnt5B7PEBBgcLd/Q+QU0qA/MXMn
aRo3JwWxzmF2NMw23lkVJE/Gyxt5dEen2A9s9yAjN1k88Ale5vqvaoKiagM6q9Tu
e/HPPbi8fLpGJiG8rI6SIydwOFlE5xzMesOcPZYpR3nBe/ZEcsrS4zj7QmTgWSFd
fwk/lPD0OIQwczR7xr+JcVUYQueqpJgY8lv2YfklsFLFO1IDo3Nd7Z8VicIvS5uX
FTufGnTBUxhPShf6PgRMscqZgPv6mQCF+H4LEPgatYLM5r2tu/2LXH1RCSMDMJFt
3iIFwSV0rKEQ6r2U1InOkIJp9XWGDtJ/prC6l6sP+aRK5PkSl1i2T/MZey5BVlt5
JnjoH6pqMQsniG1kNEOLZd1ZzLRDXNY2m66gGKh04A7qj0399Mlk2hXtfz5lYNL/
hN9LH+mSyM8F3e85fknSsgLqIo+lgzNNHNwOBFqLjyEvm8bFnMPsQf/bzLLipsxE
7dKSETBAVCs/cHLXn6PYG/TO1xLYLIdO2p+RHT4kneYivmNtynmQrAOyMfN0RYED
ijl6lBlEvkqBLby3WXhm1R152FYW+raZuw+Rmdg7svk96MiCZaQFT3hy1saAdOa0
Sc/eYQa5/AalebwRQND3SPn5Ht2sqiRnHJVKJlDW0RsnPK0VLvbsjXO6gh21sVpL
6bA6q+00MMmMYUjBHHgihvct4/yJqqNAtoANMmNH8PUdJQ/xFnV3qz0zcXoIi/LU
n0KLP3DOX1+XTKDitr9sUoqiyrX9LoMBbf3zfvfXu5x35sVFwXSpObAu3hh6XYkx
xnbZCD6UrUVFfinPQCdYq7mcz8o3yO6REqghd/Ro4FrgmZJgV6FRAElpo8s79yBa
E7+smTxxdHFazD+vcvkNrIGVE0SMf7JZKNzJnYh7ZT0zt/GM+TOHvNsHhR53Amjs
TXohY4PKeY4OCD21q5ERuZPfr3asrAa7Oi+FHdrGY6MczTVN4eAFcQzw/tiheYgj
/572cY+EpUL6u2qQ6pHkWYQhPQfuljPhNwBtdFy+SecaaTkCs6nG13KlxXefNRkx
KU/1R8wNRpk4eNsdzb3FnpzrmRZO6iazXHiELp0gGnutQt59lxmClVBO1renm7bz
rfS2j6BN0Kp5L3bN11yDEXbDwDHMq2kzNBAccu39ARw/pYK+Q/ao/l4xrJJ9CrLF
kjsDSFfir3YjTBvNVvNs/MGX/mkvuc3FN9AJ3M6Ys1dT/tGc6JrCEwoyS5Gy6L4f
hJRRfAo8fX+DCev0hiKWsXj/6Rd6jjxZX8kHRd+hjKGwZWnpF0Pqa5hyakhycliD
yHGCJ9RkWEgTC5FjmCol1JXJirLq4P7TghLYO9xHtCOGvb6q1Bhoil86f+8dzkFk
jKu0+wOoOljCQNgkdPFToWemyhWkONEQbrr/Gbx74s/wpxsakEVCW2mmEX/J6Uf6
FlaeABT4RyltTaOAO0rXhjy8jgymgFiATFAMPHOBpbxLR+KyKniY1cacfx/ex9B3
WdNfSZK5bju6+n9DSdLJrxY2zWz8kZnlCMidu8p0cAkDdXQUHEtAPg5azkySplBp
dp7jLm4+ioQx5KI9TaBb3RjQOAMfk44EJ0RwnbDTOtpOwqe3t7KS9kGN367trhqz
WT4fJ60ZZNezM/MZptaTM7XBDjbSyshuEiJK7uIt5YbbJBNWQdhOy3ZYkwirDMEF
PzykhJf1LIjy4rNbnrciE7/5hayiojn0UR6patKAeTV7wmNjelptBgbPLlodVnLC
7uDM3AFnho8K8o0mAg5Q9ytWuS3awX9pcUq59HYJqZDbPqLNY2IQg4yhuAyXy9cT
a8I0X2jqTXvkkDK1wseSMM9uKIQ6uBnTqAqyN7Up7yaPqvYarzYpcYrXp/h4YSnX
ijGbjn9Nbqb7/2op4wuov5zV1ZgampourBLBlLtw2nmi85aHiuppb8M+osOltoMr
sgPjB8v3VsG2DXXbzHMVK9sXm7kDXWJ620al1WSTdvCSw4hDqDajoL2uuuMxWyvJ
nJUWfeUIIWGcgQJPIKDSiN4gCJTu926z5hsgYSCxLb/DU2INo7CoevPDSzCx9bFF
1wDB/v/e2m93JMcX0RDJUo7D+aILF0tJOmLdnLS0n9Uy2WqvlL2Tk3TKX/v90WS3
eHKc3yV0aLPV36yF4dN4QMxtV/l6Qxa227zbzpg9McSxeglgGFFoTkbCeh/eYUwF
QHDrc/Z+prKyMNAzLtE3cF1qz70yPcjpSMn4Gwp/bOJUSMWRzl7ZLiyaAuLxQlkr
ead9F4+cbCAVpzrDZ8qRwNtwxgrVk4ipcVmMvgLi4Q0CnofnAqwml/9/dsbDfXwA
Jz8BeClVWSOZ93uSdCVSNYqckGhZxqJCmLGD6JoAlRGwnupbNewObunV0qLozNYv
i38G+GVBNgsNpcy6a4aKeFYcd2Z29sqL91U9AdYzptBgGtddRSnjLcwuTOxR4KFg
fsuVf/rKaiTNpXXlOGGDfM31bNAouizTtWIO6i9vTidfO/fYWPOef1e67/HDtgmX
TdCtttdrOUrmdwYiSb64Buo45iC51GXRwMHfq86pSunRdHFIn09tZ/9V9p9Mk8Ny
xaHO+7bqMuCJXJDdDFF76oHRM9g3Oac9z0wxNRsUgDSiRWWqnXY6CGtOwKZPON5+
r/SB8E66iV6vfIMxyIRJJImc3bEC67Oa8CnBoETSEYW0lhEjnHjCsuqx8wxPg2MI
5C5kPXHfxy66qmGngphDO6WYMFZtSVzQg4hcZOycMQ9X7bSySMe9YQTkuGKa9g/0
yxDW5HG2CFK40O10lhzKdt4CMjAWzyEVACfycgy7VYW+FYZrU2kCStTJ+iLazmRW
zTIT/SrHRhS6DTDUQogVXvZlpNsFfermGJkoRw5CYrYcefNuAcj1aOgmM9J3AsaX
xjGjyw/1h+Af2H/kbnT0jKwX/9fyCHTalgLNQMbH2vtcmcC3a2NpArMGgjTFgxLU
QzYyuFNbIlhExiSeUTm3Qvcistk8W5ab7x9VtTl9p+6/lJNSOq7u6vJR9ukY93pC
MB4NxiS9QOVln/Ty0cTi9lHKfY5sW0VcMcQxnDlypIrDL4MxNHcmDRPRvCJ1sDAe
n8aAsx+G1qDvWxmfUlqB8c7edtHw0Ln42reBelSpbkjiH7ZbNFbEuuHrQkjVUevK
0dMxvJnKKKxlnlHP3u8ts9i6pUzFGYPhUo7a9w2Epb+c35zhfnJF8OtWO/KZ6z+i
3pZLb7MdIGO4OzYuPIIYHOFyGKgnd2rZWN5Ht0z4tZhDfLu4RQSRMcA9t6K/c2uN
ymzlRRuEeAxOB7ivHJbINytxiYt5xLH6Ez73HjzeqJiJDCfzrH403APXilELE7yc
eOer8/swF8TAcxJB+4LVgowGKIw2Hc90kTXsarUFYQHaCauDxckmLW7gNUTFelhI
GcUJGQHPNYK7x25SSbYRfwigkdmUjTDiU6mP2/5D4ALKtBX8KMmOhA5+Ol6Us4EK
TzDvCgyZk/3PoxbRRAtVEFf9GbavEGlmo3WJSNE1gW7bFb+UPunU3yhV2RrFAlXF
ZuY9ZInxsKJ8iF3VdrUHopRJNLESEDO3hoQ51ISB/yKfbLOsxdSz3/x++eUavVzs
fDgPMxAZMwKSbZzuB0JIL3HPGCgAX6pkQD6C9UEQVphyjIV0zTxq8C8Ssyp9ybin
T0Ddp4Sx2mVRPSgO7cVzaYk+et734q3qHSjDNlaC/wt+2cXv/GN6gKE5M+q4++9X
SPMSkmP2jK6A4LO0PFpVXuJoJQtyGelOV2fPyCr/n21NWpoX7/sLpKktGG6vt44+
kyxvJT2WRSeMkCt8u68dcuUjx+51O2MmARsIT+7UK2uJNTEHGmSWWrv5YDElMUe4
VVoC9c7jIufY6GVbaEfOUs2yNJaCpHaWmBo1txHkElYzl1WxWOFBsf5WP1CHYx+x
dKMRE8379sTMRiKXAdxbmRLYJeCSrZExnOrRtw0KTzPzRC31+d44ev+0UCgO7ouD
djAZ/xE/TeZfFjBgNlCE7CoXonybV5KM1TdaMe8dJLCwJJJC0wojz5YrJFn4uMp2
DEC/I5syLQKoCQjoiTxafxKlfelUgIrkMh6srTHMzniiIh/qt+aGQ9OvVCFR3UmN
ize/3RZaRWp82iFfVy3bkZQRtooXqQw/5x5gqSCFcSYLZz9JSqZrQugw3LgAl3cI
dSzuSA/dYRnbIXBGSindu21RpjGQ2Wq0lUSlrRJtVNH2M4StgPsqeh4g7794uJHg
vEjmnqNlFWA8u4+p2BOrXT+AMyr/CRdg8SbBHeG8T9vKCeUnR/DQcviDJQkaCd/I
JFlZQAW7lzmD4PH4vQOGQ6kkepI4Zd1lAWRb8SVz3WCMyi98vxscT/r/8puBs7q8
bpBWEufK02WFwBeSk7OR9qqtCC4u6N5viMS2bh4ZiOXKXKygl4jmP4MS3eWuajSo
mRq9apx+pIRGGTZMOZCXqt2Jme3JYoHMj0ZIYz7EKsn9ezzVLyphP2VXgmoZbX7X
qNHhLLl+ROxP0LzVHfk3fTDvljkN9zTKpIl3UwCjZ1UEc9WW2xqTGrHz4bcGT708
19LWvezv36IxvOR0aL6RlhpCr85Zq8MuGHM8PhlIzuSZi9M7DqA48060SfJq2+Cf
krvU81IjnD0qlsIXlDLUf9ziEwWxDbU9Zt3XYmZcxKvyU26ZusWchGRX2/ucjJmJ
RlWHOs5twRVwjjJHKv6Bdma6Dz1P35x8B7vTwJHYn86f4XDRuC5Wz0LgIOM757wd
QZ0aPGeASiexqEr1uk5ub3agiXOQ6JdVffo5zjJvv3y5ZnXnsxpukR6psTmw+mxX
ZhwHPKRFACHVOJ/U5nGB8eTkGCK7Nc+l6X8YBD58broXhF7FWw3u3qntzWFSc+fn
3Zn5qQjGdvm32wHqGZJAA7yhipFKaB7srqVGhnRFlgz1o5bbwtp8wUsmkY3+BLZ9
K1/LyYSCY5y6uPn1fUBHkonbR+xXfvnf7v0xOxgWSX7hg8wSHflGuYLVfDZd1I35
qr1qwNzapge2H/Hyj1aerr7Ac8dJcPfBgK2AV+rRfkzkhytadqcmoQygkuBwf1rM
VxEDmHYSPfeDNwwGaUHMLwq0Dt148eSF6uiacLJla6AJ3M/iW6NLR5VlTAZvXzkL
NjOxx1j+sn1yPIhNhjG1gOq1QutA3gkacRs5xhLPFchHC9RIJbQNMICMfrW1ee9J
jHY2tqIgtC3Rirn3nl/NyeDDikEejf++LVMzVYsraoZzdqlliShtR5ePAbNtXK99
uwYEDSWpYE1QxpzU++yWQ/S5rohjAkBM3p13GrDg5xtF1Vk/dJTRw7ZX+QbYZnXU
/EAR3tO640wL9F9n+yf63wMbrxBTrfLEeBEC4zZuIuqrrfOhYZjmo6xLVdmnFk+S
WvYlWmUHRe69gCFMzabbZ0hs1gn8AbzCUK03bSPkWq4lt0tV2x3gTlc+jRo5Qhmk
sB7vSjbAYEiMJ95TME54pJzRquYWi95XzlrJPtc8VGmp1n6vE0c4N7VbyAagHsed
0vTVxxuCb+dQuteIoKZJDvqnrYzFo2ueLTXIpLjVfNQE+iEp08RRJzXMDfSyyocF
Llads9Urx4bNtRTctHuPhja2ef2s36OfoOjqrMG5LCoVIy5Kf7FDdmaVKsrF8REn
BBNquFUNIk0nUb0erNpeJKiGMtGh9nx7oPNcBBRlzetWYdJUecqb8YZsNdMaYQvx
1tZsLwaSjmvWss4SZ2ZyT8AIa6CTQd0U72yLXKFyEK4Vt6yQfYA/noBXcHM6/ExJ
wN55rOIl9K4+wi6GaEDzLRbxs/Sf9yFY80mTt6Y8SBovrJtb3Uwjp3qoEMWFDzFx
3kZSkkyqSGcTW7ZBQ1y1ar62btjAUzLufcmAHV42iyD3ROxhTHKeevHLKVeV7ICn
USQag39y38UOUU0u0c9AYOggF+dQ6j38wga03KLWDFokUxHEJr5v3xsKCPvOvm/w
cNbW4fjgH00AClDKALHq10jptTW4i6aVFhhXgQNj0+nl7SsWJvoaxbPBoEuYkQ4j
x/BE6NKuhDGMgm2NWNIEOvIIiNRMwLfrf8ojBErVhmGsK0mYW2tAUajDSkXgSIkV
09fr8AUXUr4FMjDN7y6iFFRtrxx8mQqh+2IWJaIa0naVrp7Uvmk6zKF9XAMm3Oak
wanCh3g9/ekienhGJl7ABE4XZu63MKEGp89Sm6rxZmqLn0f4j1yGuJDksZb6SWlR
EvblItlzbPRKVRiJOiLUYd8qHd6kaeKRsdbyBIJ2KPEtlOP8KbloedoQs/R8LpqC
s9Lh4mt/KVULxfEu7vl0YfSyJvzwiJveh/zADkxUP2nXvP80j3ukT+hvPp4Ngqyt
A2qeLF7lW68zzMoOor9qwtGbhTuuROPuFyUPwHzBL+5BPWUHbWOxxrPn2fKNknqk
dPrAAd1TmRJoapZbnBtJE6cnrGmRh58Djc0kVNGuOm9r6n38Yu4teugL/hV1teUA
zB7fH8jyjDLK6OaeKfqOlvwFrXrQBO/B3hSzLL7nKlYyUsHWuowS2Z51d8Fwzjzm
H44Uem+KmqJt6jYrP9KR5EEwcJ1fiBK3/vKXUpADlZZzxre8HxsOsJY60Rn6PMNb
7uRXv5VlBRWWxbrr+RDUXU3oPLDYoLgDZfjOPK8RwSb70avZWPl70QuU2nVIyJOX
RNK2FsLG6Cye8FoXUoeI6v1cRHBuUq5hkIRcaJHcexcVg2l2GN4IuImxbi5Np6HZ
PHqKwIoBU7MIDsbJ+4BtstAru2imSW6jZImvZpY9t55Qtnt/HLuMFx0gx9JSdJtM
ZAePNUANhAOupuY0HXmAE49HqcIJn8tPqfzgLejwhlzCYu3keGu2+QVbFUT15PT/
SjKkTGalMKoaXZheqp12MtWvsL0Z/udVxqC+adXbTozuQfZX/geLqPxsUg7VRzT8
crcom134LTS9wpZOFR71nV6TA69cOAoOujqRz5phoHqGhBUuGar7AVSoyIWNiKkX
Bz1efNzSfDuqgypzEquXY8c3ZIX/LIqjXg+liZM1486d6BNuj5ih/u8SliPlTYpM
YR9tkzg4Y6lI9erZH2/xnP+i8EcTg1nDX7skh1TjbZpLKBl5r7TTLXsv0AIdHRy1
xX9EhKQOFU8Nh37alPmNiIOFHYxrmkyAYGAiHFZKPQgJVXfu/6wXMw1yA2xx/IDL
VOYIJ2F1FxEpTt6uYvVks/y8pIqQSgiz3mWs6mTkvOf17AAjNtynn1lc2c3ES2Gy
nVgxwOCLNn1RKdfx3b7iRfdjLfoN7zz9VJG+YXsxE70vlhHU9ft3zJuIbG4oolJb
Ol/NjQhFQhH2zJmncaaWa/czwACL7SoVHpAJqsmAS1QbwjEPc4bpHcVWB1A++TL8
Qg3rL/MNh1j2rMSIHpXD3RcCaPvIw1upkWuLGsHv4Wu2z0b0yOWQ8Bab0Zcza9Q2
+DYlThLJ0HRFw7lCLBzDG3Il7q3b2L287V1Ydy973tSC5PRusGaeGZ9bdTXQeDWB
rY38m9r7JD5ZXy8IbwE9YM5jBhfuMS+QYk+bJlxcFgqaPRvrcgjnUBOkK40gv8yb
/FwxoeuSMIEBbnL+mTRE5KmdKJaDR846yn8EI9fIAXw4X+aUkikJbjmf6C/yCsih
mc8aDoqdAc+Md96g46crekuwykIVwXGR7PYFmo7V8AOlVYNoyGgsUArUNyloMGEJ
W9WM8lDQiMsXmnnrK4coYJ1p2q6OOV5gWjoTXt6sgtqEiExvzkaafWQPRXcHikuE
35zou2lF+hNSxyCpImfvxg2Px5T+CGvz6IljKgfaqxuIGjVa0nLOeOK2ZCYyag4j
H6C9X+qHZ8XT5bnnuz1bwknk6SnvzJUcXFWuI1fqcLAuxzRr9ssrbhpsRo8DVUTq
R/V5pyok0/EVS5dX4x5qOxBiLis97BVY0vLGc/GAD7haQfgaVaD3pOTjfSbxKPYG
2VJAHYb5JGqwebz8oCPjfNbVny9vjzVYmOL6lL6B2ig86tbQPhWpDe2ru28e8xUc
JjsEzf+CdfIeVldfY8fxPASAlV/W92HD0wlFuis3oXu47kYy1cDEXy8LIypba2zk
z7OYO1EuIHxWEVdK31ooDNxTuUB/UwjWXP/Xcz/qta3+6qN7kSNQkodq2KA1jx7o
CHowysWXHvYJPxaZt8eDdOwraczwKKH6vJFJYob8+sMUZ1LxeGP5Lw9EaLuIhVUr
tY39YZJKrDdNLMc9RvEb9SirfUvMd+ou+uwPYlDOGhxYztmZZ6vKLYb8vOLC/VCa
IT9jMyycFtRlTGAQP5AbFDKlgHfVIYDhd38LIFcqQrsdxHunWa/52Nf/P8VJP7y1
ccpPwoilVKoWxHUCJRm3KPgYA0/IebZOeROrHvxinVxwiTReAYcSOkufsc1G6rAg
oON9SEhkNafgjyV0I85slIyAYx2o4AZBAWOXxqc/BnksC+L4XLsMs5jNhsLLWg/f
0jJ3JjGTzjkY33+SxzCXd50lYGi+I9OKafBO8zE2IWUI1yDsv5pE3TXDDaV++/8z
O3aXmUmXlFWU79oRWVHpax/heKEZab+ZUk5l8zzCT58TcvRqqh9FtOwyjIoI46rn
ISeyDMHO2ss1j9ZgNnrYWIW1ivB1ooZHnBHumBQC31fLgNW2C3L0L2++ueQIAHi8
yWTs4ZY437BlEEcVj/FeOSfcBJOvILQrhpxBCEzHb6m63W4TTbUwXsyxJFymYB5C
zNuBysm4gcxa7mmbGrYwoWPxkKUitBbFr2LTfzF7RSPNxhkOpV6XDrqwx2QN7FUH
1y6OuiyGZLFsnzFCBF1iH9mtkfFWzLQiYQgQ7/Nd5yJugOQLY9RQ+1VPEsyX43E4
VdFrcS9fdj6yeYR4B5NEwfb9mF2VEpLcrxOlxQ0oj90T0+YiHocJ6uMxq0Fiqh2J
l1BrFyt4EyT0nD6LwKs/kRGEbkXN2x+YllYunpeVcNQ2UeBnujR6LqPtuIfVHTfl
KoeAxuSC/L3gz8y7IVSY5RJx2yF08InsImEsJOYFtg/RPazuW56yLMmSVFEQiLI7
G3TjfhyLUK9pztusK8JRJVYZ/T6KhNEXJkxLyPsAu559XCZMnRnLWYYuZ6SdL9Zk
DHWlQ069REWlhbbi3CieJj6mYLu/POFJtUFn61otfWGZRPPu4SsAc5e26aR4SwiW
fe4VpkZ5G7Ftw8SZJjRU7+1mpKISkYj+fP/mmFLE4hZbCbjh0T2CmWdXsY8hAe3F
NnKEwqaVEgT87AIcaB1n/ZkvdL7gH0PpoQaurONwFAXZ2JF2050qpESKoF8aCBBD
AlSVBkGjWIvfM9zPFtbVt9S/dRegoFX8r+OUCrpre0uazICt24I0dp4McxyfyMGZ
i8+WurwPrufyi+y8/MV7RBRkQfMLVMae6aANWhwSEA3cFumyudj0+yovXUbmMxBn
U/YCOlhisclIlo8yeQx1w6uK2fmS4oCX/EwMXjARDDYeifL0KmfEAWKB9MWkDRHK
7qTSECc9/XKi53e4K1+CVwmMDT8O2zjVkrjsjqVeIgwbIILQw6uqQkMr3E5KvNvQ
hykj5QZBckflBdG4cajJATGrq1LxMZJzA7Fp6aBLdv8X5/zVxwloKtqg17Fdrvro
G67tsnGrJ75Oj9TWaVxgTANy0MQu0IXwTbTizP9nOfu9eH/7ozXRm1yM9lJoDxpw
U8Ma5KYOaO0uDuvp7xfcSieOHArVQafNBSsLhgLGyJGjiuKnMq4vuG+mDqEF5FKe
GZHTEMdDQTmtfU5gX5cgdsQP2R5o5okTkXTQOZA11TDM5E//k+3/5TpATjYaBU4a
Xt8sdageORiOE1FOdqrHdg2FgXI+e/8oCS9/T8SHJRC+XRb/VW+WZrEv8PDoWJkO
hqc0KCOO0DGYyp9TQvXCvojNxMKWulIidbGCO8YfVuMJeJTONZXINy1nH6W3xF3X
lmFcMTc42fKgMC+wWMFtFBCsAJ9HcIJvx9dnRNoQZvntbqbrbQhhv7441ffhtf4e
ca7L1TJ3K/JoSIqfPyBJmr/vZxVZ47BmxBnqpvOChcz8M+gaXM6Nfu73n78fhobj
uMW5C0blBZ8NoF+Z4VJ78lbwzU7TunrgT/7nHjUJpjOtlS4k9DaQ2E1YMlyuXXq0
3KT5fneSoDRMvKV2/HwOazKRkzI4QK5i9i751axfOd8ZemyFpUhfe2TVx3FDgnIe
/06FMfBTT7r+LElJUgwpiJB+0H7OkA9Cty7YLzkbwBDJc01XuGtUorUDA+24HYNC
2XYSzpuLV3hmY1ImoQUt9v7PcAApVCyBmISo/khaS08S/RlxYvmhDKejpgT3VZuQ
j/NZsUkKQwyfY5ShhMWT3BAPgIJdm+hv7/aQOpoB/HXwqC1zpqQiH62Eh7ljIrs0
/11C5owldFTmYjo5DRe/lZshqXZ1ZLq5PxqAECRueNl224kfrPiulky4c6+HOEbO
IUrJsE8xjFUPvWKduVbXHPrp+HmkrRXqj0W05pXP2Wjm0JQHy1i5rvaEJ7spylaV
kyqSJOxrPBjUroSdqICMLTP9I+Cr/STh3IV34ppMKdosqzOxM9cKHjnGemGr5uHn
IPLZUezdyCnqkDhH27xTZCEgQDE/FVTQGkzlypQrQzOh1XaRZDzCR4dRNFE5Nqoi
kdkNmiOuIi9wcNLKO3xnPG/vuDrswTxsVP/7RJIFnZfCkYCUN2o9SspFijGmrqqS
/Wy+CnqtVhv0ZbKTamF6RRC1WKcgArpgMEhCSDOSQ35qZQfFi0TufYjxHZaQgRJz
8i1F8NBaL95aB/RkhgpRI56D2P/wbaKIDnsgeolvj6Z8yWXntI0wyQgcYmyoL9ag
zznN2LDJoXy5zSV3ksqTekHzH74rfQeh0glgT4mePAzg94q1LT9KqEI0tMGx8MJc
xAi8h41Z3kFnmzxxRyK4fKlJggTkruXyob/h6Y47sz7ydxUm8jc6+CMMMEfp7SXv
rlPRWC3xy0LA6RkNuE2Wl/A9nyt7gT3BeBM2fNB9vEENskt3ZrBSPuakAv5kudRD
RsdCiDMXhm7tks23Nyr8QTqyAdIinjZvwsEE3nBpcwIa/Csk3uddfs0emGothiX4
9YJ06pt/2CLwlHDxWEZ8Pc64Tytu/Ln6YXHMBbKxv5l22RZX5pox8EBFZLPZAkPi
8bG3FoRdjzE45Z6qtgEbCVyA8Yn8qGquqZ6A3XGm1IVJ6j+yoYjY32zWz0zCD6Yf
xTmvOt1INZe84rOaA5wwUT+d3r2lXSShkT3kwYEpKll5cMBkVXEro9qfKCJTemIp
zzL+yAg5YufEldhsJgSMVzgN8zAtXRAMjP2v1iW8C7IPF6SbaH7yPoJuSsB4/LAI
MAQL6TIcN8CUcq+iofr9P0R6RCinEx20sq1FpKtfQabolgiJlD7Q+Yu1thyarYCN
ehElrAywjm60Dd+/H5B/JFRcjAuxqIo6ZfqzA20kALvGrMiuTV00jz4O2RLuIoU4
JIYwNHSvKXdHrs+JC5hE6fjfRCZPMoKtl79xFIgJklLEkUzu81obtFrGlDUughyU
zEUyfyz0O+0nvBXyebsQYptbbsuL4gh1yvQHuXk8HXSfElD41pPSKBQfKTSco69H
20OgYPgEXjIxsV7PVh5HpcaEJchjObuFmqLlU28tPsLwYC+O5CTh5a5gx7AjkY/t
r5X4JqqIrNFvpeED2S3to4+x0OAB4m7g2qejK/onglGmMe42RQFCNnfe33Ob4LS/
6vAEZQ3So0l+OaR9Z4M7pTN1KL7K+kyUEbwbeJo+ScofIb083/s4bE/N6Enc3/JM
vpwgWdA4s42g+VrQhnkPBv4r3pO/8yPcQqYzX+h80YLt8pdPSLuAYslv+B3mlIYm
aGv7Q0MXQ9Y97YsX49gzltOeMuJjAQk7osiKAsORcy/KUbe1S+ACg2dyXqWIRSVS
mkXL7wcQK2elXxDDdJhh4vCWcyPC0OMhGHaoHj7XkEq3K2ddFWkWPCWqIuQX+med
0SCpwxl6KTbVkRrl4dv9f+BT8vU6Pmu80IxMNMdAKKQt1fGoyX6id+qRJoy7M6FS
7zEPiWjIDl8/TPS4SdmKzw1nbcx5SaCWi0P83NwCjC47vHwIjcG5WhqsSUE2+rvS
1dN2gCh89rxnm1FpWsuOvsvJoxps5CDE5a+bY6VoCfABv0NDaw/1ipcFJRSPfoE9
Lh05z2s6KjlL2w1mM2jm+CQhdd8FtAJnoCW9jDrgXz5TmDcEoOhhzW4lyRqe3ngz
A9VbxrpReCPtOD8TSTzfLz1otoeZ+yJ68uB0n0YkdaBmMoUTeDF2bB90MLO2QGSm
Lym98dngLu5ZN5XJuKUigI9GIFyliaJgPRGtpsU1FPfR6nwlxGL71pa3tM2ZpXcZ
7CWNkypYa72pBTnefDGD22JcW5sDwVe0M6B2nJSBx+lUd4PH3tW1ucFci7htZ7//
edq/PsZsSiWFgRTsS9o+fY0AskwlfdMwq7oWZb7mEKgJg4U1aa7WNN2+z4aplnxk
jVqkjNH0bM9mDS3TTLSB8GwZO89Blmg4mSXZDSOnAcVbO17T93b3InnMEd26WZTA
dg4cbtPu4Bf4yF0qpVGn0q6ISC9j7xbDR1FTvXGHFqweAuZI+vB7Re2zzmTHzT24
7rQqz3pfJNoP0R6UOpAkPXsA69CDXt3eMSDBasX8qIHFCchPYrOjeUHXHy41Sjdz
QEgfPFV3nrci9QPz1UbdQwLvu+wIMyGgIE87DgGJ7vKR4k3tbb1to95lpdMhitZv
6tVGQPpMf1BQcYRF35NbsN1+U8ty2TvyxsZkbHrVT7rPtlfKGKxwQZ+tClltbcXh
sTY7MRIJ6dbFGZlTv9w5DAusehadAYb1rh3n5cN+LqHBMMmjXWBCGph71wDUlSpb
ZLZslKXEybtZSDSoGu9mVGXWGb82jEmANdbQ/O6fzX5BEmZZUr/jbzm4UuoQ9Yij
XVuyWQTYBZTYjDQNORBgj/jCet5Beek+SNUcxlck/JgWNOKaCqDPkCO//kXaHyut
w5bzDB/c9NQSW8lB+EGKYyZrP3RpFDP915jsBVHKnq+YvPqLeL7aCPhJ8BUMDYff
A7girRNiYmSnBPduoosnrqXor2GIDG5PnVvuegZVhFcnQB+rcr+2g4lxcujLjzMf
lR4ngUDinibRcmW8RGOuxmG0//Fh24P9xAICxK9lLEoPls6nvH7Yl+Pmqc/OJ2im
Ztq4ApNCHMcggOOsW6LK27hofoM2/Hjosqp3Z38ECWmnONV+4wVw7m034krMQmDP
ZYugNWJmHKiPHjEr+i/bO/Lxwxbc/hVAcUhSYxiMmoC+JMkZMBz5Aq90+wZSlqwp
00WVl3jT2TK+h+JeAWeKajtM8Ba4bSGHxiYON3b2MvIQ6kF6YvJ43uh/g9oHloOt
XZXDwbNgAit1I4jQSUTpySx1pBPDfeodZNBUiBKoaS1fWe/Dh5feMPhNh6hxB9KX
DOWNrRe9sD7/LboVmH6ah9fcj6igNEL9DbmVr7h02Mitvi9rhIWwxNp9w765ICgX
ZjUS18K3yKVHtCdp5y8wyq0eIKawkK9sFy7zY/RLcUCHZ9wdbhiX6+JFjM7olkEp
jym/NqK2dTUyo+HBs9ORMW9VIOhYqkZ0U95Mb2MLISidfp0wkipT3REb0PCsN18d
A65fQ1yLw/71xno0efU11lngmx+sI2RxcL0ImtHNCpII0hWYXbp86I2Q7Vaio0+y
ujPpAiFcNv8nMJNRvaIb9EgeWn2a231z5vFM3FTQ3NKVMfIGxmhBrI2Cn1qx861s
eE5a7es4F5DMI0WMX8f3JiuFSSyi7J6sONGglt+vpVssG/6dwI8KNVb6IEeQD1Iu
yC0JXbhSgprsCs51KwmqfeTmtzSJhSSFhWsZ2S2HucmT5yj493xJ6WtC9noPatH9
o8ekO2RSPg7qTsSqYGYRIvbWsT23yXldMNpY4N1JLrOHw+ZLytiM4grr28CufBvA
XEfaaNEg4rdslJnzoT8n5gUjkFDcnPBKMMycgbH2Ub96caaNs7QMkGlq+9weOm/8
ENB2BuqaYRexQG0os+cCs5e5qMexecvH7MM62WwrYZj57ptqoCz6gZJCILnvYuX7
859nikrLLvfb1RRIjHgkokWIoH/x7CGor6lPNrtd7vg1oSM+jotaG4TlIwgKmrdO
3h1C9U6kHYQq7h6lrdCGv8DjqgvLyNtFBlLbLTVO+9VHMirmZyUCrvXeIzlQaVZm
7Q/RAOxNIUBp4gwZ3sk9h39ukpvtyJrJBvd9AobCFr1a61pXJx4L9eT7astkNGMw
5ZPu0eFE+WwNTN9fhrXvCTfTiW4mGX3me6TDQBOxOl8RNJpAadHBGCUmc2oUjSGH
Ei6XnRYXtyVvTVKD3Q26OUMKiTNTiY5mcZPrVRpef685ol5LF30mIGbIW48CjRN4
qXoKrqXfMOpZpCkvOBOn0xR8KkBvv70eFFKfRDgNiIoD6m2cYkjxbcXBCVDTjTGv
w/mVfe8OK3VVVTKqfv508cg8TUZEC2qRg7gapLJ0qDImLFwhJWwVtMqpfDbeGoNz
gVgwIZET+dVp18Z+A7VEmziz3TGYiR5z9MtSp19BLiy5HUKzZuqNSpQNr17MAdgJ
SNS6mktONszPhrDkhhv1WBzGpekkxxam4wvWRjG9xA7bZRBaHxAVT4DBkOisDNDk
8FaPmPqijafX2mvxjP62kYMqGewf7hqiIQWN8h51WHB0DoImiY/fD3ZAka3Itptn
i78I2XkDiUzHhBLJCuuc+GXBj1EOJhBF2ZocCOcHQTKQs6z6h9f+iXcTu6RWzT12
wRXSX4+Vwy+7Q2i1S9xOGNRrUjo3UbSJak37zK7X1lSqHSzAZbXJeQLsdhNdwjQm
NP+IEYVPe/xZNRCtShEVxmNuw6tQpXB0ofas+Tmmtp3NtZJ4oD5cMEBm5sXuKF8k
HaId32OMS6W1Q3YsjjLvmnSWk7R4rkSwT6VQdBEN+6j6+H/xiCKpNvR8Yoaxfmxl
PpdhoGXO9SIYTltrmtWYIc63oTxndie/zpTSk1ggxDdMI6tca6lEwyctOh2d/ZaW
sRcGv+RW9q54muNDM1fO7JPTRveQzJlTLYSYZ4NFq8mJ8Pk5cUT+9JAn4ZklN/hm
YNkfg6gd2scbSTXbzbsHiYREvvtCqI7tzoZeWqSCd9wmYGpMKdgsss9jjuqW0VOo
3+aHYTAsAt59UK2gcQbeECAkjWUCYVUjaUKSMcHLE/6MIqp8Jer0xg6ZwTE8VF1x
dQHthqB2CIKBeOG7hs416JuQUscu/H4VRe7fbTkUhNx5n7Sqi3zDF2YHYs2kNWCl
W8oVcU/eZtGbbZSD2FEr63KqB5W+aXoeCpNMPndVeWubP7nOdRXRf6JNujtWjaIr
5Mz17C8F16s9JoEJJSNQK6U3iSXWPTbAKTN9kpX5Lse3mhCdsD1g+lySj8nXFqPY
dwG/syxhJ2H/Sl6vEkg+YDRE93fFJcwiUO0Vnrzv2AnFcfTBrbAPESKzXkyvg1PK
CmaHj8T0p74YST2OQyVglstalzbKWB4GajTjya3p8jnH1BCxgmfrHfVeFDPUkXDq
2ibsl/K0ryyCvkcoWldTeptB3Nfka8ociSwnVFbpto4+9edVZkPimIVlXs4rtOar
F/Ybjx9ZhLzqiJ2HXRSVAKOdPzSxjSomAWGDaHnzPmt/7iiQtyUFaS2Tbnu8VH3u
Qnkci+R9sQtmXX+4mjLk46TSgrdMlU31Hll+cQP6e8n/H+MRFDE5k6qu6Vd6l2/d
OcVr9I7eAN0TEEkv/nhQfkwziQNNDCXgrCnTWpWM0ST5nG7yVvHsr1UpZ7cOxeVs
Yr58lutHrSHwu/2WmALexuI72WKvyP3URS9FbfUMH9WLvwGxABD4dsKr7mMJi9HY
EbrwmWvfTeG95Vr6Pq5PTe3sb3nbJaViM8rnZVPI2tJGfRJ5CpcXqP/pHHqAJdYT
Xf7J/yMbdwUeF8lI79FeSlf3lYZXmifKlK8Tv+nXc+X/7gRkULgaUSPV4OIcvIwp
uk36+CCrEiOQBwq+T8Ie5wjbHXdD2Yyv76MuWS/bZZd/TAfGWDXEALWtO4mgagAl
5+5OsQKjuVvWZKlI3SEDwvLPpi/FkdGWype4doma2q/+gj2OtpkbwaWpKAUSLx4B
NCO/o83mv33LR7L4ijpJFnKKRiGRfYyRzRCTrzPhh4K5BXxlqgikLRO+ftrD09EY
PqwVdYzTEz4sh++IZoLcMJANA/zg814/cnboo2GHymQxGinSEqUk+Om6+5C9VdHX
lY+2nN+bAyYHOfoynejQNoVLVyAwKXMlR6pUjX3yFtPLxT1mgYdQXR50K7eo5vk7
95PYUgMbdmTtyB3U8UAXNLByFvkmv111S1GABvdg3M+a6Jvl5RHwa6Gg/P6R1UAC
hu1tSX+3QmLtyeqkYMLkhZauGT5PjOFgdmiC89hXIS5ovthHCp8RGhAklWGgSjOj
ixRJ4e8VSCW8r+bOdQ50WD6aTT2lmDwzqFUH9s3vhHB3OnWbjcQesdr4T2+knGQV
P+l1GfQpn2BAUHJYfoagl/alxnAVx/jW9UDm2/q2AQ4oTkMm0ZzEswFL5U/S5vuN
N/A6ji8mkAxCpmCKgTUnrMw9wdBFFS5fmFxDqtVj+25FZ4A/57wZvIuhlUwFpd1Y
79XMHvit85/olkddGSGNS8QHDSoKgHklsKOHUJRBHbw80mNOSGJIZOVEBj56uIqy
F9LkhINMmCos/Ajlb5vIHlen6pMDEeiOg3x2qrI5+uqX6qmSEd3GFZQPK+bDHzzq
9mWVBPNzu1i3+k9ZxtNP5+vXyy0ZGcdNOq1jsX6n4L4M6uBTb4eEFA4R/FrgOsby
TsU4Vaq0RDh/D5pNabqOvo167BrWwGIOiAaOv2DRc0ZGmgWq/nix8oiWsJFzCGtW
D2HQBMDOSc9W2B1ziKocGWMLD2M+aX1PwQlZqaZV5r8DiSwY4kA+CzdGsBF9dzFs
BguCPdGConb9croZuYxuJDg2RLoPAkCAQ+pIb4LoknYb/Q0U2Z5W2Pg/f1BUncyy
pRz4aK/rcdlRQDS4ykpp2+ty0rD7Vg9EGoSlXpZL4vsy38wrxk8tNzj9apb/yKpD
aMdqcAkVjVLPmxmLPquKpP1NlrFcgRNkigyur1QYirAKqNgLUh1fsVTY3ZkhTgmS
Jv0XL4kqgthJKlVyKeFfn2J4YBtv94TpFMF+Tl/CqH92Fw2ilhUNDpJfXorb/EN6
/RChOACUNlLIErE6FpA3luI1JAV5LnaGzDwQqzh2p1HmVmJKncx+/m8HToLyFH9o
GygO6mdzLJ3KHgd0WPdPtshZN8pJXgJcj8emtPTWTcc3qokblCpdCyAtqNqPq8sG
MUhiLp/xTLa4pG5jLl2dSjZHnq5W321OIWOySMHfM7RjKmZ6Tfa9sZM13vsRNIWB
q3kvh/4ej63ysygaztQy/71x25X9S2kgk2aAsxMTOIP7uCV1FRQP/zhsAjLO9P6/
BjJZXqgrGD57D+U2RxkVd/b4sgSR/l0uTK5UJ1jqlEpyv0d15R4Wsv6k6l+09Ryv
UtpCuVbz5W5a5A6RHfSKHKL2JrasVsEiW69JI7hsYL/FhWugKb7WNQHPkCmfcey3
1aATS3WufoGeffJuTonEYbqhHfnU4abRpefd8L/qYwhI715u9nmvyQV3Xp8hnfPC
K5RDXP8WmXmk5Yeo6rpGS6CDaQdfYRJWlvtlKRh1Muh5JyxWCCgbZgTGLTxQuAOi
JkRAuAecD2pLIbJUSsKnYG2wZCRDk+LXDPOdu+8WCOnwHy9uXVw+QNmY9T/HAvcm
EsuCXF15KzCRCU0gVKkfBUnjTyvStpOappY58JTa2BxPNsJ2bSug9QLE56UFh629
Xazi3lLcSYtxaQuJHlL9V5uBL1GRpmyMT9gzK8WkBH7vAyjEacd64OEXP9BNVdxh
06BoAZg65mdyRN3a/EMCb6SUTEuQvLRwS5I3ofndzgzyM0/JRn+p3FvBtlJCe3az
jqkeGp1ZT0VEwn1KefR/WHYQ1IxIBAb/29M/dQWnbeP2vL0UZp1mOQ7856T1DgAl
0eq/iCzuuBGovuz7BHEyGct1pamaFm9dO3T2lplp9HJhb/fDLw569jNhp2+gcGGh
wzHAAMGtb/VajSANBm14Ew7nse1xJr6CNfpWf9yZAXTnHxXySk3nV1lwiBOEwgFs
qYTzRQuh+aS9ejrs1D2W6rQdRgcQZT14vxdeV1i5d2oDlZBUxS931yKxycVnx3h9
8HrXmzYVY/Yhq30+UAHylgWuYdiq4rywMzMEvIJc3HgRkw8lfOFbRsNy9KQ2IRpL
/WzY5pGxhyHomKz+Xt/eemQr8Nuk8aqZLoBc3xUzkqrXD9ZsVfkW0Tz4XY13D/da
IUGRc98Ki4A30i2TXy5RhKZ2aBab0miJtFZrcl+1Jr80CMwz+2RG7ZOgnBgjL4Gv
Or5nL1NrfN+s6U+7pY3fu26kxSaWdOPCoVncMFK9XT83VT4TEkIYPrILAseufiZV
eIwRbNHPKgqJiRYFzndSddkwhnf+JHD+RK3EuPaYomFuUJcPH2rUzVULvy9OWZOJ
3LpTXG0dCF1sX61gYDXFf0pZJcOi0awAGutx26rV9xdmFKggZFh6CC/0OykgW/pe
ogw6+G8TDvLqnKvxF5Tgq0FP4NPePDA+VvkSMup2hlT8RivWCMg2uZAiwQCarsrT
bOUnyW/frj4MxaFYew1I9uC/iv9FF2edeeQCVBwaK0q3dT5gFcqt231EQ016gpNR
xeB02zo5XmLbEqRE5VM4MfXOSza/aVuqeqcMB9n1OpujaSa+fcqZubFdsF/P6+RD
jYFOLD0SNLmJL5T90YW2orPZ3ZwAtZ2IgklxXZmypMoBRq8WFiFlSeykAKkhBB8u
WIZd2f+r4lHG7NN6aI2cL/mI5JI391cRZCat8mAAK9ljUmFU0ODX+qgaafB7wY7s
ZwzKhD3QOxhgOQl5S6bk/uctxts0ixvTZ2365KXRPm8LcY2G0E7UaTGJSXHHa9vy
JYwWE7Zm2u8GF6pp2jLHO0XeEwLs8QhgAEovOKAg/JZAzrlnnEknhLNOSdq8Jy0C
tsUcUCGx+yZ5r0YZn5IHk4aRjRu5HAz+yKIoRWrcgxbKHwAdgODr1NJ4xokeUQCq
W4Lkj8FIL2wIkfO8BKy8Pfa2jUknBwFdwG0aUN5p0P5RHf5lDzsVUYfJGDNCMmlV
ICaUX+fpLQC0CmiMVWBt0uvbvSoisCbr0Nvoq3JAoEU/Jzvm9Vv0W9ss5zB+AphW
kcsoeMUtNclQRH6yAM1JBlgYYIaoJ92s0KXsCxBnDgT2zACy961XnAnRw1dEiO7a
J4+vrRJppuBDgjz3PflsVDtKDKm0ayhH+/PrIuSta1afPU5RGh+a7c7ByHK23v/S
apxtPADFvo8FxbtTzp5bd92YFIhrFyvKiYfiiJakJANP7mwVxltEDh49n+3K8ZiF
yx1KANdeApfjKrkKhIbP/RebJVDdvouVW3Py+Mv1GF6d/fmGkTWNPC0y6aLfOEGo
ANfQgh3TyhFh+lPwASTIotDWqgR+gjNouX7fmDKCLMZdhRkusTlU1Oik3zWFEQjQ
RNpJkQHJg7oz8ONKOXJo1ERZrv4846xr/Y2BJy75EA+uXvo+tBoW/Orwo6Cll64P
7QSogIYXH8oJnZLzdKZvkRLQ/rsmfEQ3ZJ6zR/9kACDCBrfrfhXAA5iMn+nTnXL7
27Sfn4RY9IS62Js1gVM3XgPyX34+oCR0f+dhM4Urc5NaI+erNMsOVJzDDQCbltP8
i7m/bzGJlUhia04KskBLgCRg4u8IG5EclIhf8ail1OxFmfY2mP2LwqtPkBi+R16b
jkn2r3jOFVXpomY0Ro6oBb2XWrhnHIqYfQ99GN26a/EevpE5GyVDbWoa9yxwsSa2
rNOKtqIxLUPx0Qxa76CR/LJXmxKVoTLyikm5BLVViE/U90uo0K/Y13dGOdDSHma4
Dzp4zDjgfXlWdxm1sZ5Nwq6Vseh4x8UlsYY3SeP6ixMxKSa+odzd4zmzIMUiMsr3
vOJtuCro03K9dKOIxlsYABlwbY5WV6H4vCS/9Oilk7KOVInP8z0wAnmKwhwhDyBR
mvLk7GBt+CSM6KRa4/35D6ZtM4jwm0LA7srG24sdCCvFCAL3WPQR9y/dBPKW3ESC
LSqoTGKs7VRBqaFhHzFxSdSytd4JThjAcosuYwEgID8U7DWKMm4d54qu3/H3LbGq
mJPTnQDKLh8UVHU/pJoSX97OVpdL4JKymemtIaI1KHzx0pzPfWKkCo89tiPMR8VV
/KLcgoVPPFJi3/Ba0Ep9hmkOvuZtULqqfD9PyYbl/LO2327KROPo4nEdn/Saq9+r
YUIMQtJOGA0hzIgotidbSW7gWXXFPM8Bls98UpedbyABOC5QKihVHdrKfoKdpxpi
LF+7ezH/zbV0cNozCtCKKyXGIYjbWMUy0SuJmWFbNW2Rn4h/alU75wp1sctil7vv
AOCRVq80Bkh0x8FS0lavjIHZRC6jPz5098iW4hOTAIjIye2dXIWHoe6q0rMdT9Fx
+3TTICRknJhSIHCecrRJEIYBg6RJz7bfPTrgoJEEOlGVoMavQr3dc+oW5IyElS2c
mdheJngEGPY/EpWI5dV8QzqYY3kyKwSg958Tux6X3P7B1gqjkZ9XnTDO7NKvnOlD
abGHeQod0qOHK0/0TM58kc71z7rh15qbrEBSCwQAd0IXNOi5uCf3+C88gdOo+e9p
DjTzZ7prDNTiABS/rj7AI9U2OIDAgYOzGlhu/iTKfuRdGjLMSKCR8XPAgeiQ7Bxt
+e2m4XX3zbRWCZlxnarP7qLF+RSN2eV3NB3mJaTi6IkOiq1PUuAEW0VgHVSmX1Ko
RhrqpOelUoXUeQrofMmrroN3L420OZ3VqcSaWhazNQrH9LGH/9UtwYOWdEqUpTOF
O0qElYwKGpFNU+pp1AiJ2svTbHZGzko9mxh5UdWaiqtPWraD8Q0+e0lh6uzk0/2u
mpwzYo2IupgU1PrYELzY4sDDPPaZQw/YGuNz0Ko3mPvdrAJdr6lceLL//TvVHIT6
umG18RM4+P6g4H5JCIjUJv/iLpYe0yHKnHf/QZzFrah/DWdBf76Z/ayAoDcgk7el
qgIxAxGsG2OcLxrWb9a4/PR8l2h4cQQRYWb0DfRyg37xvKzC2PYLebRVLJWiN1ao
ITkguXGeaIFQG0KA5suS9DSosFRAUAS6uh2l1ENnXN52/U5SIoVH+ZM69BGDBPid
vkfFwuUYMmMkNc6u9UhUZ1EMlt/QnTHPhPXh7wa4dyB6toZTCwuHcyRxQ34hH16n
J1S7mw9rWGpFjeKjuMr7fTWvtBO8gJjDOt9eACLQfZooXWS7IOJvYehMKPNlBO1H
b0QqhtV2o7h49BYRmtvXh4jB+sQuljyX1tctJhNy/zzsW7xb53MjtxHrTihCYQoW
9y/FJ3YuvTARgHU/mOQ1PqGYfqupyOXEO8sfLcZR7qNt2bUkKLH1E3FSveKn7pna
IKKRIeqxI/TJsyeHjk2RxjKewYy9XHYPxR8TxMuddVErl1krbyYlAW1VsWeA8zON
mzroSE2sRXFkuNWR08eACSc6wOrO/Eej7N9Jw4eLIgSsI/xUxwZqKRa0Hr2cTjDy
HFL6IyzIgnRvQssSzy2lvITsm2e9mqFsm2dPicugo6u75ySW/YQWGpPZMhHSe4X9
l8NOOPq7oV82G4hbiOww5VqpNHNKSzey7AGAfcSpwG4RP02tI3SJduSsCCL9toXp
Sd7Z3DCI0/wUvqDN6wwkBAnJiKO3taNrOoLZ4yA2XIYiVkl/Gas7EqPjzU/e+sMb
QiLamCR7+C3xcDSsL1eDUeRZc2ozlvX+pF451EuaTG6UwUfWUnMSL3VuhChMdTcn
eqmQXEL16BSc9lLExYGEEKH4Vk4ZYkzmb7H8kCGK2D01W10rph/Wi5nMEX2bb4p7
bag7+ixse0zz+k/BkBGmKRR2+eaisbqZiIoFktx1daPLgeWHcSNEXMwdi1Or/yee
tUZKDni3ilwmEprWKTTLnPxc0Fd5fv61t2UVwP0BHS9MhQ+zXG2qonTJffqNirSw
Ql04Ov2UioBuFVuJxma1VoIne8sCXkZePFUQ0nYpEWNaXIaGiMFwPGapiV5pUnBS
2iU2n5FbuuNS7pqGcapL3A+wZXhjeZq6olmCo4u2iogoLdJUF6dgD15hziwBECxq
Uhs1Vqk6IG0IpVfEbu4xKlYYs1UsJLVLZSkZhxKGSNaUUfh7OaXzqZv4eXJ+1zYq
A3WeTzhQIYG3NXGl6wBVqF5FZvC0lMGMeU1CjrkBZZCE55qmepfyo7fUecyLjq2e
JegUu47OF2YlPp8fe9leDXA/Nayxw10wGsmXE1yqQLYt7umH0b/t6bUrLXsbgsu8
FuhST+c7aTniyeRNivl0G3fEZjGgAUBIe/FgEvSjsNNfEavXkaDQfAzT2nac1m9w
Db6ldKmHo5/cBx1MYARxn9JuuE+1DVvWRxbAkXJph/tgwaAVXbdaeHGKI/yiOw2k
+BW9sulvpjs36+T1Jk0invpjmojmoTjS5Lj0Zn8kkCNLCDik3DXZGuo5ufAG2/Zk
U9ON6m6el0ABzjEZaTyGmw6QicJdvauCjcRyRGLbO7UADUo83fyHuN/M0P1iZtZp
HvxQxQIQUFvRlF+Wtqwhr0Vq/HV2wJxtTk3wr3KxJ1BwAVQ3KUfY3oYZ1O105wAK
fQRCZ2toPseh17uoPqmRvPJLJv235RRblrblHuM95/qquDBuZrC2KhJ1UvEu4uG9
0/VydI9H6qMyiFy+NPgc+vwhW3KeC/+OArI1XaloxqeVk+9wKSQ5jVYqNAPUoAtR
FQ2WzFsezvQSHbFdMV8ftBO5gP2Hiv7g82igNJ88DCCU/p8XSRYQed/eoGSSGYtH
bnQeTXlyACT5ZMrlrAMs3ZtyyUmOMsuMmsIh7tOKw3kO4cQINPP9BHgTL7vSFTnl
cYfCAvYo1/taj+U5nx7SnIRHcCy91v/dypY25Ac2bKUA7RRAPhDCB4B2LS61a6bk
QttDkrt1rRVK4MJ8T3kJDkPo5Os5rz0OccK5Bg7SqvIf/GL4gDqikVAvG9oEh4vm
Uk2uhx1PCgsYHK2+e3pQgO/Deg0ECrN5WaxF5npUcgxUxaTGFRfAsQMQnlrliCuL
4v7/GhXQxuTPXCUBbvPaUcJJTV8bEWEPYRs+nTeYOCymq2Q9j63bS/ADxzl7vmtR
6H1R5A7zc9HtN+VMhXYeIpcuqgLl4C+WmiQlmTgD+4XBKgL9m/EF7KYtsjcJrgRU
hCRqWbatx9GYwbbwZRqEOKE22tygJlwl2N3mX6Q5DZAem/LwrwxqxYL9LXryGRGL
gIQqU/hNryT9q87mhSRi9R6683TgCXwc1XunwUg/eeHglTqnONO2xRPSlFCTzgqj
KfpB5eyVkmSOkdLtB3ZbEoaxvfpg2WuJEHqy7OaTCI1TmfU3dBKXbZzWX2MZwYAZ
m9h25Gtgt6GsCQstsoQI4a29/g2MPja3q9VYrYK6mzaSNP+JlEZoiYRt7KKABdLB
SLmaOXIArEhmd9dNaN/Q01DlvR+wGEXaWphQwqcRQp+N7jKZKP1KqcUdHO1Nphzd
lJrQD5OITeLsOydxcikfxaf2tJugZxiXWzkdKnwHbNYSmKOv66RlS12ocwmHp1JG
HFT/X1SWSI83gTHwKclRox9uypxDPmT570Q/av7Ugs9ZqpaJY+s0xbHgji6P74oG
r4jaIcoIG/EYe9oo9NmXbSIj/NZIjfPHnKTv6eEbLIGWLYpQ44/tbG5ZJVBve0kK
7aRSlq6m7wGZ1ly7zWZYQEumcH/ySe+uj1aHka/6Tqc7tI8l5uRHUd7y52gM9QDS
7ebcyW3da/Mflou6P+dZCrneguvsW1ku281X+7+uktMo9iV0mhdnINP+jLm2cdwM
Z7oi/QWFay1DL+/8h8IRJRSBOf3ohRmHsgPKoZMT6ROVTPOXiKTvnzjVizYNchz3
70sYiLueGIrtrVg42y9QWQu52KcAjFY2cdcNkycmOrdjEl7RWJIiC1YOMlC3yoPo
5boOmtnLZXy/VqQx+dqn61vp9hqsynQgTpIpVgdVJUZsnhpSo/lqLPqeLW/SwfWT
oX33hmNFYGG4jWdDUp7PzVuFOShGcPMzGAISPsSR+gO9UM3JustwzakfJ3yc96Xp
UVCsJrUmgJJ4zwpv4rcdZFSnicIysASGBqZJMj9d61CpHNhOISaCpx++2vLPp59s
RtlUGpHIycHdmNN6YjZRIo1VMCGgZR4JuPoj3j0/18UwdnDZGVM1oBTk65A/aTOQ
ui8W1WGxoGop5hLVXLNiZD9VtGOdb2yMIvk9rKuApY6VgZyoH8ZO9OS5siEuLbmg
qDdyLDALJzbGQd5X2clNPNU5I24WnQAG3TsO/5HelQQiDF5f34wxDJX83GrGuJOa
1hxNt9wGzTaVXAeHsiqgzsJP90CgEIY6b5FYOhoLAv5yLwELIEdM118vJd+ehI+D
sqsAJrch7AAcYRTG4Lw/ZkEI1Xq0BWmdpK4zcArlbvP0lVFV6ctcC5E7NUKVSgxl
T1F6IxHZOU5VeCcrkLHOP+RnIF+ntjhMVQd0PGcIafy0C3s//54M+ierYFWcsH6X
2FAP/qHMlw9hFcICr03xjSTQG4zZEec9kHc7lgXRAAZuXWw37AEvBWn4XQVNbA3s
n/79LRwMhA8/t+yviQv7gmJCWATxyS9D3Wm6JZnmmFdP16v+CwJoK3ropAyZ9kqn
DvBcjzB/kkf4DpPJX1f2j8aQMyCw3Bdzs87zazHic38vpkElDx1zPZyixgEwKKut
kFF9jRrAcZS+iiBpzfquOWQzDYVEqFHDJCWxgAY/NkGKiCKJwdT5LXPKRl0PAchR
WBacY/GDvTiDwXHnvS3RYP6sPOmj6mRBCXrZgunsBDLy28n0SZk/UaMa0FqJBmda
AmBmP4yHh+1V3owXDHPXXywpypBBbsrW5Ngq1Gq436UDj3S+xAHdEbCs7ZSrmUlt
MnqDZKj0WKJP/LUjouT0kWB0czyzsacyR8SfnVkMgDYwY7IFIW9cHSJDAqaA26Bq
HBngWlUEtPAMwRFzPvAkKhSo/g9y1MuA0qOcVyGuWR/xHOl9kxYlHBmm2LD1nlA0
CJFrynQTKAiVxwdSf3YEd2g40RLPOEMXkAkhQovpqd21XQy/gR9121hCp+J1GRGg
rwoVx40yGqZIJ3wgBexLC7PhxrBj3a44HFzYoyoZK2PQ6ZeCH9QstNKhfkxiTdWR
62fRkNXKDuvgU2z+EUtFLS+aFZ4HEwxPf+79OMvdoD3uTP7Rm3ZpvoyY0xyyycgb
WzN0yQN2JqA1zMJ2y/Pq2Ftl1O25o3NaImucL2o0ijHaiTF6B7y+yFnq4J+8v7sv
LC6VNKtVPmVUe4BdTRN4/QdGkawsFk+kVO11hB0rHHcniPTe/e9mmJnpNvNTpe/x
87DRG/U0JmWU8D8y7BOwA9aeHu74vksJv+Q6MBYdZEF5g4ATMvEIpFpZd9f1f07j
`protect END_PROTECTED
