`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sb3HUPtC9uLbHTq9Fn3QIe+a42k571nSTclFAnJqMNi2Yt/C7xGfRt9kq42Q0t7h
kYrydENW+RSt4sBSQh+2wTxfk9Gozk/hHkUBj5pi98ysXlcrh0ZI8jVDHkxDlV0s
oPQsy08Rr2TYZQyYOIZz+LCds2vdF0XwpBrLGA88KwXQqFOayxFyXSsBgADvpbvw
8WXpkUGjpkzDlPGg6FaB3w6fUIgobYpgaHikbfyQ5c55Q5UCElviBwzHSsCXBUpK
N4ijZ7dQPE0lt7Y6cUrMuarwm502Z/Zyq0dmHlGYrIrHp3z7yv+et8VOomCVbKZ2
AbrXlAAeOMJwzG7yrryIgQGwWit++I+MTS+VTXavTFRwkQ36N+qwrpEzASUWxymq
rIKGWbBTEmYbz9MTA5l8GuT4uRyrVzCwiMV4EsnO1kdKysPhJX2nxSmdrkHUiXBS
1FzSEQ12ZCsATKmBTXbwvRuGwtbu76PB7ZrgFGx/6dXD47R9HHaMd/guA1u+3zQ4
elyhfGZpslA790M87jMLOXSu37GGnXOsryIBCfnRZdWFi58F2qRIaDa8ayUUEJdI
KDQUPguPbS3nhBDnCBZT059w3zO0jyWxfyFxACC7jk085acDBczL2aiVu6vXVW17
xj3N16hhPUF02FAMCEkihBefcmK4M9oD2EX4XJN4M8+ORZNFC+7k2ad3JUD9ZsM2
r91DNC/yRvbxWjibRZyvoSck656KvseUxWEfuM4ZVyCUutNqpHnFbKjZyVYzw8W4
8DJYUlb1NSPPitG17qQP1am0si/MpciqX5t+bAws8sugLvYJeBCxqwtYlQgzsWI7
Rjf2sso6AWtksawjnKtqgsrKkoar0ef8qc/iBjXkkAv0ydWlomwjaH3NBRsB4K3T
lMUI2bZTfNFAUJCGO87n9A592DFPis5EN4HLpIonPr0nHUgGv4S4bcSdvgtEcPn3
/2HFKL8bf2+jBnzsEP7F1LCsVJN4sW7s2DRlpjczfHzvvOicZTKtDhY6WcWC5A3C
i3cMHt40e9AX5vACfLb3L0wdhnP3V5bnpoXCc8/yI3h2vNj7kdgN/YWk3ysbiUQp
NxwJ7PqsaqjPk+FVjz1+8+5xwnuPsCr90SmcP+qB8G7W1aCCeUOComTd5EheP06W
yEgxJj0SGTAMwcpZFaSf0fBoywqXKXuKmuqZOAiahB5VY6fxehKU098Pgmst93yu
m4jLa53AnfQeTXWLv6PSWCwUm61/vdT77rfTE8lWfjbOLhjsLtGlcuZJMX7t9hHk
D74j70ftNr4BNhbJJO9JSiV5j/NBp0DaOGzGNl9+PaZwAn/NLsjWiolD2hBT5sg2
F/5zZu6DhBOQlLanzNuJvEHOt5EFxXpJiX/pqYnf7i7CNgfcUs/xR+2Yp+z/Enj/
9ZBdsUipfmpjfA6fMhYB/uS3yOWWMWddvgG85Hj4ESBfbOeNRO28/X1HTym7S7sE
e+DhM2t9M54tIS3TZdji8iBm8waalR5ANYGp8Emh9VjaGAePW+Z2ujw1XbUu5Fav
Bne9wOeYff8mNuAO+yY/hhw0QnE48sbFM24/ZXSnPeJzj4+lzOGaYsdqW59It+KO
hZeG0o9lRvP5ULIvWwjWcihlG/RhL8xBkrYdL/xk4H6xz8obt/Z2oGVrIuLmb9Yx
yRoROTY2pLj9JuiY29Eifc7lJdX0OcjnsOm3lmRocWJ+xIyAhWn3jYxojftqRWVm
uHk4PgqYEXOGCXZ+9GNSea08irhHuRXH3L3nfaAp7WtvEVimvpWHJVVogb7IFsjh
vXUPazsn4YAGUX4X5PwSO/KCvAes1sCqr1f+vVozwx/ed0dAKkMHjJQ2EeAKbEzh
C6eLphcZn88eXQmQnqgMeqCL7JXUf/iW7w7YRGneFgGin9EfdM/zrsMkV7Tq/m5F
3ENc3Et5bCt1BVqUVqYyA2c7vMA1k68+Ywi0sECd929PFHi6UNoWI+xY25asmNcd
mmE87vmNH/WVv4ukhzkxpUsXdwN1Y166CymkBFqvEKsBhs+11xbBScocFf43O91x
er0+5mQcJWJigA0sEp1RyTPm1UmBh0T44szvLZUWFCyUWlyIlxek9ZvuyziET3en
Bk4HdWWY+G23Koz+OuTKLQQL5wwdLAGV3bLOkY6gOWE8bx6N8ktYfG9sAQrpmqQv
WX7sPd3AkTADialbVPDOdTI38yoPf4+28ottOettM/VIMykBkjPTJadePSKs/VWL
9j9eDVoUyjkPbUsOD0/9whAIgnhhYIpTAsBbkhKG8vcOi8VuA1Zl76b4kbygUagF
U5BMBon8kro05M+FZaHgnQIs7hDKF/bVKXF+pr8M/u7qQ/Bf0+SB+emZ5sFFU7lM
bT9BK2reNROWiOgmCH4OMt+TohkdtvN6VkEMNkJz4c0DPko2zKeaSn0oZ4tJd9IL
5AaT3MN2PvfpfTn9GpZqD80mOKoij4fTUsuxiVyLOqhJK++jezynmYwrZLoYvNth
Fn4ZcLEH+RQHhgYzODDr28Vst7E1HaNw1l577/1lHNOLc6++38ZMb2JqaVj+dx4p
/heyn/lcDPZLQ2wfPXgVaMjusd8/Gz3vldble2nkJTW8i2fwiSv4QdiFbQnTs3Vg
XUi2H8pjDaBs+khR8ju5UBSlCjWMEaEMXh1XWEPkjDSfb45Cz7lwe6SisU4fGHxm
vdjvKj8VTkNJnrdzR2Wmj15L20eh2m1nD3RpYNnP0wevRQ5agBBXPOLFPIcEa/3l
hpwNeqCvEFoIxNA1hWJRUmwga3EErhsFSY8Yyc1ZRzCYzPiYC9yDGn3zMr6XF6mZ
CQcP6CsOm7/z2+NoL/w3FVC3RoIzUYi1z9sKntkAAsLcS0UunpI6DIEZc1ynawhC
h4rPm2mQyZhIKhL3l4f1Tatz9UXSmBA9C3hPE/5o7w6RJOZvRqJFyQYzqhVloJcd
nJvijcwoasGLk4SKkCnpkePp/G+A4RStN8v7roEy9UoZF8BF/5dlOU6Zt8GaJecK
E2TrAydvZhFcQY7e7WcMkJXd/tTT61rpUoBq8sxXUiprs+Yl4iF57ueQm5j4r1LF
ywVLamFxDpERwmf15NRarQ/X7m7lUd4Nmt04r7jI/SbTaGnUvWbf4/Vhh9eMpMdE
CiExp+yFao9Fu5i/VbGmTm8uaaXxc5dr3oCurp767FYhe+ZxzrcWJS4vFBH3lEwA
sIIuUSQ9T0/CMWf1lV7rhL1i3ny6ei+i2VPotL24DFxEy05uInPQrXqSVF4mWZhP
p1gzzcpHBEBdOF2K7c7eoRFsVoTkx8Si078HSU2HqTZ6x9H5jG5jzLs3KgKTlOqN
Vt+GHuPdhYaIpihl1346CrM1LzWKADt2fenViMRVRFsHl7C3NBQdva5FLbKhhUUM
3JXDybQIpBrc1unw/dPVRmHc4F2/5RWTRYT/PWTvxG7w53NRxw0ZSDun8VvhzHWb
UTyPLaD5qjszkYVFWhyHh8Sn+DvVURT7ilrb2fESVXHmqMx5zNXeGreR1yLhvGK+
OWLuj8+zwmetKZ143GlBNdfZIGhPQ4Iknw8LORg54A+3Z3yGIo8J+sq5W1t1pfG/
ZaLASLtT4OmKlo4bVD2E/L2s/4mhrPYW97X/Ciakx4H3HFSqHnA4f00NQSvEw1xL
XJxEF7tD+bZXAhrp/H6f3PraHSts+UOeSJatW0gfDYvzuB5qpgTOuhzFnHJQ/H0U
n524uZb1+ITMGMNgviJ0bKvjLyt+njzKQmF7ThNnf2tw0xlVrXIoQwFf0JtWELKe
z9ZMetbF0ndGfyZ46v2F+8uVZpQdXbYdMs+zLbGJc5gsIqhyCaSMsFwEq3sLDFgj
8qphGxiSCQtzO4ZzYrxj72+2m65p6xE83KKjtvbz8Kle39RVKl3z9FhLjgEOGGmd
9Ck7ijvTa/5wz9lJV0vgIV64zjhRZ+hpRyAXYQV3eQTjNHgstEsNB+gFnbIdP0Gc
BYjv8WgEx3qJH4MSOiACNsyeeat2Z8IvEFS29sXOdXFngEtdx8acPFzyu+J70BC4
TA/8rLnehiQOm1Ngzxl4dj3TrD4Rub8qprC/XNRXJyZt3E8J0U2f2fR6auhBkLuu
+kVqTYQensaGVKpeJ1fbgNh7UM3DMFYYirn8B6uJbud48UOqsJkxzDwFoOBG/ki4
LtPRe2kau/AlWr5KwjQSNn+L3fAqjVqlC1E37t4/8fGf828DkXHZSfzFDN8Yhkkr
bf1D336yRA5+KQb107LJWA+XtTuFuc5qjRx3opvK6TFOHe3DMjY7L5x32lbrwZV6
cJ1rBRXns/Htzm+OtE0KlsY8/8iAE5exWkPIYCldRVc3Do5HPm8Tv+RDC1I6GuQg
fho7s0BBu1UR1DIYtOIFHVHaL2awgXfN7NOORMIH/HdNE3Kx/1/wuOIHNgAz/iXR
8lgAhQ9ojrs2ahv6/7Q5BlxyU+EXhOqsaIzZoL6IbqeNNBnRRbN8u705rHZUFfjq
KAoR3lg8XU0Y4GiiBZ46ygXTg9qacMn/s5zNFNWs1xObVUlm6hUhT0/ETjlhE9JF
QtYuKnsjBWSSmQXznpwvPQfoM0aB5aF9DtZsFMKsolbzZyHDVSiyYkIM8KXG4soo
s01DUDdrCO0FVx7z2rUqKpzA3hQM1Z6ht8VnA3syeoHQ4jx6sAiwXrxNKCl6s9un
7tm1H2lsuwA9vtHsYDlDcuHX5C7iHlDmvbCcAK3VX+a9qOotahM8C7h9TaFySiQc
zjYQL8XWzSnrlK4ebyJPSDZVXOh8TSb0b+2AP0hftyosyoswqWtZc3Oy6FZIECt+
qzF3+dA84ByIxFZFb6JhU45g9WEcftH/+ePvvzpYA5zUeHBhHBXQZr3v/8lzbyiU
DT/6fno6UeyABqZm30rh+TdMpLlUZjKUF0P2jemGdC7gTub4wxwuohE95oy8aKzr
ptvWPa16EWtVKJBVeHjasDYaH896zV9vIINXzgyG6AAE7k8EnEEHFx7fJFXIhVZi
uyX5EtsCXqeTTc/mt6EeVeEBtk8dd9vzDTcRqFRk7wIK0SQFIqNziH3lvoXq/v7k
B+QcF8+sr4VGHZ62QY6RvvKUhe1yNSrgLVbHHglvRzPqzFvWGbW668j+HboAVyjM
K3rtE7HT0me0X3P1mnR6m1N1KGlPMP56lsMfb4/f+CFYjOIsw0I8oKDGJXgCs5ab
y7m4vwAJRaO319gmw54zrcUS9KPJt1FCyY7evruE74nO6f67JcTfRGEU5DtfgwmG
WVcvDu73qIlaxQtEStisYPy9g9adBHROI/+GgHPmF7o2UZ4ExVxmd3UQw1PGWxpE
i1DdsSSGGks5vWBDr2dWOvIXEIcdOO52A9pIX4Qd8IZ5rZHP6GvCw6yf/7Fgq4qT
P/MP3NinpF/neu2tu57U6l+sg/YpKYmaj7ZhbyLfipUvwM3OYwaQzbZsdOHWB3SD
1t3tx86m4puH/xcSIWvTzHMyXf/V4Q00OATiBSmK1wBQS6l/l4ri5bZOO3mjALzp
sdq2kMujHTRg7MIZWhOoqnFW0+2isLIn9pm9Q7SA42tON8whb5uIUsLJm6syHei7
pgoCoYF6o8VEKgVSBAKAmoJMz47SCXGrDivDcFlXUpzl0PHlSUD2CUBHcy/gaZmH
mqACBsafakuuwU5pVLBSSN1jKKpRLgEt/hZLB+05e7Kh24xyF5xJCIPCKB9oxR8L
An7nklU/b0vqx2EzQ+Y2xizJOO84pB9VOjZED9Tn63GsnhaVdPEyFEJJKUqwJuTJ
vxJFNN2DnmaakRFx29JpnDWtKdDtqc4L//UoggaVGyOmq4F64jtVwlHU4Md8G2Q5
cJxLBpx9+ph5CYO7GzUOMo4ZNi9Ao1j5nwF46dLjsmLxlpQfJkELSqtq2umvkD77
ymsgQLHNKvfE0BRXNeNH/Xd2d01ou51KnxBk693iVBdC5wH2KbrYr9p8dpIO6Fyg
qRDWaB1cNi9gJUpumDThEANFxl0EZjeGSVj6Vgj0BH/yj8DmKKsgOf9YbynT3Vci
KiRF0B0Sg0XUNodDViFoQ4ipSNvW2/lRFNpR86cGfxA3WEYeIlT7+PNHCszBx1nt
3QTHLa9S9rLX8jPvHqtgMzvT5HZPDFYGGGyKo+JSPFomIutIGYJXFFDGL1bqSoaD
xzk0/W3v2fJqnPV8w2FXOy2ZTAMD5b2iP5uN46OfZ2WsYmbBk+AIMFaNZCnPP5ww
Lumer8HhY0bz3y198RfPEEYUuoDlzzVB/vAUllcOaPR5rd0g6+PLOaJ9rgX66OYD
e3YwcvjK/voOf6Gs7+OmZRpS0y4Yt0tO0g85dmiC8NN63zBlWKsIDZYO+JcmO0AG
T1IRUWG60YZqjCFE4JcAvQ==
`protect END_PROTECTED
