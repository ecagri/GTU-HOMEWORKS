`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cJiCDUJcUOnPH7TZByvJSYcYhcdWhjyMOYF6Gr640JkhkoNunOmPSO50rf04eIop
h8Hd9zHjK8TBz24vjLVYnpz2W4o59X54uBocZ4vqpZnyyRk2cE02LkBfqdMJ2NEN
eo7atWYvEDlbTMAUn+L5iDjoa/QNjB2ET6i7N5ux6Av3BjacHYpgmAKMQ+FpZ08E
ImVftT6/IKTyILThgJQYXEmPmIyPkrzOJSCLkHYJ5oZQr0b/tzUWKMjmiXU7mqRK
2jFZDwI+UUmheXxjTrHizVuXQrSYpJWsJPZCey2hnxMnHKywuyikamlZgzJu1iXj
ena9D3IrQPBQ8OHsPv7aJBnvG2eFd6zpXYsnBG7M+AFdyAgIiJBXxJsM3AD6q5cu
rCgsfoQB65ZheEtZW7wKKPXXa8rqm9V9az/RQHwxaPj+VCRz7wFVCw2O9mXxA/m+
M9XirleB6QROoX49jKCjIjTk5V/7/cVQParAn079mdUvzUGBvknkZb47QnrJ2aPh
ADj1UHVEJkfSl/scT8ZKzO2ScjzLGrNujBW2vvcZE6Ma7DgdZiYjcRum/DVv/SW9
s2PZ9oGRJsttF/Xl7/1azFKcnygsymX8MXpFGrZgV2PvWu0RQ362Vg12YLBjqZ33
d4719oOlY5Z2XFuE7Yq5u8YJDnakFphAcgGe+bwCJ6cbjoAr+arJLLz/Q3ys6kML
cDV7Ev34F7h1pOPP9nm7oU25S0foc0bYPoQA8PRUmgE=
`protect END_PROTECTED
