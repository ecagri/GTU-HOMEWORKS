`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dQYWu5dmcHTWidZM6W07k9Mua91f7lmsFhurQJSLbRn+/CaMtMJaIszOWtUPyVMH
5lU/aMPWkOqxXuuZIzJ0MaO900mCYvMxmxP1it8hToukloOWc+n5ZOecRzPdixBP
HqRdTxT7zFClAvYz+3ivo069I0ZkQk/aEyh/fM56w1kwHUxxO1xYDZ9u5F/3b1sF
2sajAIN3bNc7rZBT95w/3l6GDSIvp0qag2m3rxvZi/zeHAMJW2zEJvmYzU0iwWJx
cDF2+mStkjj8Y5LiXnumyt+567/nohlDc2O+Uw2oeHbUH1EyiA1MOO7GpXPw2qSM
4yKP52pGicpKysZlt4fjrsfs5/bpsUHOOkcb33tTQwO57PMDlXxQQNgC3lzgRHlV
Afduyqe5i0O20/Xdons8qDNptLV8Xo56xg10TVijK+YQmN6R7YYybXxNGtzum1eT
yqfL7F5HdykHWZrHR1z2mcLyPH9GIka8OhMlITJOsm/vu18EIMWlNZ9oHCMBfwBP
zYJiYUJLqQRk9wKiqDCXUTNmGRZR5V63gU+ZkrE5U/9o2H+IQ7XOPkPUkeboS6M8
F/Hh+8lbQB6HDkKqLMepeLwr5jDfnwhft1iF9dYc+hAeuRVXGMiVv3KkKJkYWm4A
tXwOILEenMrTj0ThgA+PEr8eabP5ibpgnRfCVtqghhItaxRK/cdhUVYLjUncGH2U
BaGNfNkQgb4RwOWMcCJ3a6yQSh5UyFvhJtyHjaaNjXM/iMym+LgJn2oEOZPevXAS
sZhtgUHOOZGeC+J6ucS9Cm0lp9pNAaISLdPmdS7WXmQeBZM5wTFAqsndYrSJYCi/
Db1LhpypkLxYEl/Ia9FTfvTEEDqGxE0W7YBDYS03m5IN6/OJaASdUbs9tKS15gyo
FQZ3cwCbr+JH5YfYBGAvIPvfKiAFS2wQrXUkk0C1vfnuqQAA+jpXxUJiznC1yBgp
gteBAfGpJniEnUIF6e9yCwhFk2urkDrZqP4s69X30Shvec05qfKkhoBGdpGirOUd
8fQX3leKDxhuFOaxdyJ3V1YosUXauS6yz4z3KBFkwKKk7ZFmfgVG4WtT/TJxWXeb
tnSQmgNYOdGwEJC463q0Fdyyo3ZQig4iA1qbbXcz4bucvPCfoXBY/1P54I9IIeTG
imiLg1AhuwN1xPboiFUn91xHQTnSCl7+HW7MYzd0Qn8CZ+NOxiMV3nUjA4afESVy
YbMBY89TYGYkbpEi7zbP8dD2wA/i7mW45rHaVivuLte4q1S5Fs3ZAS1co30KQOs8
dHXAKq1bEncunbEZVbNR2GlX37J62w57Eh/vWvywohTSbRvR7KfB8WKjzPWU3ZQ7
jiJrZt1dIVvKKZ3XHv0cLxpwSH+tAwEBm9PKqyrJKZv9J61NEm+ov1M4pVug5JpK
SHdGvB6+mUmwPPPY7dPdCzv21vjFMpcTImqQns1MEpZX3655pn+YEnGjOOv6dQM3
4MZRYHEqTyi/9JhxpJqZveM9HfNIgbL2zhv4D42Teo1voIfBVotR6kyboThGakVt
7dfobNMhX12Bph2ThSS3EuJwo7Z3EbGZ5pMwv9lgtDP5/BmJgdhw4tC/FrB6RWs9
/IdyfNT2nD/31jjLAST5TB32wgIizPDnUj3LfRA2ko6mVQHaxAk7F7jc/KhIYbbr
HAMeNmUn4/U7oF/5jQ5H8tho23+Hw//4yg5A7rcDtL+zsY5EjZsHBp5Y/Fxed4Sk
6OXTVGWppZ4o7snUzyUw3lOAswCx+xuD2NJxQ0JdsGGfcBbBebxUZ4LN1MQpnnoQ
0fTEChDm05KZKutnGb0mtqSnjUHzfVz/W5YiYNc7dZGqDg/2P34QB9i0wpYvQAQ4
UA8vU8aIzt75GoOrIWQt4Qkme5Po5M9TpEFTZksKp7BlqWQKRt8VhWq1ocgJFE+N
QFPVukDWAfrCUZsdhdI8saY9V9BrM/VUBBbDGEQ1Ccikrbhv06lZKyXZZFJ/5qnl
tL4UUafoawcV2LSzwrMXJnTKswKJT0rLPxt0bU07TpWdPgbvGjKkRk2A5L7JX5oZ
UfoSuIDzJWRZtV7CaaCN9reAeEPyXiQZMaJvvP8d0L6K/M6qxZNq+tLMpGI7s1Nn
3Wel3VZksIxGPo7LpODubT/LhFica108wyD7Y+NsiA0N9N/DCjSX2H3EXLIcbVbK
m0xUAlKPBrnF289vfJzc/bMO0t54DMAmfUcwYpyoJ2g6jU2hi7Dg6QsI9YQMeYgq
C8XWiWxvRcWVQvG0BYP7AWWESxOOiF2puXlSq/LGSt0eDeq2+H8Q5NDW4eRqFv2g
6aD1lF/UcQKJep5HF7Xs6dWQh/2klov8xUoJEewoMS2bTVHdlXdYXn+6hOAmYSWK
YEjajzry0eS0M7fqLtXhdiuA1SkTj2y22R+ZLWlv+kWiOg/ee9A/597Fe9haHnf/
dXMyBw8BXqockKO6j37jUVzM4bCNux3tEoP6QbkECfX+yj7ZJvv8ftS4t/zWrTML
x1mMgG04EArlzKRtayE1whmTOjVAxFKjqFOBGow9rkQ/FMRI/vTXhm25ZYoRV4P+
HCvlM25dYQdJkoCrikmebSZRs6kDfYsqdaBMqfiPkgtftbvTqXJmw72RFa3g2Mlf
62Ko2NtPHa28sY5NuuO5Ri6ggOgLWoi22OesYCgxG4kqkROUloHgoGPwePQzsYWd
nnFakIBaO7bnUOInb5YuU3HCX6ZcYxsq1JFP4mkb6PzDgkvHGOEeyHCROUSYnPYk
gDepG0Ue0zz8MspEIQi8Ep53BGnfaG+FLYYMGk94N6KJAhsgH+n2zO3kNrunjGq2
sVn0goyCiXspTOrdSl9McYBSfqo4oeP/WqLsZ/k5wl6bwEWftEYp0/pDc9uQstQk
MJ7LV+C1EoFNGOU6+Jpi+Lq6mP/vuA8GkUMfFPQsxEStFYB1AkhFAHsB7GN3D0Wn
vOXkp8VQax3nNujKNsFjduYxQt8mvV7X+AZS2r5xcr+rRENEA+QUH9QndmuF4ChB
oP1Pgd+BT1OIspuU6Vww8WWCSlEClWGrF7fkSM5ct/koYF4UOYXvGS09jgJ3AMdi
R7lzODlua31ForTwGdqgKFc/QAp6edYbeJfZpTV2oXHR6TB7yjuF0LVxPpUSyb4h
raIniaWjYabZKuwtb0SmEpCIUPpqdW8tNfASBVByZaqws8L/U3bbsZUBMp6MQg1v
QUlRm6O09bFUgFxqJaBSfoA4O38B8SU6YEyadL3Py3txOUXOVNmKBL0qOY8LCaRW
OZx5CJ+mVUkB5mBo0wpxXXA/E1AUwtln1tG4N+jqEgg6o8Lbfq/w3RlVaF8Au5DM
MES+JyuEuoWJ4su2Uj6JuFvoIeQcPR7BxwNV9/mdvV4wI2TZVR2+Q2ZLhyhhS2TR
gFRoIWeNGjvldyVDAlKelII72tiHo6INWTnH1cKHH2H27OYtbTTPSm8MdXYLkQHc
KBiBdpU/Ylgy1ZQOSs09/0SAzC7rq9c+KLI6Iwp12r2mruHUDpqu4SyE12BPPqa7
mTIFBVsePhIypcgI6q/liud6ABgbmKEah8GcQAorXIHO9HmBbbnTVPmGzRp2CFpZ
w72gXaucEqoEJd01vVEYJlIDSd5w+jU5VikpZg9kK3EIa507w66sp9ubOtVc0WNu
HacpPHOpoj1iZONna2Rt5alo2WY/8UFIQ63CrA7RtOxccsYRn74nr36zE+i0izoX
BuqhGBU3K+O2KXU1oN5Yn6bJemo0C8F2IEmNoXQhI9agGU4FIQcEkUmA9qSndwAt
fxL+crjWu5FtUOHLqNaMiTfoGRsKadYFtCOGsJWk9tiTNvcWn0SZmc1wN8XTtOS0
OflEBlzu4P+ogx7BvQWgo9NilUZw5utnH7pQzmHa/hlbJUCJNkwrT8/7v9XWtRak
l/ObdDTotvsD4y8ZNfvipfqiONrsv3ESSEJ1Dt2PPcwANo69nefDGv+bMBh5NXi9
6svO777ATL61Pct0S2CXbt5Lmme/H9JC7trg9UuU5TONQXNeAgjTzMPkfVNXgq1p
Oi4KIt2NIiQtz473PF2U1XCJZbZNW/siws/5/ksLxDhoJL2KoRSg80yKgh4TBVzp
ZBrjmIXLG/JT9JzKwbK9aUom+AAfWQCyQOGIXPF3KrOIRj/syi8wsjsyx2LWUjh1
FionM4Cme0uG7qfD+M3xRDp+QnCDjycqFaAdygttxMGCB86+OJx5xW0+TfMN1El0
obniiAdSHq4Kmc8z4WeHwDPvXEQwvoycFN0z42temGHLtSqMHwRnzk+SSKKZ3jkH
6bHZZQ5ZE5aecws/SSi8ychj6+qIxD/8HqjiXB5uE0ftpUsZ9E+/5u35iKS9mpus
PsYD/QLvBdGX4Y8m8/dBYUgUhbi8gZSi0/7L9hlHxsZfIjWn/f1OX5z3RH+N4St9
8cG+MMmIViTZPueb+JfjLEWTkUQcdmTTNukmBdcwZv2+3UAHY9sH3o0liZNx64Tf
4gnn3AJDZfWwtwU3rpQ9Q/H03qC1u0J5ET1d//k3wjp8gD0+cH95oC9l72nSGUqz
JBb9K/dscJgyTOqF8VKTRzptR7xXPTFeT7oOND1qAt9H8M1J7D/vln75WhZNUTbN
o5MuxibgtLuRbHjif6qePl3oD2vAv8eJk1Z4J/ivM//oi1FGpgZDqIu+V2TjPjtD
nO9hRUwkqG0TgqScujqQWWAP62z/Hp6L5hM3uJbERnetqxYx9Z5qeyGfyssZCkIG
z+EjpdeE9yX+0jPZhh4CksDILX+wkoz78mLiBYSirZjnojB183U+7lt7eTZBGNz9
wg1SHZ3Vdk9GYAUM4iRCRp8Y/BQztUhM+VUCT0W0ztq9JaNejqpZQRBNlkHrgt+n
L6aJJuGgFVzU2eD9BeiPr+usxfA5jG7dlumh7eblsVLsFIB4jF/bxmvDJ6mzDIPR
l2brR1jE64XXNgw4qwLQtI9Qu/a0Oh2FtSV9K8H5wif/kCSditQNZzrUH+DEeFA1
igJVaYAOaV9TntbM9xrjUPuhdxsHR/5u7IJc8gALQlXEUEWyXIftrW0YwEMGhSws
1Mb8Nlbf3voDd0i/fmmnUyGegMzNPatKi1F3fMtsbkeSPj77f0TM10nBTgK9chZ6
pUnU9SUIbT5XYC7q/9O7F/2khQ5b0qJIeXpUo/VEIhZJ2XzAlrx8jQw/IwXKk2nr
qOqromAUFRcp3IxnRcluT4Ku0zMJ49tINKcKGKeAz4HXqyk1Q2f88IdVdTZXeEF9
dnSQQ2TIS9KGPykrSIXqdZZYMeAVt6acfmLpsg+xZYxfcx0mrvycc9Gi+HTVyNNm
xNml5jh6zZBL3gvX8FMUBtCpyISJv2wjSvyWk5XeUMbzRT3koHea3iiDgATuhFRr
yifbCkcUMk4sJuirk+xiC3dhw0kA4isfJ15ixVni1BIHd5irZXme3JOEdaz3ox56
PuHPFNUV2s2fVNeLgechjblwyAYYiuf4TnjXRz5JEVmrfFncdZbbSqEdPCabTXFi
sAerRf94pcD+hC8IAz8v11kAPRadu9iDop7sZ5bBqPHNvnd6VmN/gulmBxzIqh32
4kuXgKvYDYdW3kH+2nNKi3UNXGGsBO2WhdKxJtovzSgF8wD76FVtuuHkcEnRX0Ut
uW4UNVIku/0TfHyt+ruYfcRMIy3vVVHkLl2QdQ1en9WXdymCyU+Lb0n4QNhw1r9N
dgLy5ZvUVSZNYwAGs561EcQf25GIXfCg/4NXnSkjzdnCcmJ2Z5uIK0hTwya1nUcj
p4LVPWPemYdrMlFr9bm9EDRbqc5kt7YtA4Sz4mvRIg1zh8WCtqBd/pxP35qtvRpO
ZFHBCy4XNk4zCmInGML/KU/b5H2qn2o/AihKvNdvjbfgKhKYGPBZ8sGpJL+zN2Hc
IEtLcyUh4iA3G6+GgBu7ks8D0VqJuJXTVtXUiDB4B2f+YSkbpEhXCxJh74SGCY0q
Jw04gKjcU3xlRjEZ9vhfQRfVKfley9YOogwD/uG6XqY0Gaw/xcvDRlRPb3YyCdll
CCSAkc1U90+hBXAFvvEezRHy8YfVtupAq3BTAW4//qmOyDHH6jaLQjjfyOwKZyw9
QnAz0HbDKiedfUsYMq58Ig+Cq6CbJIFYpdfjKwH5TXASbKO4Jz+/ZXWzPpWr7rTu
LL5WDzcs0TnVUTrR9PZhHQ3dfBcTtVOc5PLCuUic1E9HocfAEDEBOX8Pnu5hPy7J
zvHrhkTQMbwIrCa+tNTA3PCbWY3d9Fnwuoll89wokYLxucWY/tJl9o8KFdBBbmGG
IXZEaFRzuk0WP4bmflQJaCFebaxSdgL2Xpm0kfTNu3JjD7ok/RdOrXv7QVtY5PGX
Op2lVtxV7E9Hnu91qdt0ftULgDlLBedcoXdpf3Oi2J8=
`protect END_PROTECTED
