`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t3AZ0f4Y+mD4iGefEOt0IGyRnb1k04vB2xcAP3KFSRcHrAizh7I7bEwljdtG/3R6
pMhQl8qTjlAa2StMk2GPNyeG+UeG0d0UEDYGAvC2h5W0lAjTAjstZ2O2BSkDTfVs
8MsA8YsKaU6/9zgXAxughySts2h/1AOhTty9uNWMQljstDxOU/CTvBBMIBxEQ6iw
bHn1GJAetNaLqtYi7ZmxeVfQ76duU9NbyV2pv22jVzEpB0pylb43fcQOr1+1jQsU
Hoy3UvXbdRNTJYf0bIZymhGksVKHzFGqs85Zd17RYCq0o0BrnBaZCzsBwG1DRfNO
aQojag2HepEkiEgGWpnCQ3iUn7rMS3xb7/FgmfH1sb0698jB0pmFBR0eRYrUMG+A
rnt7Lr8qO00c6deXoPXkUsOJEPOrgBz1nOsIRzbx0fjq5ribjCWDC80KT9QHkVo7
LkTdYSwrOqXsKEEvNSPitk4H73WEmkj9m0fbVa8C2AqBy9koz6UQ0DM3k0ly3OV4
gj5/ZzNhoE7iVD6IOodKoXbbWWN3SWcy0nAvoDe2Pd94OUcMMDoOafIuzT5Yk5qs
xGfVOh1r9L8RqbhIZnyDct3vhpc4WzlV3YqkZ3CH6kO8IXpTBYVRG0+TQ/+q8maH
Y1sR3OmV2823YdRY84Mu/Uj41GP/01ACMm1g6OGWk3Hhi+5zRUUjEL8Km5K+UuIS
jy1OC4ZI0hORbp0Bb5ASV4YmXF1o4tbmBDiQlSrS/PpoYsZ83Xv7bx2bK7C9AWQc
EEa5A6/ODjgsa7eonjJwkXC08koosHvY856A8A6+WXWUQYpEo9Ep78NWilWewSit
FQ35M8VaP6aTLHitfWKJsDqEJJUPBdciWx4Twf5XOAOsRaApJokXuHYOPhpKKpk2
EKdplymZiunc7obSzJfAK88QpkOIBHBWQ8sjV7T7S9le5CMpZnXFgMG/ZBS0//p6
cS1EDyM7WnPrfdIryoIXwYQBQMZWQmcqrOIR0bEE10Yaw1DLn/5t+XhbCnkEeBGf
PjTkj7qcnTeR4ONBo8BFzksI1F5JjGX0fPlZAsPJP79tTSKboeJ/gdSmYN5sRDhk
UE5Xxw0MRJJlNYaJNBDYpqAPJrNRQe2q3tVqJGZinFe0l3cOcgkZEIx7ob92NlCA
tSqgrSQqzw/pRWMqUvFhQ0xNtzWjmU2NV8P/81uhrpwvBLJPfbk5Gvgcnj1z4qkw
QPlzFJPgE2zy+e+7R+mL8vTcJZXRwjJJ+bV8axz9Mpdftrn0ag1OUFcdRFFhr+PJ
9Mw1R1p2izsx5q3cCWS7kbUMQu8uziYDGmK3dnFiTq5FXaZCiYVIkHFbxOPjofOH
7eR2d7EAl0RVg38fS7kYoHSF9vkg5rU3Xrx7dDGRA1wziPWGEkZmtM26u1/dbMK/
vCnCOQhFZGxevNN3E0RHGoAcu0YMllulESp3ftBVjTX/cN9NvpfvPEoGCw71EPML
kF8jBBrmDkyD4aseumA30E7RsTjSwHTYLXxQQyRPADA7Ntfvkc+CDtboEcBtpiaB
7HYS8U/l3sQ32sVYAAAftkdnAR+2B56r8QpokOx9TFwmIyebSEQ+DiZdlCbQ9cfv
DaOSXYt/+nod2cMaWwZYhJSO1GdNFVIxuCdu7PXnjtfJon7bfB38CJMMrOBj6AxQ
7mpg5qsbDtagv5chLjmdexiac35kW3XdQXZHoCT3UWyN3UCha6KkUsAPBH+CwOg5
KnQAcFMLj7lI+3q6jfnKSNztEIIZ5KymdlYob+9B5/5E0QtwaGpp65H1FhS5cBnE
sN6idA98dDYR+FMy9VDC2EV18wmx8YBhJSlVoVipypGGV807TGWVr2MFWRFKZXoz
LPuTSFtZrAVcq5oB48qr5gMqbQlxgrbWe8KF6skHVqaJm6UNfEQ8hMa5z5KlSJSC
1oNLKOdmRCyOoOyZIgdx7fHYYl8KcJGCpnVXsAwjBl1nntxuVuEqjo76LEKbDAss
9GMQBsXTeEE8AR5iP7o9Ohwi/vK03ESD5xOdoEc9Cp8gVLqWK0DUxBXrmMJLZO11
z1D/okFm82PPSJGkSFHU0TG8PuXZv0xYli4nge6gae2tdQ8LgGcKJZ2hhCi++DZz
27YH3Yl94lUWRDVoxTGjhl2B4oNguJaq88ejlFSKCweVGWuMfZEVBGzszq7sNJt4
ygiTaWOo9g9JmadaKxXDNMbK7Q/+x0Y8FSpAKImoKjLbZfOcKXq5Q7XRg+BUuQnf
eD/iDNQw1TwyoqgCiKtFSw7fRaVvbo8xlUEfkFAtK9m+tRAGmKNoT8XscPJ2f+SE
akSdNG/FY31jmDF+37qKO5pFTXSAb/a24pus9XVpYRljeA5pEHmc/y8ooyoRwnC1
er88L0wbuNgeJA2jZQG/dPqjXAOXlfKxTxX7Dpe8A7gX4gPc1Etf48q0TM102QZj
Do6dlS/faMWkbv8/T9t02FKjoDDnL6Er0mN5EllA63LNr60DlZBN6AIdeQ3UtD1t
k/0fWEaJPqLvJwKBDGrpxuvSki8VKVyXg/rz1su9FNClS8UvZWaYHI/bM5mnBn9B
O9E039TI/kusHYkRlB7vHq+RBPf3JapAD9VMbJNGoww8Krm2nj+RhXftmkvuuQqX
h1NFASjYVJ0MQl44kO1OFefaeJ1gIRMN5tTb5Cv7MBVdfUvWkS54kLi7LSxoDGyK
ilQxC1ZLbQ5RbHb7I1CYGDPKutp+wGVApTZRLMDCp+QUzxcKDExjd1CjIgpEAtTU
pSkvi54y5/PHpB3fxbnaQX7C2cwSGYfUROoEzY4ngKp62T4gpaR2ldILGyEVitxo
lDmMxuDNkWMmt8lw7M//Axr6lHNyfjGYIZMlcnByWxXcNXSLeaJaOXZHHFI7fGjr
nmcGuOFjznbdbCY6TY6mPLx66De1Y8rQgNQsrROsAFpKM+C3lgH8s+iy6NYfNdfl
rZAATl4M7uMaFZrA5NES1OAbJWGIWto2nqrHcUNxXv56r3rL4Hkncbd+BdCopfAW
pH+JKa0f2OnlSnTlyxQka0Js2f1YgdQfMrec/z1nrkdr+9k6iZ6a2MFOq0KkOTAp
gGsqpLPfe1a/Is6kuOYn/tIyZxtbEPz1SeAmk7pIvvaYbVrjXCQ9JbI2rzj7Wqcx
52qv65Yg8RtTc9CYE7rV+WQcRkw9sx69D5l7SWRdq6HCA+yhlXIP0OgcNcJGDyiB
saoz6xqqNLMi/B7knJ94H0sRU9nfDpePoSRpedUVQxWrqtotKZnanGoe8+SJPszi
tDPO1ba8jUB02fpZldCG9V5s0AdIVWdfbxwfeEGojiMzBjyXcIUDKwYgAUkrYF88
8YnN2FHYrjC8HYWosOelMsmN7ciDa6RXLEa9+B4jliiRQZxyPizPmcNyrB5tfURG
gfwbld3v4z9ArVaIz9/oio/Asgi2pbvZE/h5WP+Psw9H7DZXI2mg48U/2tQbdvpm
BDsKgNUyMm70S4Mj2a7Ungu9s/aeYEmGnbJg5MeZ0iTMfu7nc6m4nIMZDiUeQjH3
LH1nvzsLF8rsW+Qj0H4/Vfgdpx0XW7cdpAe6gGYsZiNWr24bIr9/QL6kr6EleslS
Y8mY1kNv5azzpWTPW4UovOnZ7hyB6ahTNnutG5A579YHxd19PGAn2KXqLuCbHtDS
YfgdHPWL7my7tz97+N7efW747XH3aH+2Bcco6KTlBjeI0vJShWin0fsH3uAqjT1C
cOOGP4xet7A4/i87o3SaAFs6urH4yZPuAxQjjW+/lhl19n8tZTr6rRgUBh+pP98Q
uwRD7JCUtu8k7ATE3tUM1I9d2N9INvnvlZYAeeXKmUJpS78J2E1nkWxOxDPy34HA
J37lVvu8IL7+vXzXaEc21i09UByBlalmqdPUOvARVzAtk+rmzwsjZlmJ5pFjwu6+
6P+IZW0uB/UWHSScLNfXvEXnO1bC8kcHgF4nFU4mR/p9lswaQMMC4aueLFrq+L3a
5eOFzyK9bcdM6YWSr9y3S1dMXRuEBWlHxJvJMoa3lBcj3U30KUlSlQQoFdK+F4ro
mSPYewYpoWwWelc3AyOqDZ1yjTcy1y0+sA4IGFBQ0Pw89ykQc307DF3A3XW9GgdD
P1ZMpRE4xSjcw3mLzziUK5Wfy5NPuzf2dWGcDEResHOjiAiPxY4zrHIGLid+LI8n
tnHx2AbfqT5jbFuSl44kXBoD2PokV4H+4bgB382WkkEdxUHRMnxI1Fu5onF2PTwe
RjF6hvNazAuwZH4amn7FyfAybSyFDNybU2vvRtoQmNu1oedJHI/kK1oXHNGmECBp
`protect END_PROTECTED
