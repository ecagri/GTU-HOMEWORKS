`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RbWvqy29KaXl/3UGEhcZj9QHCpL/uxvEJtqZCeVrKgfb536q98ZiTFJPAaFUay1b
eOqmd/8VwfPhH75TpdCl1VZzH9DCLm4GKEB4HAP/rabkxGmsppzXhK7zQs9iGSko
dAQ8otNAoXymnobUbw3zT+Usq5PAvnKbtdjETx2kmCE6hhY04nbS1Im9tr2f4/zA
d9vyBoQey9PiqMJAL7QcwQq9V+s5RvR+pY743Q/kC2dX1pnDypaLIorGZQ1HqDBQ
H25NbjZ9V+y2+JKk4Y1B1UgVNsU8ym0zYFQ0pgBz2mkhyz/mwqs/24ZVkr1mqQ3q
A+5uqzXGBMgK7E+n2OoMFMRegdMj+CfEnmM6wLnclffg3qygW4KbQXjcORRTnNS7
LhxRUW33SkLMeHFHbnP2h8R4rGNBPPJ/zCKmYmxZVsTwlfb36yBg1qZm/+STBJEq
KtqOEOV5ah6Eaj7F6GXJmu7gQDimrQKabwXrS7OCNyaGm9JjOlIWjEWiA40lkWLs
3XhhQkPRtEsbRGyOBWpEXs40kf/3MrLjaBnfsuoq2iffFV/tYNBtXEhXJ8gze3x+
A4bWXbkk5rLzKrgdTaUmu1bk33kDyhfT55GjxEmCM9vRqVQ0v0QxbVINtJvjdg3O
Uk6HDxdGE0bblSo0COLeTpT9HfF8xaVBAOnobuGJzzZ+YyELygjCScz5hZqU5J0D
jcIn1CD6hebw7AHBZm2JKKi/CcVSS1nUsSQptGOdZQehcmm2iJwGSceqoNsiX60C
kzd4NjJ9AiXTEb/rNRLqHlAelGg2uR4sRdRwf/oeDIiN/nJnT+pXxVZ0mvLLayMd
ANpF7aryFDX7/pYDsr6iCFtO5v9Z5ZXXdOIIFWB6uj9x5bEMXlt2j/TI7dkKwr9T
TexO8ikGJK0GlCJRTZ1Rd3sdUI9os4IRo12YuXTDYuUccFAeel+WewMUH+csGHva
gTeaDhJHzT8LjyundnAX0JE5bRWyfOTtitB76iAqDtHWpjk5CW2EuA5sHvEaP+8t
GcX48uIa/QH/X61AoP50WzPb/c47/jTA39MnCB0lNbIAWI0/kequOFKCrjptuGKW
aoGDkOz6rFp+rftRhkTvg36Oo3flte8oIBxeJmCKGrqAkBWpy8kY2VT8Rn7x8yKZ
PNUR0u84Pu3uDs6M+o6xk2Skf5zrlzHaTn8afck+U/AnUi/ZMURn9bqI/o0fgdRy
YtQ+7Mh97D9DVySJsUwf+dhJL+XHtFsrgykIUpwM/ABIaNIOrBixGU2Ok0iGeq6f
WFEoNtO45Pv0m+ogLVNdROuzkNY19TzKEaUHsb4Al9evFYPm8FhpEBmskcXCA6q6
JqBrkbPM/+w7tAnoIonxT/qN+49XEJgEGDJiQELonfrItp5jWzEpD4IEkPxMi36J
1noHtQkSPvAyiwhxKoXLlm/AMVTWjLVIYXsPObM7BwIhOaDqayZBMH8+eI/ug+Rh
0GL5IrovIKvykK0J2+PdRndCXlf1W/8jqn9cF42Nnt5MxOvbyWcHa+4rUYk6gjHz
Mpq9mosRJ/IpqDuNHiV0VnkA+9sVyPewlsyPanYlOixqrIDZqi5+Ko+Fih2izepD
bBCHciHiq5upfkT0pAhmZkv1hZaYZ/6XIJm/tCG9A+apkBQ3OJ/xd2E7bDhDHuXB
Fb+L2HoUSiTTUsJlSArJDgDjFNVRwBz98ShLynvsfOkgPSGF4Ks6z1WfO8HV6OjU
gTOyBDy4+zLGzirU1t88xyxuNY2yXaBaDkOI5Wu/YBfmmZYj1BpyxAX4jFqFiL6T
uZe1qpUKlTyyWwQ82yDA323EeDlrgbyFkolsAdgTV5wpnbUJnljtpbaw6z8yXPas
yfZbb2IR5O0ZxbvZ9nJSr2b1/vUhsnOWo8oYOkYKVMpFjmQo+P7crXJb+NF5k/zs
Ip0+tL/ouKZEBQOm3FnUDn+P3YwFLmOT3WZvHeahJoObZUW/67iihufR6ftPJt+t
yyX3uYys8PGchsbWmQB6UQPb/HdH+onRU3aaHdZEixnRslab9OFd2R2hKzr9IZ1M
3qY6XeD2GTfL2x4anqKQEuZ5YGF54Eu2fma/bXDXJZISwHI/3HR4y/gl1b9sv4LX
rW9W9TTOmOvF4bh3BlPCtilgo6xMCeTJ8eJl69cdemUngNM/PnKp8GAHFYbpcH6s
JzgVw0HcJIbZ9j+/AmEne7WRavECUWdcEzSZ/dhSAAk43i8klJlztQ/F9rz16SGm
0PqHp9lr0STpQUH6NJn6EKy4Aws+fJNtzU1AfhovXeQXBZE5MQdGGbH6nIXDOOpW
vw7BTQ1d+gwUE2EX1ywZPCCOTdpP0KV1y/36ByRtO3FzSo/jccLQWi1QyAATE50J
gCfYiN0HcAHLRcZbk9JPBNMudsxDQUFO7Vqi0zcsdH31HkHhBA4kNvUKmf64Uk3g
kCF13FYMcVhPwcMGw3IWXR1tiWayrYgXDIkG7yuZZ6TxonEmPq0g2QA+gZo37Zei
KpEBGup7ApC1XGeItHLA5cLVosicZemQ3mAiUhylLlDjXO5j8AoPWpS+S7qMMDUr
6jvaMAzgZBt+peJddfD/mKFzmD7wHQhdT4aFU/UPAKvtvGkGXibO4vVYAnJfHY5i
uWQ/zSFYnZTzCVyQCxoj5W57+DO3pDFWcGg7ERhr/7hgn01Es963ohHDrMeueWyY
Fy7D7dzwZLIs5Ju9bayozVRZLEjIUTmuMdCTgxnYhwfLIv8Q3slh90PSc1ohh62c
Iq5ODfKswsMfmC9nc94jg8dSLZwcmvGG3UuXNIuSwCoOZNo7fpDCrmLAm3q0DQms
dfHm0CInL1R85Y4gx2/eMQbhaAeZ9Z8dEUZueMdU3QeMdN+wowC80EG+VUsAd+zt
pGY9z+sV7TIHAJA3f0VRfjBpAPtvjyu2lsMyFSdfJTg9oV6o5kphf1PjFufZk763
M7P2YoXAUD0TG3NT6ox8IU5qk4XSOkkdJ8rR3sdDgzDiDi9JxoazCP3M6BcCCoRE
IP8Q4seo+3y87PkL1lJJXZ0Wx2q+9Mj3jfSZ176brdbdagj+91hvWf/RUSDYJVwF
lCMG2gLW0E45uDfqP98zrFq0hc6DNvziZvwaT5/fGlPk3J+WWaGzzXEfQzpfIrse
kIueBrty/mtHnhdacGB9sgsvXKOqtFBS6GTEgwHXT2Zk4ykW4eG0BPb8GKj42aF0
h1fD8FM71o9UZW61FMsAjbG9/hl/WV+rBE3LXQXUWdBDHvHAMnu9UgjBUsypJxHy
ZPsseti0SsXqVjgJe80SdmkYmesTagpwSDuBcLt3Q6z1eaBtDGT/07jXrk7sDxiA
CCCDQcYDwjYAr9I7jFOKPWihEvP0tUvo+57kdzUBVcfj4QmHb7fkW59cr9J5FaFW
CzJoL9VuyoK6bJtXQNlbHUdLbbK/Mn6dYtEVukyYtu0dpNOc/ccdNJX1QxLWbvsk
NoDre8o5PlWc04KTg/hnxlK2SC38NPfBrQLbtyyEb5U0sbg3q3X4BNeCp50UQhDC
zdB+yao1S2mWFAWaRz2LqvEYj1bMdIzA8iA2dvSfHQg1/s8EHG9G0+FJwFkWfAy6
/W+al/ZiNuhgtKz0P3hqHpCXw/hpAXIWYpxRPhDgx0nt8BkpiiZIbmjBlJouuDxa
piA5mox9861a+NIRO69K0WQYFRtDt5CNkiCVGaf3URO3qAgt3oMqfDfBuOeCrUsC
J5Bh/XfEzC+NCul67gvQYHctVf8AEo1kp6E2NqFGuPUxawv2ei7H2uh2Imq4KYoG
nwizI4SRsBHQD/W0Fus4CvqL3bMSpvPxi7dwCc+yz84q1WMs7v5y6QqYiSd4sZjT
cwOJ73j1xrN1sJwLgBT+HUEunHAAbEHqVm9kh3UkeZNb7xAHUKQbRcwCOY6NjYc8
cWpuArwIbGSJpURcZG401vXAAG3ffLQumyEyfawtjbUdGmGhWnz0pnfJZkoaMN8V
XiPAukCu3aND8yYXmrUebZObsQzioGMl++qmXO788WZ5vzJ5zEAjPikNCytBjMnu
kfQuQ858/odXVmJmuJDd7U61Xnh0hEEnfC+wk53XUEAKnzkOQWrC2om4ywjgj3Fm
eWyzyPe45pqf1tjMi4umS0+ovyavaRVwUZJm5BYi2gzQV8meizYd/grzr0luoPid
QcqdZF9Gm3nXb6dmWViKjd/ooYRRHbg2NayEvvFbkKjs6VvE6T8HbSZSdrQ4l57e
vvJ1Qas3mDzEsp2MidnA33tNTZ9z9Mw09IbxN7c1qALbBrsIjojk0ftxCBCsolbu
mlcs/5xAZoL7voFPzWQQMddtAjbO2UqSOTS4u53w4TTZeAVovk9XwIb1pk4Jl4Qz
KqIjQJ+CRuia9GC0QO9Org09klj3QIu3rvrZFoqrfptKiB6H5OWdksMIC6Aj0MQt
HBISEbMhv3H7irBMCjELk1gSnziwvZ9FriHD9kh7a9Z0NYqHzExtcFZ6o/jH63+M
jMDuapIvR7DYfLTOsvJUOsMBaadCX9B+h7F/dqRsnMluMjM47ghMoWRu6vIJnEBU
35FYwtpRux3WiQONtLtURgo3A0cJpl/OPdzUjZFRp1i1UfP9SGwRRYKYgPqkoPD+
vKp0CCVAfTdoh/lIU0YY6eGbcGJ9CBDJHg7bJF3G8hDw5ZbvFnVEsdYydZs7Jr72
D0wxIpM0L00WG9e7UTa03fNpL1lu42mHNQ2helM0eVKIyjZ8s/spDcyZTjrpSH8m
bEU4Od5wmr/mtlFnl4DqbceQKybaUCg1KGCFJZo7RRaJf6GpYp3w/AlyGJ+IIyxg
WsR5jOc4pMvW2nI/f7ne8bqZ6mHm6cpdE75ODoe7oj31ogsulRyX6UILogthsLQR
ckkBwhzy9h08dd9Z2W/95VtVv8tTbXmnqgY6pp4uyKDso/3u2tY1aYqQ+LX0CkWG
xPg3X/WZZRjaqkyOeYNvf6ZP5m1iYdLjk+nSyNJVrWWcBwzNJHgnF11mDIYFGJ5r
bK3kMiGzoAn+MuCEG3YITQ6fta9ZCjpgtvexc3cqD+Eq3k4pL8zdu3NYQOIWnAmz
9nrF5wvigHvaqxAhLitEWUm9FXpcxaZo8ekEgqyv+f3AGdsuFLxIox/K90v62oI4
n3K2SFo5PFQ1ZiFCxOKjhkj7tgE94Scu6SL6u9mfkpjOpMFQMAV/bmC7NjQli5al
FlhidqTvHkB1+0QmVctmj3H/xEA5KdehJsOeIwAQZiioDo+/Dp4w/omBtK8uQy1R
dexd2sUi9aZ8E1WdJJJ2TwTeAHdMGgecbnpIcxVf1PE/bC49MoYzrFLd8zHZ2NoR
3r7YRC0R+dDU2Gjp/pteMVXtgy1ZvDkTNnhOGGQgyZCIWguVw3qGRjGCDHnZEnwX
E6GlgDk2yBg2ae5oj/sfqwMRTcwjlBTe+1oD3wrub0e1TZLB3SDQiWeV30va+UCh
Uax6zmqaV/6paexagwLtfNqNQZExikNbZ4OC+NYfcvgKRa/QNPw5lKqgAje4w6ZZ
se+h/BQyzP1WjxwisfsAvLLkPpwb9sQUmyYVbroKbW3aOFHubvVPqnDzWfWaAvCj
VLiM7xCzNvw7r1MGU/DuSBzH8CsBB6oczVA3sAoL7tiSh3ei11bprNZToMf41JzC
+bT+BX7QhoXoO224CowQmg==
`protect END_PROTECTED
