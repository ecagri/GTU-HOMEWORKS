`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MPqQGM1Nmu4qj7NwFzAHJBThLlicyhLTNAd2lU6w05HXoxpfTFsurNJelnnRe24O
uc11fSbPWWd2bqQmCevnu/yRopUhzwo4bjKsKve53tFGxPnAimnStUC0Ks9UHGVg
BM/ChrTQquvY0pSXnyyH6e0ENpjdNMPlZlnP4tlQ+VtnRzD5Lrc7LImXexto55QM
MxuqJ0b4iAfjNiLz0fWnxJ/oyqOc4mo1Ksji7cucHImGqIvqz9dV1p1a89Ex5XHq
1IwN2obvqOV0lmEsGF4CE3bqtQTEt0vEqwZ6bKaLBlk4MD5IxhT0F00Q/mi49FF5
Ak+PrJyiRP1GfPvZuzZE0ZiSz1m4a9Dd2ILxvAOLZ6vvAoaCo366rEs0J+lD8DFo
RhcUNvebdTHmhwD3fNXloXdsnv8XKECV1jxk3ixqe1ifKCLVTxctQGecqzoicJhw
wpNShBKPpSxmIuNLX31YprIywMbyvhivNGwocRobpufA4pXus3dhU3M98Mv6Dgpb
rh5fl1WfRpF/L85r43aPE0SfeHnPE/CCthqYkJxzY+yzxE2LqHwB06Px14i/vacM
c0U9MHBvXtKoeyMHjAPMWUkQkKenbra+7fDxQsvVAJQ2wlK48ibTuI+uEwUSDP2p
xt8PmUCJOf/Kajk1TrRCRnyABtnsn8azlkvCd1MM7714gA2bgeh9/4y2pfl+v9Eo
1kymNAoprpTZOLS4nOeqqbGdJQewtYF2l8qCMGgUoANnVQ4VtkXLJZRL02fSUFZs
5dZ8bCNWJo7Ssk+fg5Onex2hcalwIOO5Png+yp1poa0=
`protect END_PROTECTED
