`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5mj9w1sns2OWqZvqDryPImyWI9ACXYWm3pg2E4scFTNsTExbvyzmRQaxQ/dcanJu
YViMeVvYQX+OR5f4iZyLK7xs5a9bBNPBVALU33Ro6rf38Pz8hqv8ISmBGGqiCFRg
tPXtIBMjh8paGAV7xMb4ySYG4TODPPhiF/QBtxPWyHoZuORnWUuzXklKZBJGUd4b
N/ORYnpC3uuz45crByX8b/bVS/+Col1+nOADZVcrY1Qj/o/5Pq/G2xktItAvZXqA
dBtH4y586zNWI/H+y/pkfA7DMKnGP7gs19IHR/yZOM3AOqBJfITAC8Nabq9A80AT
FroE8YLpDTNXOtw+dz2w9PXAcxkLr5xfABCFKgZ4ODjZTkNCDdzVMGrEtwJP8E2T
3rB+9zPdjcMnaCx+CF0CHD8zn/Tiakq0KPVAcgceKK3v/6QNjyIuwbF91XV5ddgz
awFLKGAzpGOZbDacnDytP7phAbpgliG2m8HbV7aboSsGnnCu83CgQ3Ybwyh8t2xM
J17MJC1OM6WJ3odVkzifn917sEyBjf+Hr7V//eXP1LSaFnI5K/AZ/GdQZ66OJTyb
aWgO0g5xZPxC0nIVAhEOzOcuyMHRIBxOzV9WDuqrd/PIYnurND+RZUpmBbmF4XMC
w2w+Sq/BRm5SpGs3ARx+klWApAYQu2vFZtCOE7+bp9KNTX2JHa+gHXbB+/v1POPl
qJNenC+ChcB2KV86GAC7r+AcTcrJi5+KZeHBqDOex8DZu5j7larJ3o3FGWrB7K8s
gMEz8WUZTKbRgW6zfA4SJ/UssHeuxOcE8Gq2V+gHFVb0NAGIWC3Eccu4wKz9w2m6
GtPKck12FH2fmlz5pMS/UDiO2YvgdPEgsrCEdTYDskvxWvPqOxphmDI/fbCPsK0C
B/dciSv/R/ejdmXmkcAbmEtLNfg62XsZsT07oD8zyTTzLkXTi2ux12Hjl2gEUm5y
TEwShgCSn3UJQ9J0NZWI2Y3li1hcOw82t0v+fC+kxwG0mU7g9rRMXNMQpC5flu37
mW+qWADLp4tAf/XCx+VhGVc5alF/B0IsxiVmcxUlz7DGwTXDlRSXz6S/PSWPK8FB
DRN3CbgGRVCuNGrrirW1BQZ6TyuEWxqkYs67fOXhnJRSKtrT5b7TFmQzq3Bu3tb4
Ph9jXUfMDBW1lshHu+sVJnbpEV+/oKjR7dcl2oBzkA832BS5WveHrdTWEb3wlMsg
kgwZDwX1bMjNt1EsdJ7UclC2tH/YU60VZjqOD31m8g+mH710Ldw3pfZJqjHF7gty
2J59viqDlx3cGeHjgSjUw1JkJgPYfhs51sw/+zCHUzDXooj2aX3/p6Yij/qH3/AR
sx6pIBciHjVYk8YkdAYCjIJN0dqZXBNCeNCEIqHe/iD2rPDqoUUXa5TsL/CObb3q
g2wGTidcIc+U40MVTM68+uZWk2+wmsLM5yFZvi1AMfASKunWsP+IcmXzkW51Jqhu
OJUOG/J3IrqZVXO9KTFfxcUyZIjBxrrovctky3ygbsJXZQ/82zPkc5k8B8Z/Dnp5
1YC87FMr83Le8vPzcvyp5T+De2D87gVDEYtwiTYbjb13PsdrpMomkFCZ18G50gIU
/HnhepxYp3vfhFF64Mrt0oAsCvVmrwU2WeuSVGDbvb00rv5fi9RGs9dlwucT10ej
mb2d58yZJfVRvxkO3dxMAS+Pfx0L7x2VtAzKyqmT5FWrNuyVIVnRb1Ki7zYaUGB7
yd8lic0MLu1gDWpIQhKok1zDqF0gUnYyIMcb0tca9frz6Kl3JWQHqe9dpj2zm/rL
xTswrUMUXWT/wtlYki4JjOL0rsoWglA61jap7PVvQhNhUtY03j7Kglov1Y2ZuaYE
twsPVOozBTxsxiGwpsScSmEUd7XdfZFDPHsjN0aiHxGH5HwNWTQX//EYgSN4ueuH
3rdxFgXudXpaaTHDwlgT3uWH70SF3E9Je36Dg62JvJ8zL8H+yRhNk4VwjXCsMTfj
n/bnK34PobMr4cUOxPIsttus1kEvxrfIqk55KOll3jkca6T1dtGnwwxKiID5fH8M
2YRsujK21/n1g88Z23wKj5oHCljSSpMWRH7BTQpvpEfGa0HOwHmQ9nBfbqEydomS
5TS0QWB9IbRMqaKXBBg0Aw6y+QE0FrOXhO8enwR+rmAFp9PZFr+WlJRz/k0nt9H+
zWV2T1J/35eyPcOvFo9LnTy1GGFBYyQ7yz9PWpGMEvbF9yHf8DnJX9yjU3Lkf8PB
hCL2uI5qq0gScitxqVxpWeEZNSseXyQ8CGTt3yQNf+236cPrhRuU0p9H71NFSL0o
XiJ1EmHmkx/B+tTIP+65oFWkUCgtzko3i0sVLcdiOJ+HP/+J1ZOltTirGIeh8Ug8
Btz2F0c6oFh+AIpOvgUrXH1Ijg6s20RNSP0AKKRpfWZWRnkNXmccXpfz/rHy8Zcl
lJO2L9qPj6ztxW9KZLMUfcl3lc8QhZrV1RgA5e8tbu7vZca5LJmAKp08OqwuhG4v
Hl9FiT23vgA3Hb3taurn86zkaZIYbf4MivhPXh5DdYgAwyRlPW5hjoZr/AlRnbl2
C6Uq9e5UgvSYgyVVAABhYFITpNxAphI7usQuoX5hcwJgbXiX/qtpYACcPhcCCwry
mc//9qb86tMd0SlmwU3wrPlnxlqF+M3v40+8M1TisrJLpRc8VIwNhu1zyMsvdkhJ
8xv5AVItg7QmpWImFMCUwzn6E1SauXS14k4bH4OR0eLGy7bvxWhz2kcWC8DPQEEy
x10HK+y5n3ccoEw5OJTE7BbnevwFP0Ut75nNiL3gAlOgQfTZpXyRpFuCPtyEtr0J
G1HbcdPVGSFK2k5G0VkR8FQaARH5nr0EBc46iFnXG2Ct5Y4i4HIURyToS3/04hHp
OIw2OflxkPSylzLLz3vUmoFUr0NIOrVrHDMuzV7oV6e/nrZSTdTXI/tcbDeaZkOf
gVuLDO2Zqt4E5VQysIAQ+XKglJLWOG1JqjXsaBbufdw4KfMYRprldZXaWTcfvxrH
dZ4X/jmqev9azp6CLh66RdtJY79Qs7WVYON1+FZ0wQsSEYdHaLM8XCnNmsyN6bq/
ohWsF+zJ3eXZqqaWHyZojCCTx1PZ6hvXdq22QOtps1ky8H/LXE2sR1SsBz/rbX8o
3WjxkDzeNU9qwbgb74dNQM65+0Pb2P10TxM2jN8axMbCvCWDjWh3xqJ2p8QdPiXI
c16Q8cWsBx2QugojpmZhS2Xpk4gpANGvA73O6LXN3DZQSM+752peDq7sFFxDYeJt
xMRvuEWsfRd9hn+ZQGKi60g71a7QS9siXYx7r8N5RNzCM1kRp+g9mJw9efn2jz+A
Xxq64JQn9XOEhK9DKO+/4xNgSrzJDafcJgmaBhX2AjyqIp9nxGLe07DuZQ/sRRlx
IztXBfupysRMozt3kyIBuY+kwaOd0rCjGUR/8UiSZmdem4RY3W09YW9TvTn/BIE2
iTE81GAXo7RG9IuN0sRH4ehLK7D912GMf3ANZt3ifsmQzeQystvGjSUON+qYc+yG
BfnPly5V2bUcIlRTHmduhJXlIaKAZFPOPjQgZ2d6EkIFA8hoD/KPkBFIf4B1b8KT
uckRBxscSiXrG76pYnfg/FHxr/AlsoMnztYvIdAGT5Enr6rQOMNjmuZ9ISs75eqA
zsgBeyKLzcPbTCjzpxICkL1pCJM8gnxV7XbE01KcNJnNrmTWkTDidgcAjH24DdRF
cWVjxnrMjTbnuQcElSXYTe0i5f5X3vJQDv1ouTWHhqyRk+qB+JSToijzB8QWrgYO
vh0eIyDwf0XQRNZkzIACZn+oCqEpweGKwV501QjTCK+PCjRHCQQqpxoQ6mr0Y6O8
s3iLQhalZP7r19Enpm3lc624PjWizH+h6lWUy/PSxwJSE1IWAwOkH/ibOiqcFBlw
AVtXSoM+d/zXz+8FxHrOyEOyauyMTZJKDN3UhRyoijSNw4pbP26B+EXueDn+qu7d
nd43fCvpxT+zwD1yMfRf0pNmcmuAqqY9x/qguaNrG+602ZFN9yOkFgdjo02uhNrn
GK/ljMnSwUGPZB+8uYY8sHkGu8h2uSjsQqYMC7e0tlSD/28MDPkVci9SP3zzaIT9
UVdFLxA1gsG8m+t+OLJ3K4cAaZQOZ3VJjQtw+uKkXpwmJq4prfdYlpqRSBCeTCG3
46KrFZAJWPx1MvrpuOO4DyT1dRyDtp2qPIvuc0c5WUpzOVWNZPki+TaxPk266pbI
6k9AhiGTeD1Tul84N9hpBSAf2aCYQeKUdEWVfXJ4bVMWjK5Xmag4WFRUNJhsL0n9
14jei9zAu7UjVlo2PMZHVjtftnzLt20t6p6xYPuSFSTdAwIvTG3VOsMHRusdjQ9f
vgFi0xocH8ySKBdLUAX30l2ZbVfkN0jV4Y/PespJnaQkCjS9QpgX2p5K4M62fSV1
hx3hzsfmEf2ivd/TL9NqYDkP3Cb/UprfNxm6rN03idol2xJAPfyWYxRh8Tdn8v9i
BOVDq7GkfXSGq8Lalc/b+FAzVkKJ7SPKxGDY5idUM09I0sa0f0mPUG4STbwbkw36
pZfUYMDhNiWz/jYc3oyIrRj3EGbfBmPJHHfiqLr797EuY3nw2UFaJiz7ZWDMxOX0
XgemjCRcx2CxwvjlJC5pfeFXJxNKmsJEhHxC6DfsTzqoCk9vexIuH9JfMqZhvrKA
7hDKNX1s/K8LwQKlN8DUWfNOUtjUaBsoQ4Bx1gXZOwTW+tYEznXCF8tIb8Z9374S
Y037WEmuzvHH0Sf9gJuFW0lHJbSFiM7fyiI9BN7oBq27gR7RS0oCBAP/6L7tmsZw
pPhFlLskAsJ8azTzpAGbVgtqtIktGrz4wKD/VdMu2d9qeJWPiIWpONzY7NKagnld
E2YD0J/AyOWhBCBfoC9cYcpEqyndzKNSDPAMQVwZvr/ysl/KIEQu61QhYEVbemzm
+M9A2wKQd48A+fTxl60BEdug/x2VP11rSdZFU5AJRrU=
`protect END_PROTECTED
