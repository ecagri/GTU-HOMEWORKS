`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3mo9TEj7lL5pE8jES+sxPKAJ2pDQpzkbBT+d+iPFcD4EBYzF6Elg/eP5QcLJ2Vi7
tl6NXNCDwYbnr0UQrCSWreBZDxZF7w/2QCxJZkG63jFg6HjeXJASkiuG607SNX+Q
XfMJyzGEFCEAPXK9SdSK1k+KsmObZZT4UxpV5xbhzEX3iGZEYAA5RELAd6MeYM7e
G8IRtHrR3YNcSXLJR0twn2xDXoz+BrdKx/MzLpe6OiJ1PyOza08WpKvtOBGvKefW
TOBuULPpr1V8XwvbveCbj5kXCL2TgO4SHATUfJO0z7y97wrQ8NhWmg6eom2qTdPT
h/5hRRCBS82M+U9rv8lJ1YtObjMS4WB8lLlzu9AeIz5+fvu7KEcWaXS7hvkf55Xs
w8PSPlicwGklfILYeWG+/b4W4iIqwxS+/qYudgnvJ/0xNi5b1q9cUbojSkfV6ISV
BLyEwxDivC11TqnKmA+EnSRIaQyz0IeIt6JcEiNSQbAoh/nUFyUM6YrgQlfpp5ip
4bGTl68r0ozAOsJ7GCbfOu4jAEG0HsPq2eDKCbFGB0LEEwdQK5aRpfIKz4T91iqI
ZaIUJkN5kJ5xOyy4Hfsf+xikQrVwCrwGPgKDQJhem+i4VTEnIbag9dy35NKJ/HO4
00tLLm+j0poMBYiJ3eJ5R8eg6uTGS5znrF/MhnzQvoxpcfp9Uaeb9hThHXjQCNLs
nVlbkKUa4HzwkSasYM3lTnvc6t01quQ2bPry7w/jA5/4c/JQ+inBt1IHBUQbfRrd
nT+VGlPt+g4EXKbJLV0hpGbjeq3mTZ0sHKt3qzxVU+Fa00T/tDM6SCEy9XoSlDnN
Jjd6uWjK9XkTGwF5YGN2KXwwgXHmsJdAalOoviOvJebn9R3+KMIDLyz+JL3Ntk1y
sGHE8/cfNzeRXbFZHe5guegTnELzyc3r5KcHVRuPvCNku+8jZSpwQhvAzdmtpwgl
MaNeVEyMwEOhTcnF3Noyw3kCNqrB49KrnU2Mao/bvQZ56fOVFgqQdERFIG8+EJiD
l7bz8Uo+3Agi7NvhM40B4ddtV4tcj7ayvZRycE7nOGV1BHYYx6zViqhlQWaGiPR0
6cg2Z4lj2iorYX+632b0oRAhr82bHtvWfIYSi38N1zPFPQE6/HJGv0dVXKTpKtJI
Zia0SQcfAj9ZlMGXyQMj4lHbk4VJGpxVyz3nCT1GdT1YXUj3ZN9WiDmqJJrSYHi+
rEUNC1bN4crVXtyDkWGQNbuPb5vYmnUH/0bdDxGiZYKEmRvqmeUfOOxR3UmrpeRl
E3QG3NM3V6T3cdrDOjbTUFsNuHbWw944luSM/IE+AifnVktMw14plNyEhA5PqllR
LRJbu1d2eLUBA6+wxywsm7nIKsQYGyhmLKNs0m+w2o8yTk1Q0/cFM4Ih/EnFxByJ
yJOMeueSLUNKmRme+jfk6tVNla31T0974uzsOyhw8xDgMJfLP97CWRwGzYdUx0t+
1aZNngeptaFzUqArJIrA9f34FlBI36VNKr/IEXZ2IMHVRtR6UzD5C6Zy/Qhrk6/e
`protect END_PROTECTED
