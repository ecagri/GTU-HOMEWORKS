`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IHkFPg1H1lGEeh90UuonuwOCf7QqV42l9kz2lm4KjVHUZ20P6okQeYVsHAER3eCa
6+cgYPs4P3UaPdAzZFSrgeXCu8hImLdxC12uNc9Z5VzfQlkIZyNGccMnhTh21Eor
6drkf0mZqnYiR6fk5JX152nOx42RVk39WgNleqe5NS6j4lQA7Y9WDLownULOjKRk
lyP1H2zTgb78sttHEYO3SIDS7SHijm1DF+dOD8jooKdsON99znwD74IwptatoTHw
9+jcbAvWLUUTk6CFKr23/mwIEreTouc7p0awGZknsi/i9giBvtEvg6F/cz1hf4Bv
Swzhv+XId/Um0razsXTGavX7qz6UAk9R75RUIUrmpL/VchGwM7OopbgCNkJpxAlp
Cc9r/flAqnuxaeOLlErOtoRUKE2j7pH5Ap9RUTjNva+2o6USngB4/bGbPD+MobRT
3zwQDqxo2tvRI7H+sSrUnGLBr2BilvXyq3MQNCwyiFecuIqKdKU7tTVrNLu8TncV
Z2SGRTt/6siFIPAE/XyoE6OfJ/Dw5jYuKIFhaB4PySBwYA3cZTLPLBsbJP4R/dvV
TOh5Qvf185Cz+Ci3/wh+HHV5rcNVEWQBRUuKNIs12Lc8LpSHZSkkoHAUJE3GLCt8
yGmUgdVwp1pRfLvUHnCBMu60Gm+qnx3T0pLe78IsLETPmod0seP+COlPGjbLlgE/
SqQqDI7dtcws/xQrqjbUCJjjBVzMur3VLe2juE5yMiA=
`protect END_PROTECTED
