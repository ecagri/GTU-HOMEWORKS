`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IxMDB+IeDGHaiyW3VdX0TDFuw7dE/j0XJLhQJ9dWb1Po4PFSmr+hrX26Sm7YjEVX
NzTiJGpGqC+jRCsYv668gj+VTA4HBFCEmqgsXStGybJlhCvj0EK6rtlbwjcjFWcP
j7s52LEX0iXFAaSR6j28+IJc40RYjhplzNnf59I127KwcVD7Rt7DHlAnYLhDY15G
T52xu0cyMuzOI/i+2Iul9KiXMUBzosJlQ71LYAulvdQKyGnPJr04FJZ71HqCwcBW
0sKNes24ei6CcGTx81Zd3nBIWRU8pKTmdrJKjvMJYUZJzZACo8EdanX4OEwEeKrg
S2/Lw9HCBd+oL5nKubvcCqIXEco80y8HICwySfSMlRqNP9jjlLWJ6ul000JRspqC
Dw41t/BQw3rQ9naQN9ZTnw2DGLc+J3ojuvddK1pSrc3qf/AkStvv8vEEBjzz32CV
xDxcjYJDJSyUaBIj5fRxYxfGFf8Hgx1/VL1D3TbKVq995hqjeFllpoxcaMYd04rA
HCAVHVlHGpxJ7VMfy/BOipQvP9VPR8yBSiZbUuDAbynk4zMh55Ig8WLAtM5bUVk3
qs0XVX4rWUHyzvwRnwcXuuiQmzqd7kyBOpslvIcawZv3vCgA3DhaPue/XpwyvxJF
I37YSHtbvCWzAxVDZkCCxn8/b+2CnArq4mfM0/lcm1B7bYTVhAJdec6fy1lQ5uzJ
NNzOo7M1C8mLFd0fQGknGy/i/S+Z/OsJOE54awrsWk+4J1546q5qYZCBGvpeLhgW
dFJFqDhf1VV062d55o5UdWNbkRoA+EUQDvyFQx6xfJPbBbGljrAbCoVU7hzlljJV
N+ws9DC3nALfegWhP5oAnlhunf8Tfbsp47ADQby6WXKWt9+4CqxVHNcG/gEIycPu
+/E//rNschUIBVQNP9kq1ZqfGKPQeg+0d4ddY9742ARWRiGJ8pWDcisOQqz2bhNK
gamV7k5C7OBsU3ERhchVfYJvAVsDOnV9HP8xQVyM4NiNiGBsSCuilsqgwAnNilTl
W79xeMY8Nu9+DEVEZRdfdYI/JqbTkbVJjo4aGceIIJ7vv5BXksBW6AbRgpR0dE3o
eeq4NC1PqCZZSPpgu8opTCJWaGoTj79bSfj9Qd3004s=
`protect END_PROTECTED
