`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T9ZiiM7wOg1ZOmcqHGOxbkRUsU4yx3JlGG0XMtEXrR0aKXzi0wqmJFaaNiNWTsMf
AU/Cl4spA9DLuC3oMxJpWMY1VXZULjolF+11r205SoISLaMN5bVy3BEfDgy2d8bn
peM60r/FkYiuT8gvyDysRDD+Eeu4lVGWLDghaJxqvw6NOQLiuXnqZEsWppKHytMC
FRSH3HlINgO/fzdfMm6nB/Yx22edby2aqbIF1PhGbm6xnow2dUT8IR8bzXxGDtcI
S1meOroz+KZ6gP0jXKRXal6uEkU6WemA6wqyXpZ7S01KTG3DZcrPHZAVNorYXLw2
pP96e3Skw/ES00oxP7bNB3mcFSDGZD1ZFLD990UnwTWmTR9KiFU0EUcNqPYNW1qT
Wx1onXSwV5dPyU1zH4UCwzQa1zNgUH1rqyndHY0Wx0uvg6bvUIp9wgqeKM9aZSQj
xm1+2yzee/2ZRc+lsx2gMLa1sWxeXmAT/LuALMfzStnnaIr79t1OpIlSJ43ZDzj2
jJOyg4A1XSdjBVATNjIqIJtLbkFJTx2zqeepaZddloawmmCLVvN2CFUk9jUJmDCN
ks2feQz9+2FjDxr9VqoN2IYFkHzm8uZt9MiTaK+fCWTeUwU2icXkD4vaEUlOJe7Z
FvYMhGgjERyUguf6qiRMaqoB8qWrxqbumb+80sQvwmMDa9UN5TDXh2Nfyn9DQARO
dHJ4Pmu8VAiDDwsdC98zEyLkii6XW0orO84dYRcziMv33SP+BqbsZYauyX290OOz
GorvaLADyHwGtj3Q1CEHE7NpFk+HUHUyaSEGG156Ub+FFnF9Vr1iPkvRAN/bZtGy
JMtYKUS+epnHtdC9Vj7M3NHr3c62w1d7qFyCnGAxiXetPq0Yxl8VxwiCm3r6J6jw
yc6JyhVyxFdO1RSr9o38BaFqJguymZhB6HZupw4/SchwOx+R+5gCWVlJHkos5vZY
6mrk98UdhW5VxHdCwwPuNQXYKoQQyiB22OJZcQ+i41/ASBEyKjiNC18tEJb+deZ2
s0wjDF2oyHJYgdjrydPJfhqaxvogzheEnXsm+MDZNzxOErhmXhtzg6BNO0gSmQ0w
5PKagp73avFyYMMNwyOGrH2DU7DhFpsN/CtithBFjkno7Zqh0kPvD048NLe33pL0
AOu/1f2JgBwe2faw9lv8dOjrvBNkuU5PImBLQ70BXPmxpBBfONPjTe3yBkyq/BsY
g0egPOwveXHUSlnCGBkHK6PwuwMtFgnt5G5AoC114E/ZGmAa78dQVDFafXmsyMWw
VQdUc6+M+8gz1HrFF68TGWyr2i/gDMNa6FJtg0cTVRJ/ALNJXv/qy0wGyjiZlFJq
abwTq4B3+fopPPBX57vaLHFRG4Eg3X5nXwaGPOfapDVhBvqWDvtO4lVGfgE9sFy8
P3UPyQtN4S87tC0n+s06m45KVISEsdnG51XfkxzdPfU0x1yy7iRMG4s++HVBjuJd
hhqZNjJdZ94U6m9v5B+I1y6BSMoLnBvP3j5rgyxIPR6+LnJw05sUn5eOa8gvlUHa
5gZ6HvrTTsc503P7c4ZcaYjqLVGK6v1Ak2+73dikZ9fKvl/YWfDsdZ6nLbGQymWZ
jeztbYaV+9Djd1oRXSDhbRO42FwyLqFccanM35q50IfJiuia4AHXOhN51lRqeSXQ
qySGKSg3mp+HeB9F+VAXghAY4+yfyEcMEnAaTSOSuU/U9OcLmCQepsY2ut0sWdXv
LkBm/Sv9ZiNzNlT7GPhDX06XbL46WXps7wDdrCqOo0DcmzMjglmPv2zEBu3Qa4rY
4afIFOBssgL4K/NtYe1T7j1VU/Tj9LTuxswBowrBUxPZpAY3a2gGfu0TzsfHdEIT
zMOegaXXLexXJVQGGmwcvrG2JnW2hqP+ooNJIa3wexnYF2RycrMqBrEqQNIrZzrI
z5CSijkSkIcKgqXexqZJteePMGIttAKyTvfyj+B7v6pL2TrHHyY3tAJWyjtDEaAU
FVl+I5eJt+KPpXsKpsZj/audjCUiY3t/Mizko4GyO5RZOQxjbjlZbAW8qOwbb69s
fyOkBb8od/csVUUV3fBmio3V/T7Fd6aHVS5pIBn25CWd8rv88jlzR+xizkz7kpng
5pi8r0EZqWSnCOaa9H/TrQmm+xShQj+0aVi6/PaCu1iZPI7U+Ls4KbdLeGeC8CBF
/kufejIlWn9g66SzfXU+FVNy31O+TuBU7CQVxiz1X7Q9wndgwxiKkl2ciiie3sAS
2ltTOymCAhUi9BJS4nYvZMYRfckiIOAaYCpigq4EoiHhns2FljvIO9O80MstOHjd
rKmuwSesl2A8zYG9Jq9W/kvQXqGDBPzFgzzobGR12IKy+w2xB4iM6QkGgWMUkIJn
dH/ZSqt3Skhd3FwurXhLdtXx3mHY/nBNFnqxB1XnhvMeW+/ArVLfSUwO92r1Dcq8
ssxLjDH3QikUPHZN5Bew7zJ0aviAkHFCAQL6jg1mESB+vlkjNoxUBkV6mpqqR3qr
X/ML1L2us/ziOeR1vArfqRlbL/tfitCJ7qZu9T+XQGO9dQMrPevwuxc/r3I4V1Pa
jagXoKSTBfwJwBJ2ybtJZOmif60IRZwoWqu5X8/uoPmWeoqu9H1E8vah1IQz9leK
db4UY9v5Ks7Q71Rx0nbYhhu6tguLG5AUxS0AGeOdspHM1ovsXrz/lrwuTBq3oqps
IDOZ96AJ8AJEyxzZk/lWW3LWxNbeLroheoEHq8DN4hnkH6LCkPq6rZneRxF+GZmd
OFVp5N2MsccuWYa3OYsnYlnYikbmE+F+kCeNtX94LaG4Ta1Zsa2pHd7srOUGT0fC
wDA678ILTxGcpUU5iXXDZZodstA+EIqIO1gEu91rqhGgjnC2t/qNzITShbfG1tzO
VASzpinazVCvEOEyZS7lJq1VuAH8p6r8+t+8r5qeEhrZ7gCw28x8e7sY4U59KfsO
lNBGGiFUSFtbQ/U3UrDCUAYJZqbQ+zlXiazVagHBOPDV2sxQiqyz/X+5QH+hKd3y
KrQp2Za1V/zJexDI3E/r+3cFiDTIwKlRiUaiEu/MOUx/GMMBeKqKASv3PRoOz1Kz
hOhkxDiHMqOTDU3V/6fAOYBhYk5tZakSg1lw+j6N2CaQ3IoMcWIF7q4eJ/S5madR
6yX1oWtBewb+aXQAa7iekPzpdosx4b1wdpiaRvkbT0yoERf9yQmL0sZclI5NzHtG
dIpjmHUTQVSxXcs3JfOqi4pcY8qPM/BL45P9DGbx+6xeo9kyVLYLy2J4ZPm1bbDa
3vWdSRvN+ExZnBbRJyY+alTDaL/MX097ilLzqLUkyAhX9J/BK9pvi9EOwuwNz9GP
rtjxs+Y1MzfBor8juweVd4oqHa1cnBlAfoWGhiNmYMDlcRFRiSthAhgCqsb0YbCY
NMK1fCla2S8fs6wgEeU89wDYLBx4XAcQ9hguDk0+AwlRN0khpgr1WgWdM1IzogT3
la7+lOORUwjmeUGl/KJcL3qy9W1LoPBxEOPEJA3RtjASHyVeiCV21p/uQlb7Usys
XkU7+BqNs/63TqSAIY8jr9S/XWsmmTnIhzBO315Arx1zCNOu3DuQEQGtsXUs3KT1
zhtK4pUiRE0jp+qQBPe42Ekn1GqIaLs6nEEp2nrJPb/RPgH7wYayiW2M3xm9Iagt
nshaLEwaorHqJ0VU7o0upnEyv/ybyaU4yJqpl5RvmPxzuIMvWL7m1XfEvzpNu4+d
IYwkAsgPbuq37WrjFU6KW/8ai+MJX1AydcJbv0pc0abT6SxYbYoN2jXa6WgVbxU5
gqp2KHk+UmnyOyXONtplj3/tKdo3WtgHHR9gziQQ3QQ4E1kblRq8y23th6L2/J9s
4MQeRwu+c6hkF/mDd3uCAjjOJW0sC3IqL2jK50MbMPiA4Ogtx1P4qbpqqmUXWJ/g
tZ2u1nMiFWBh/ISKSv7piMNSCgrAskdflfAgLB3nZEi2qx0MiDJHkn35E0/Of4qh
7E+JtcNQ8VlXrE0GaPaY0V4gP251cDY9UkhAIm0wl2bQ10snjyvkbaKQMnDhtED0
8+LPkyJGQsVAUtXUbkQ86DoIelmGuylVpt9GqdQJc0Wp69qzLQJAdmCwOcbTVWIu
qRxbniqxJieBLTj3qpgOuozWelFe1IaaQbM3+/RVqkWKF/gySvaiLNHjM9tGB4/E
IfaJ51XOF1BpxyUTmFsk2Xx3YyTNjFqBRXFT0BYThntqSkZBA7TlhWoDsJv036N+
BL+b8fmwU63gyZA1+hScBK31uqLLVwCwPe3viB1NDGVp3b656dAB1zrF3eb8ZSCk
52VxpcXRzlmo2vwAczCtVHgbaT1ubgQEQpvwFHD/WjP2s+5HHPQ0FEH2MM1HXMlE
UITaPMBj9bcWl7UKFXk+3Lj7NcPpsugLtPKkiosYGvypRsZWsuj2tv7T8vwaVrNc
fQEH1AyLRUiUhKEZZiQRz4vXACpM4wWq9Ol7cvGitWmjukbyStFmSqZmn/DbWulA
kuSpI1HOzP4RQ9quVDHP0qpsXHECxxhpy5ChWZjxfGJE3H51drItE4Q8baxXfZRv
DKbyqSHtA+7ektJZeUsII2dikL6beoz+0rHIS3Y8i30zwjF2KAbSKO+BlVAcOBsZ
F8OHctIWE6abXp+ZqUSM7leeX6NH4iTCBWnQ1gyNa/So9CSO+05Ric7NNPK1/LWl
eV4G6jNExT5kkpvPDgzTAb7wh7+c74wQv7cu04KeKqFP2ElMRuH3LbD6np8pYt7A
Mqn3YYHBDNlwf2Tz4r2m1XV8DCGU9LhAdeo6ERy1QxDZP8ToWcP09KNUeIe3FNzl
gPW2WwRVQyFxBdrUIXkLLCdJp5xG3Nho4bo8R8rCTj7e1q+TCrW4c64BY5DW8lP2
RVOzK8La3CpszwX6o8UCLMU9vKCChB+CGOKzMUBZmvO4JRabkc49mXq8E2gbftd/
P2h+i/Oi0xTyhq7uuqkwvLoRDPcIeB/Luw6F3MIYv82IKZWHveem8JgZU+mACTsH
22wB0ICNp4t74MQExl9/h+W+EoCjaGpiuGyzv2E8jWgvNKbjQw1G4t3lZX+RMFpx
A8lWDWJPewnW4qDEdazFro0h0BXW8RAT7NGFxmQF0H0lxRT4De5R+gab+FLGKF8G
llFJZCCVxspnOLgPyVaU8bGXZB0NM6b2S1kbLYAzSWeopWbjwRsm3YKtUI7bPRnE
UJrMXB05yafr2dMEH+gtEe3b3tLz/ehDsU3YYKFuQNsKS00q3j/b6urAgtiUAAYF
Nz7Vu1R4nFzDBlvFmticK1ty+MW7heTkx1zHkerJdjdZ+7Q/yTqlrbGxkYnOP58z
wfwX1kkUPN70Jjx7QQOeoBfPRnLwtpWalu/58ZIQryxEEnSIlqKcBx7pxHkIi9vo
khiy+nlHyIii7XYjiTIMipE+57BMykuzYl9ediZlRtj3VD74/zkbAAI8SVETLYpF
Q9ApLBaBGsuy53XB032T9DCPcO9hbGrO/EkdmzWAtRzkMlXvqyYzR5T4YFtaKNqs
kXekfOz4dSShs+lPJods8ya12llYNiCP93pCYYxf1RHfkrFP1SQAb//ZVtN0YD1f
RPWn4ff9pELyIZJvt0Anp/+LvapkD61Sm4oLLx/pZ/0LhEDaJN8ZGKj0R94+3j5t
yYKspJJ7GgH2lvdmOH7d6gvg9G7KBzm9xfY45B2JJhHUNAHnKTvmSrCdk3oHNGFi
19p+a8fnGvweJ4ztW93/zi5/i0gkMkXgPvRJXfaFAhC1Pr92Ge4hfzP2Us4sj+1h
V7rOhv//6ATBwBlr4ZaGH68y5QCV4UQ2O1lcWAgfJeBh9kurWPWakVXcO3T4CItE
cUTXaHtDiLO9wwrfT4T7dLRAsWPAfI++oUtQba/kxeKzlr8BF/4X01nT5WcCHnvX
3SSMNmrLvt4OzlKRvhhDA0nVms/9ysxAO3oX55JbKRm10J6tcZxtBzq8W04uPyNn
OsbYQ9hTzLv0eI4mjnh0oUqbWoEkd0BhjKivCD7G2hggdJWUBPMuygFjPt+C7hma
ojWb+zNwQ1R3YClqc9c9PICWSCdeYGyi+WlYYFh7V0Q=
`protect END_PROTECTED
