`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z2q5Ez8wu8MpwXosjtrQSazbqQWKskBuZMCAm4FsnPiK+0m0jCeK0jj+aaLS0tV4
iH5LEBet6txeZQ6Hc65a2+dQ/UlRRgeHV1mXXS1v8O1La4b7QgTyKVteZG3jK6n5
5fP4wEMDzPnXoaiWuMwIXjp/aPEG3e58CRMM4ej4iyOLiRxJu+8iNTuoWvwXkpD+
35RkiYwNMsRlbrNpomPvjU0gqXAkMf+JnrxYFJnAu8RrKZr8kNrawXaAHnSTaDOi
AvK5sbtKdcJOZ6VdK92T0HfJhKrouJWTCOOBVguD4T4guHFa0KTQI5Do4TFQ8G7o
3UjeZ2nM1mCm/wmGPkXVRmzkSaQ+Ytv3sWPcCQemVEP+h5tVKDoa03+h4N+m7vP7
ZxzkHVIriFnaCyHNs4SJPE9u/BaHUAPa2ysK8MQC1EdgytAZ3MOI0vSZqvy5oaud
6F+6+bd8gyXD+8IeHnRracdu6THPoHmnCJg6P/eO4tTPyGFTxRAeqSrw+hR0EJ7J
oLTemG92TwrNs/P/KLtL1VIzujzEPzorSIb5c4Chuys2zotGCur3R7wkoyCXYlOZ
X350Fnfm8S+jS0sh3TUffLRsENS7v3vZpAOumJftTVxID2YihYIloBWobyIqORgZ
3f4+V4EA6Ze4GuCM3kLXp8kxkztXbvIDbuFOohK/nhDR6VgAn4XK/Hi89DCwn6Cv
uea1qe5emf7Ys3kos5gqFquRDCRwwpUbDi/hUQO4eJtK4Bw2qHMbJ+EUn+BVPXBg
SdHjaWKbzZ0FBIYeR0N+xNhNuw9F6bS94nlEOKz7sbKNwpegm+8bQApFdAXFb/Lz
Kqgv8WStki6Hcv7/6cB+ZB4ThSi0OecfNrp/UX4EITV0XlawgSH+9o1CoFC0r+Sn
UwjXBixCz5+IdoEnjKaEEImE3UF8DhvW5uhEup5odJ8xHG6TT3e51rjhhkNml9+Z
lN4adu7ar1izFkTY5zvQm1VBeEQ3exjHcXDmtH35fmLytbrcAzK95t64oRHTrQTS
HLpVh0qsNliSk/SW0sR+GyobHWKQqiVdYywmPhbTOxOOet5c7mFpNfZEnrRlNUyo
KTKaCFvcWuYRKSSz4BBUDQ4Kip7ltT9t5W9iMUoIt296gees5HogyXmWlML1up6u
R7kBaPlJOSwKU2qNOC5B7rSLYpf9lMjRHHFJVwXFUgoxultGqyLtg4W1intI6yqP
uHGuZdiiCKbhsemOQdPqLXPGvsRJVvgh9uYAMzT9dv0VZph8mWEgYwDxThPtjJ86
qltT0jtOUuBBLSlZhEBwRggDwmgNzopbwInlXKaKY9QPf0d5RqWixuzmlKR+Ja8V
2bCqremN/A7W8CZn6OTgU5+0+QoiuQvmwdrX/1BEv5RrPeUqDcSRFkbqPo+wokgA
T9U06fYRDD89htbPKl5mYVXtiJREGhvR0xu3HLEucPFCQNKcos9H6cQpodA1iO//
ZLk4tlwQJ0R0mLYBjyY8NZ62u7i4EtpNendrXRtXSOMbqqA8f57q7c4pUyhUzLJI
RBBt7U2gVztnD+pBWfAbffnFhPkduNYv3SYrLHHix0VDyVc25p29g7ZNSZwbEPe+
/wtZ7WT9VidemtWZZdShvP5PKnSxB5bTgu9tzsJTOxXLOjpWH2mT4DfELNLnnbQI
WT6Zo+jBlogb2vOyxh2vvYPN0/TSu9To0FIn3ms+Dw8xei7hp2KKSfKkZgvL9lUM
Vj1Ht4VqEZycFt2MpBNzEhlBUT7LZTV60tHthT4IIKBMrycgeqny/DflgGGxsPyo
dD9GVoDO5ZW1Di0v7Kt4cyeEE17MU0wo6ixXmNQv7qPq0wd6Jd4ttBXr+bcT6hhI
MTAu+K6zBg/aeEymw+5hOMZh28oIeL0T0yQqcch7sL786xJA2VPTzYWORyNPoP0c
PmrTeyDhRGg67Sj+LzpNVA==
`protect END_PROTECTED
