`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NJIAPbXV36l2oApLjigcuNvtPE5YWVzJi/isuKMfIynFS8h1M1811oovX5SH9TAK
lmJnYUBq4fqeRxmvPzXsvUDX7EBDV9FO71AEbLO2DjM7iurxcO6C7U3mPobiDVyF
NN0BWb0NPpiPfkLQ7uPXK3nZTdRMw7Mzv4/1FvnmiAWobyMiGCJvOsRPB7x4mO1/
jfk7dHI/LWBXBDTeP95hiR/Mh+z6koQXVaaC/HOyQiBuuEu9lM6UmSLcym5ZRGHC
0U97+gZot7X/04lm4oXd9XdJdMdNmkkhqDlmLPCna54nDGBczIaXMa8NLqqRaVPX
P8NGOcgv0Ag6ZMQWw8k6e4tGV2WB9K9klr++iX3niCL0g28Q7TOH6ePzDqjaLaTT
1HlYiYfuXcvF4EZJXYfZ6yY6JM9SKbvh1bfwCOxpp0xlJ0AoAULX6vMYRfXYNTUR
JdH75X9lkFgkBEdAhDOXRjV6RKfZVpn+FAO36uEuE55rupaJYAm15Ih43TQtnBmH
/450PROfZTGxdGSWN+3a74fIQ5qpSQJq9RMj7C615StMrlRN/h16ne1Gc2D/d1iC
dsf5+sqjLJqVcsDAWg6U8et2uX5/fXK/YKzhi8EeTxysDE9jBp/2Yx8wwWrcIg5W
IoCH8QDpaPxd1E84OidQ34Kp7TkHInJCxUImeEnEhPq5vSXKn0Q+UypyBGkJZ5Y5
DF2jF/wJY6IL83T77mPhMJq0qd0ATeW0lgEoBrMg/Ba/NM6BAHzC7r1YTTSUUh1r
4rzCDFb+S7ljX0IaYUzadfXPFxfCS+veVeAtS/z67qPqXP/j5xac+4wU+UiZECTI
rDmHlAoFgiiDLvAyfqZ3mqCvBvRYHJiPpyPwnoloPCBS+P4ZPUjxk0Priwr9tWh0
qXnXytAbpYi5tGZU4WKmwNdVbABUWBzEeo+ipF31uCses92b5Ql3uZyU2FljGByC
L/QJQL9X3hqB2eBTet2zdzmA+ONj5AjQOYc4vzbUPcyDTwHc38r7qxQJtWpETm/j
u5fwRIoggk/kKm8qGokRIc63HpTA+9WYxD6aw122vGk6F4gp+KaEsuybmHoEhwTD
IV7Pt8+/nauw7urVhZqnWiK5gm73HGHL0ScnuToGmWpmZfv1zDaXa4cNCU6p8yFl
Z7AnAGhPPjyx1gECLDlTtSBeNw+b104ZqEFCnKU2+MFTWqHWhpI7FFX1e2ALNCKc
feAAnwit9dG9RGnTSbNmMmpSaMOdDVEu3I+6ZghqHzwwI3szwGWGlH2N0+xboeih
HmNPhXlnbzs3W+lYMp0aQx+qvuAmNbhg6N0pUbFDTbhfzF57m1nAgoCSftw9cQX5
KWPt6o0FrhIyeKZtcEe0h0BGB/8hxcEAWKCDFlN1nBAC5zxEevA0/trn1apuhbkH
zqiAy0cWKakRPR/2crw3BJPxdKe66DxwzQY8huF2U4Tlqum4KxJHN6XMDEzVaief
bgkWqk6VE4YwY2sDK9FBvYYODuPuAdyYQ47LfacPkOqFLdzbGyQUyvxQZrUFCY3/
yq+tupuZEkNYgA6nn/BxZGyFXCPNfp83WaFHX8O5AjNlbLt6h5dphkTv7BwDIbZf
DZLfIB++P9pOdne1ZveVX6Sqck9GxV58CSRM35y/nst2NEcypS+nUAvIolIxDrOP
jqZb2ch8Ti4+K//7SPlbwLoe3+hVM0yEMaXhCxY+atnGpzqxZU8IFtTAUiSR5Cwh
jLPGDeK2g7ZEm4tc/3oT4aj+8bpp26qmS7WQUcsDlrNZxN8izcdP9BgXVojZ8Izp
qQqtvJD1q4qySJrY3NE1FLzmGnAW6fzzGixZG2pqikcgi/pA1AqDp0DcKPi5FhLW
QxbBbORc2Oe2Bor/GWiGup0W/uVBnhfp0zhS0cDIwj+3yWTJSUBB0MQTBMMc4YWh
+HC9d95F5KGFIi8HeSU2qJ7909u/P2mmxwc5DpRqunWfziYb+g90i2Gq2I2Qvasc
oGdEItfWrwqmazTBu6bJm0tvIL4+zb7oODHgRJ1lTrel8qJ2573/Z3Mfnd6hu8oM
8RtV+UMCo+OkXCDr+Odb95Ekx3FyQUgF9TtFywNEPbv1YpVUmWw/JzLXdE+nhi20
DnNmEN9P6sxAyQfPoFcUzvDuV1AnmwwQEGckuWTDQ1Fd7PEI5srdJx7Ugvs732ad
7enUAT+3bINdgmsoG5ccDsBKT8Q8qqhGFROVbR7a1m6UHQ3QCucTzYGFS5sWgw5w
vxZ2rtdjNg03GdVPN0aAII9xNSik5VfziG3qxHTd+elfIgf0ivqnySm+2ooGk4oJ
VDSxaYm2UCd7R+0PMoWOzik5cXI4FEgwR624pCt+WSWPZewutRkVKF3QN7CqmFnO
EFd2oh7M8jYWppb/Zbua1Z+HRbEJED6hFkneloF7g8A1KvLCvBOGufc5smM5fI/h
`protect END_PROTECTED
