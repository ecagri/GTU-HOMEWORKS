`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wwz+leqQKlqRfh29V1DV5HJN2SlLSWUvsaI0o27A/iKMlWcUEiSK+tNZVrGM4ypg
mY41d3eX8N/qMLupNnrOge6pPJsLXGlWnUbEZfmiXUy8i6kDoeQDruTzPf9tLovS
p71avvER6WlztaJcyGlZLmr6KLniR/rUmberatqM1eXhAm/zLJxr8Y8DO/Mo5JWV
Koz0q40lLVGWNT6+87Gf+y16udO5Ons7+DGEnl6iaRogaRL5j6/NOHA/FaWtFufg
5Sy3uGXQFK+210GazNZiIKTQgpNWURDyBbeV05KGIf69fJ/DsxbMex7QDsXPgJvb
LBmW3hOPI/7lE+BOmOmA5S1q+0zih9q7m+zXSclx8jI6aOR1+F10ZQ56TEiWVWFY
9z0irxj/NVl6ahpWZV7Jm2FCUmeUnRySkHIp6uVFn9jKj+6kcE9SbD3RqT242zO9
tlZCiEnV1qlqAFZ3JZMSihuDnBucqBh6oQhfNfk1ArDx88WUALV1L6Ifltelk+O/
bSvSb1SDfmwAPJnRtuPwipwt+MqOPR6lHe61iSubR2oXSpeEW9DmpVHs+tdrjAfc
1TXnoaSdX4uBriwhWV/XqA4jkmmITzmjos+FA4cV1hwnJrNhzIuAR5GJ3Pjk3MBv
lG1T5OvBRuJk+bG90vSh7RWWa/WuRKNrVWdOgHTHjQ3SepXj7NhGCo6zBEU28d8b
1RuBxIQTxyqoGSoclVESbOlCbDA9UYTO3VKEQAhBU6GppJfBXGXQMPEmB4Rtgwrw
RA1k24xJKpVTjBE1VE0gvXcQKhdwiMRso6RKxtr7IqJ2J4mHVcMTG2lPsydoD7Kz
TAatog3Jjdjpkf9TyQbOIkQes5iq6fWfW0M91/TGLa1psNsTLiWqC6+w89yCvE1N
SB4SIYtKLQWAQKYTHcob4yFqQqerQTDCv8wqyeuH15gIC+WBHK/jEyguijeY7kbN
VuFrTjR6ib6B0Ibfvis7W5S1Apz84cXIStb4u1LeLV1o4fMWRrjXEF135BT9VHF8
lKQ1naNT6pi28cBZee1SiWFWROSte+szNrRa/w8HOomWb5gPVMV3Uo/ZwSzfeyrC
zUt8QJvzh8+Hwxh9yX/d04D/0NgG3H2BzmVYxnD8uVn5EkoePtdU5xjzXp/zl4o/
rgVBAJSLuBOoxhHDTUrVPONK9TVMH8VYqRXUNV0nVqlll5Lqxr3Cw0fDZYjincQ5
uUxmJMvfIvIbTgfIRzUeBu3YHx5bDnfTgu+N1tbfKKBTax86agXX62gaELmxaS8y
fMa9LA2wBQU6mnFCzZtvWtHSa8iEs+fU4pp3l3G47NEH4CgjUVpm5CcHGsUDHtip
tXhOZw3qm/2E0GpjmNyDgFTrfK3wN0UE91zhEXBp9eJ8DNbP9Ug+7Y7aiZ7qmbOy
j6AounlxfpU46Hj5TTG8nPcsaefOSyLe870DeY4J+KQrxpWxaiGZVV39R8yN1OMC
l9D05eLJ5PtLjUxGTbgXQIdBmrN9aI1CkwIjsPIhmm5uYu7mC3zqcGeR+M2TGpF2
uEALtHizSm3irRHBT5kx/gRk4eNUGz1aNI8B4fyXdW0SOunIYZXqtyKxFIAgjui8
9jq82gKyDi7nwxDD1UdENtdmoqx6nSjh9gj/8kR0BfiaWKi6YcfLzFh0FDUgIO6B
Khy9HrYpn9YcJ2q04sYjBp1wwyhLp4dxBNbFFiwEZRXY9Ls+GA8Ja3Eb9v+N4Gdg
+kT1qcYS6TTTXMz/oIKVFxcJtSOPe4litWmUcpVc3q1BrB8DSH7G27QO9gKRZpZB
70121E7bMgbUhZ2ipTGeMn4iMOqOu+TuUQdMIHZ8tohYNT3Dh1QTg3deFitUPZQ3
hsq+cz1R1s569tHEy65TYRlPfMpIb4M1XSkjz6zZ3trqi4owxYyx4YrFeSyXr6GL
uQJbhyDCtckOkfVJ6swG7W+dT1D2TwUhH/v+TD4Z/2LxrMN7NbzBNpzuWyXNr4xr
BoVcUJXtXhKMyI+ew5XmSizjU5ca33I/7EXxGY1q+cghAFGqxaNqxQTcZfIiaaif
2rrpJ9QzG/Mx2tg8JeMb97aIrWXb4ETGhA2yaeCmpAOrFdbLUvF66blKLZz5yhGp
4Z3nISWtqiW30cO1/ODSabLSCRvKTqEziQ5yzD3tZi5+BhSifqN8sahx445+AhNe
1IQgM+xt0+5bY49ubUtK1vOYqZEbflyHujFzjszjjCjmontVA+9Y8nTmazw+TMbt
/9vamYv0WElEdZ/e1cvnPdD5GDxhU6EfFzrqIlEb5QRFyUMe5jPlD21eRVpi5kFs
fvSWELpK5gEnNmJOkD2MiJcUbu/T6ejy1Ck9BDihNA+jeDI5FHfQ2adwzs+5A57A
eiiN8mEN/6cf7Lb/14C0olSLFVUGDx2Jsn4f1M2zFmS2GBrKpsgLjsCRwXc6+p7F
YrEP8pADc3ZylwhusPKerw==
`protect END_PROTECTED
