`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gz2NNdCwBUDxQw9QLX1Ku8rZP+OtKkYT6FUpL3ngHo4bV1fO1E/pj4bbHNE7HKJq
3+lySHZBVmNQ9BZYXoMNwH+hkV1kleHar25tfsT7Zb+uXvUM2Nw+ux7Fi7N+srr3
CO9eAQi+DaWFLQ8JRPQURPJ+OUcDivK12okiZ0y/3G5DI/2VBY8bUq+9iykEV++Q
QNlRAzMDi/TPPKgW41CNoY+1au7e/ginTT+0eh7rEqKKoGEzI6/e1mzQwmXRqAw0
K3qsi4bpV9jxoHZtfvcXg2pBJH3v0i0xYuMoOupmJ9KjSwzXVBPB8cAHSAj4+uF9
ZeKiVf8BVHEk+N5GWCFm3Sq7+IJzyZLwfdWu+86qzDzWxpBO7T3rUi/+NMjTkhgA
kmfAZ/Daw8H+344Ix+2H+GOr0ls9Y/JZYOABWbVQ4BMj8W3cGUd3qbNGzRPY8r2T
Mq4WY9klxv5rJlhLcdEAgBrwoioyDmMzfVOq8hv5/8NVGBzdj1OXH4Sm6TZ5IvOc
Y7cGpsg6bJVdesfRgZnshSYYfJi/d95NilidT946lx3LF5Cd59IjgphO73V70zYm
jcHT9WoJRN6Zv8mysKXMrmZMNiUtAPJZFZlMuZVD0hXMu4lzlvmZNcBAR5DanGhP
q82WzeMSY4ZaXOh9QcFB0/fLRXhT8ZJ6Ke/XspxvjRce8MLG9i+ny7U+/XmZdwMg
W79IcRzYAOy6gFCf/rIjWB2dukS3T7sOrVyuGyoXj02DGVtVAIkS9yG+4xT0fHpu
LGWnBTpUl3stUM1UBwviVrZsMt65dY5a82myuq1oqN8wVV8dIwKx20w0RHZaenuL
Bmh42l2khgCY0+TmpNF1UmszboXT83FdZbvzrXmaoPZykUDq1fH5+g+8mlCS6X0n
Z+mu3n/73rZLrJELjGngpODsjqj/1pHFHt5aaUlrDWTVrhhAJ1AKrfKmGpJga3Sx
hiMhBAPb5X+DDRFX3bbHSOUqfEnmLZhaLuNBLi4qTaIadv5StDqgulmD0y5RqgV9
FcrT6J65no6JpcQwEMt8mmqbMXXLMT9pB0TYIHX2pHIr+mbjZye8FkTGuU8SzOgT
h2eNyfkj8MHYeEgPw48i+zCZipj6wJJkF3e3x39OwLv/tOyrjGn4qpadGDh+mePG
JsqqZjxAXywM5DcyNzEZgiLU6cZ15fcOD14Xd8wyKSv3OiZZnG57UJ7udmhV2gZh
8cA0HpFw4FPoj97vOq2HFT7bOs2ry1O9+9RFTxd++OIQBVYDMbw+WzZMPVfi1woo
8XX+tAZj7CDapMCzEk8/6ecte1wnltr8lgGYcA7NLMpUhH5VEqSHf/xh4y5PSCzh
PqQ4V6p/FpDA937zMMOj5Ezakz8Ay+l1wvhlio4MfhF3CPH8SUDAzxXsMu2Ukh/U
nCQ9xmHuJd4mx7GSKDkS0e9kZ4iaDPlMBnOvfFGiyfQRBrTgyEd1zNLyIMktG6aN
6wyrlj84mpUYvE5NZi2NnNKq5kvvLesAY1z6KFTY8YE5Ob9bMkKEk+ovaQYFIGlJ
/OHXuChTHU2ypxv8O+cM+gZnPWnDwFnBdTO23R6uz87U6wtEOXBcsJtkKflTYFrV
G2+BHoRojCTB7tfonULsj9zLkqpPNZ2HRhIfi7UjgjR4cYehEZndMk6zmO/ChJRA
tqAsu2URaQZwCz7rSmpP479BWe4gVFKU95Ql+g7mpKHUMDzKIWWeaZxvVbba53mB
A3LJpKQRMCycTSOVTLtNABuz9MSCjnrQ7GTwBa1pAkcXD/pmzipsqoyRgXwIL5wY
XDfmfgRDbKC/WHX9+nSK+mA1CFzO7cRrzCNUXhh7/uIKeQ4MceZaHjZpvT9d1xrb
7ZJxptb85ETeQsZLhrJec5bcc7FnrdJaCx4c88MtUWickklHI086+0urWnHWswxZ
sZ2kns8Y+nK/dJqm0SXCX/GQ8vdBsrqQB9OAlThJTclp1QdGKPYCm5rpIn5BhPSA
iwO51Y0n+1UsfsfIMrJWtxXJEgAVcy2FRA5RwdXLJ3cWMhE4tSxMPKMPkWaYpMUi
08JlUXAaFF8dqTzC98GMK63oAh0PIHdkaHhS8jOW8ORlDxubUaSsUDVBsQsCXypY
Pew8n9IeWiKARhr4lpRpjWNGA9mXOSluiI6g6IHpdD/jlDwZdqe+ehI4FOEBoXAR
TgNnB+2HoPuNiocF/Z1jFnu5lBYAcoLjifrxeFFAa/p3j4UQMReMxnOGBY/8nC4y
tNVgfgA5mYUvcfF/Cy/b1kLgMgOpi6SfUxRFyKCjx8hxTHKI2DtJ3LjalBsk1vXR
1hzonzW9fkMKfG+DjZZxkbynDyDrUK8SyjKnGmdY1TSW4xwfsZmqOc2RvLmNmEL2
yRTGrmUqeThJtQQOW2g8Qr4z9cr462M82CNXgW2uR9Q=
`protect END_PROTECTED
