`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C5j8bOzK5GKrFKYICUbVPnaV7xQkp9zA/C9T1Y99XXS0BRP4nSOul6oFMLcsm6B0
xXdIMz4ZfD3TGk+Z7WXZKE2ZaztpmiLzjfmfM6C6Fl07nyM96m2zJ5CpvxmUw7gK
DbvpK41tEYqtbPHgqEX7snXyU7pj61SrXqWooOhs6PlQPSqo0AMzM12SXCrzW72M
iUdniVrBLYB+1SgQr9SOHxJoB+6abdMYYOMwx2QhFE/45CxjmQjOZpxQikmlaOZI
mTA8ip5rFr6AaYcXIaHrbnFMOu7JpjQMnhNudxkkD49Wz6LNd1LFkuNaveaN9QeM
yDeN/K0nVyjI693jDFuBLrpZACemrx+qNuzJTmqnsvs65vcRNSsfTCVeeDnhPzt+
lipRkwEkxcWikb4No7yCxlf08M30sLAuzHBn/ng0Oi8wzQEDpXdqik4+nF+xzHp9
B7fzrgXsvvoXNhkTFFMF/ZW1wqVDk/F33VuTG5efsi1sj1JqQu35ToxxUheWrsx6
1q9bsnJP6Q/LuoZLon8S+2bHZJ9rQUenAV+NHNzY4ux0rm3P/9a20u4S/GFNdcQC
DZSMHRMRwPI7+C5gpHGBU0MJgKsEu0Q1OCtlZmohdcvv6fdkj7qVA3QhsTM3Eh+t
fM3JUYWw0H/Pgd7WNn2KIsGa/Ta/vdavAhu5PLGxc2T0KyNVUow0e1ic99uvDWUD
fekmcgFw5RqwdtO9bwOrg/pJ4ruxYlc7uSyZSw4Ot0kFmsZ0kzLvwvj0WuxUazAk
5FRd7JeHataID5zED3GweE7koUavzYEnYEk0jtmMcfRn3IAmUyOBtMiwpcioa64x
Luuh21kX0PyQgkiXU1svVf1tqsGpFSLTCQMAA2HaHkFdoXX3xvteSs5oUBVjDYfc
d+rCL3GdyDMEUvrQjJbF9F2vzIDgXbXcHqPmIbJHrQh7Ch2gnNezT8qceXfGVnz9
cLHimS8munog6xNSv0FVMV97mGfXr5az9cAojOxiyvHBPm3WXGKr2xOWxZH4UBkr
TQ+CMpPvCd47ty6AQ98NwVNwmK3w7hc4zi1dQLIkV7NMqRwABXD+BhkJGGTnj+pZ
q31R0xynn70ZA3iFnMeX4LMQdTvCtSmzjqbgIujymIo2qbyHo31z2+vGtZTpeaxF
tZkdAg8CE6Z1stEDy//SbPz37CVlTfjYv/Ldl7M0CJjGTrwDL9vhxkfi/dc4dXIW
AldVLjvC2ApM0nn8hqthFmLuXzuiS72nyTFpWI1dfprGVcRqCTpZmoBvLmF1oonf
/wen42QO8l6mfwh86sonTpLTUrZd5C7/RKBuKCOGUX40rQuZUIV9q6XrsybKCGOR
FCaPtR5FClXgpSG2ZHira74GmQFPLE3ykbsetrlcMGXSwqNAOAf5wx+vX0RLRjxN
vq2trXUUAUD4fi7eKZq5BmYvyagTg3W/h0b0E6CS88Dm8FTT6cP511FpEs+nkEml
`protect END_PROTECTED
