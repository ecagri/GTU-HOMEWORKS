`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kg8W1wVLjJIuxL3Lwd2KXju53moo9xBFrJIsxKS4nJ0fC5rqIPG2KF8UUcOulzXn
BprED2fdjse08oJSJKq/qf9/WgLjA88pP3ksu3ddoYlxOfmQXXTlW/6xsP94A7mn
VNX99W3JmbuLyJQtBXcneW2T34T7/miYJyUYnJJPlhPvfFGnJpc52LfWHFANLjFV
391fknM1/iD/6PPZ3UM5yFDGv10RirQ+BKs3f2N7rGgzs+zajA/TxAYLDhnFU4Qk
VEIViGfZP29Pdd1nWYKEh8RJ33wzzsnvbLKBTGvCAKTy7ZHMIB/PgSmZ/jWXpmBz
VfxVb3FW9FhKvq7oD3AI9htQhtX2f7178uJP/GnDikpRSgEZii2LgyPhVViHMLsH
0u0sf8pRXWDPGP3NQ8P+bgZMabRwhlaHVt2gqSDapU4s5FzM3KA3OBDLo2MDAU0U
vbT4YUKtMKo7yd7dXIJ17Fif8M2+XTs618bIqTq/ybsGA0y5jyuL6AypBZD7Mt+v
/Vi7Z4s1iG4/zKfEutPT+CSmeuvPdAd1BbcvLbdGvJmmRAmj6a2OT2EeYxg302x3
R2fqR7KBf4sd/O+rtwoV0leM5DBItViJLkCxEHr/2SrwEqxRTk6WBIEi/LSz6bXo
FaUTWhjmZYeSJnVZs8UYo6AVe/88QAK8PCwg6C/ggUd+7z1XDKZWClhD8WWFS5lC
CV2Okn/iA7n7GUP7DgaqezqcBztQhDZHK94+AQqla7P2eTIHd9sS6cK5xtYtDdMs
VJVgsbKc+yNONL3ybJMEqNsLNctE5C65geCE7Kxp96LwbA7YS8h/4oVe9kBYJKWx
Zbh7RTf/SLv6ABL0Qsi4GHsSQUHeZZEAuL3OGLb3m9UdqWqdL4nDbOcjZCMhEwv6
3cVxGY8WdtRpIo3lhoQ2bSji01TR5YojAm0r08rRlr6FA7Sq7MQ1ozQWSCFRVl35
`protect END_PROTECTED
