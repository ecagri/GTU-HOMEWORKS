`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ExYU6x3d9YxCGMwGS+FHCfNlEP5z7GjFyEmVF90maSII3/qXgMYTDk37PXECd9pG
wQq5eVdGach8ad3e184EhTU6M6+VogHn5DP6R2XXnYQQU4cGRzqaavwcJzm8URBM
Ce3WcwNZvfgUaQ1RaDTvpT8NMWnzfkTOU32hvrSwJcABtautjrTwRon4vn/XSZLP
brlnmSaxUMD0ptglwz1LcSArLliBR47PRPfymZYdSmJ9EeSOaP5bla9Gts6+1OUS
J3pfhqExuCsubtNvygDuKa0Xd46nabfs7FQ4e1AohzQu2jHlnPL+Iyg9hp1Xfuog
6DUYVhQRUAsuuiw7QIwC1q2vpFSKLCgCcdkg4Hv1oOU8SWsJQLeLrBJIkK2I+FSG
55I145A5vJWBrMP+Ilr+QSnGwaNKNLZ9BDndpMM5cXNCV+hbXYsF7ROK//HtfD77
mZUy/+m0NALdBq/2Bndchw/H/J6EqEqubvO26qj3eEIVjUp3mDAgPdB1k3VRYitq
VexxlKjRgfxNTp5H82LwdIRUOMFtgs3fxy7hN7sWFx2RcnCtfq0Pp6CJ8TCGBea/
gKNIw0SmQWyhkVDzXfOswg==
`protect END_PROTECTED
