`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gr38JpeCUqA2kIfmZx6OEe0kMo2mCcFvbnJlrtK31VjaVu9os3hvs6pF0PvrzbXD
Zv/tU17eicc1/FuAXmekaIiMaltM1aGUsTaNJi6sEE3afiajfEvPGYchI5p0lv7K
lFKZ6U0t61RYqEZ/D0nYF42zyX4GDGRan0sA7z+6lTHwenKNOLG0wb7R3nTT3vEg
j3QafaV5sj3n5FZ7Vrd9yMpj5ksUCp9DYedsD6pljKCxra+75vFFeOovjiholx1r
OOXb/wy5qnxh/ao5rnjUYdBa4Pg/vsxTMI4gaHnPmVswWm7jcS/aCqqZTl9q5+XH
1aJ7jr6gPi0ajl3ckEZspbJLprP+TAYZStRmeEmiI7BayR27ceSDDzh/8fp2YoA2
AxAsXyGG7GcCJQnJs5RjLhNXH+P8PZ5ydRy480bX9I39Bm05Mjosh96kWtMEKG0X
FLhnGffsjucBo5sRUEQWz8A14z/13avYiUQGNpIGyLSOLnAbV67RjKwuzENxQhXV
gtJhSy93iSPit66nGpp+Wigb46Qq5S7iRBfTKiLv58ZO4S6tNMrf2iJI4x4zTPsR
vKLkGFvERoJ9K2cFmXHxjG1XCH7hmLrRmPAeDveFb2lEkykcVQvIj96oFoCo2/S8
8muKsN2MH/XZivJ6rGnHnCketnmqQrvlSBU0K5Meg9E5JtOR7p7CDvxbLDBRl5zC
`protect END_PROTECTED
