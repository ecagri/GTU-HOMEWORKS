`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pDzc30GtiNfjt7qstxV0mS0RYqIX5fL75ahZ89bvQ87uoGbwPsdUEk65moetKN02
d72RjpLyNTUBjCm70hh1xjWEOxa1MpdMxynYPdXMtIQ3BtHFyVbI7136JlGzHw6N
KSxFcFR9mTayaRYud+hDo83vA8cCijm6LBTfzawqWvieXgC4d1W7B8sCMYBOmHwb
96tfzAVIfi11BawIg+LPgAw8CvjbzhIq7lSOExbEONAwo9QUrN9ZnGG80Vna0Haa
3uCzp1NdMox8gY4xtZCSigK1vF+mnkCzs56T53dvrvVyEYZzLl/PIXTSN4XEeY65
IZVSXRm0iqMlvvNhQZig5PklI3nYNuZ1yo9ivUh0ei+xnV34/CvInHoMsARXfiXh
8CpWGBaS0IM/0diaihrFXSiORjfhqV4lFVKSQZfEoP50gZGR/C1k4IPlZUwowOVJ
QWwwWqif0k35bXYzwqyH/uXTQTBkCe8He7pD+9Tf8P74GWtfjI1/QfgSW8Tk5qyi
heJEiCnrfefLASLH95VoZWyXdt0KSSXN2o8JVIOcoSO90IlNriniAe/Buw1T2WI/
IFKmPPtKto3MCiXFIuKKxnrK+DOxGWIo5gQNfW23ZbDgGwqu33ljtckH71xRQmcW
O7aNdDVwapvsJHRbqSak7OswzdUkBQthGg9APVhz1evgqnBo9EYPzBP/tPTS7MhC
QKgRgAbr/og1cU4kbITk8RHzUCfg2j+e/sat/xyHcJIne02IDrDEFVSmksaQL0ik
QEppPpDj4hJCPl+cbUYoY1hg1/2rPopBTjSCNlkQ+Krjs70tMbL1V+fJBwMw1CQg
G+DskNjuktrny7L1Et1ztxXSm+36OOqytMUUnAcoht6uttLLXvtjV/ujTO6fPtz0
ei3qb05DHmYYLeLaoxixJVgph22stAR5ZQFcureyG5Yrqa7dTP1NBc8U0xtRqbYY
PO2eBGWu4FRwP4kSPBZEOrNDyRkCMwJJSvieQei7g1VNxRBKZfOkeXMJEU61l+kl
sBTTFz3TH8Cjfr01VBfkIBd39C5uyk12/AxnXrDQuAosdYo3SZ9LFEpR4IQvk7AN
is41urfvcB0b8UHewL5jl2a7/5yHFrHtlQhDLQT1R3XA8vJ47gB2w8W/iIycoEys
tiej6FTMyW1FBusmcLKywmltJVWHDJsa4K+JNC3Tp86+IjGKsYsZivmtMMwyC2gh
SnoaBp9CNOnt6pQEiK4fn5tU5K6CpfbhA7TqjFxlXmNTz48ZkGqsbvuGHq0m7+uU
aAYqn5pNXoHC3LKsF0z+TLdCLH9r5JDnP4QTUclZP6M=
`protect END_PROTECTED
