`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M3Cl0XbL0qpYW20R4X7mF2LX1tYLPt9g+7DB8p6o3NzBlJRDQlf3cVH5jTyId+oW
VlOnjkGwmKrn2QtpGXUokbRfF4lB/xPfYX3gS/rNaOQRPgkq4w+ZhDZX343i55Sa
gRDbe3tIswyykNYkflszAtro52A0ig4IA+sdnQo/pTuCihj+P918A/vO55m6r8sC
tgtE/Q0A6uro6q5PnF5HdnxqgGIYbzi9bzoCzystQZQdCKbbi3iKmgFtReGWA7jp
8YVQ+bEUc9h5qX/CNlw4/pkS6G/xK+grZLA64YPVXNH9qOoFk7UqhTFlCieQ864+
pxXKmDXu7eSkJN5wz3lWcQZ32gm4RI03fhRi4efmUWl+wiV8UHUlcPG+96vwQcI2
PRSxjK04uoT8LGXDPexSAnW9705L7WZsOEj9iSxt0I8mZGGKz5Oc00f7GI8u3yxW
yUaNd174oGF+Y4xX118hlfQRJVZyIstt0Szfjw6TLBSwKD1isXIfGpK2mtRiC8Zx
LIt6GkFHSrJHW4xZ3YUK61kruGtUSuy8ZDnVOUIkuM5YR3/2nNI340FIJNqdQsDk
02IwWmaKLBRK0wynBPy6IRpvEQkr6NMjEPjpxTSNf5peRuXQIlXRvlJbpiVya1ih
rcDActyndzMDDmRYeHy+Autg4xzYzxXH3LSltP5MW0bpT6xQ31rcis62NaO1gOaX
4lyZV+OYShhK/nbl4m2PZcHDIbobnJMw+X03PBW61Q/RZX8FA8A+e+vM5MLkv55G
SFecgMFHV5UlfwQeGWYbwcRTiF6hgIHP3P1ssZF+R7r/l8C9Ww5U6ca7DOzErygB
+sM+T5iAlKnbxwNZrZk69s67v/rZXy3iDjuZv5QCYcqY4aM5z3Oc7ZZnjC8VxNUG
eY5vKKptsI9PbrmGTGyYxRpacyTW9JFmkoQFExtHC0fR0SIucrNMDOKtRpK0H88S
77xRi6gMhNgYJXrj6CMOoZIUGBtCwhbk+/PC2gupmuEtV9JEnDuBAJgCh+aHut/4
efdGIXmj49gTNeOnVFxtRkmG1lxWsj1duqy1r5Tese5nyec3dju46ljMR2SR4ZRg
4h3F0Y93ABe9ZslRzMPVSSyREd615egwcH8HzI8cSRTa2oBZtg2oOzWrU1s1sRJB
9Ls6NIRlQ11+j43pEDKasP3LnuiyJK+JEhpYt5MoQOn4UXgv8AF+rcBxuAvA5mk4
Dp9JyhD0CWSYvcYQ1faCF/JD6KETStM4ZylfpXZLaiGI+zCRO+t8Zdcwgy0eeH1Z
pyWcwk2u/4uD2YfXZG8rV3b6+LGk9MYo7FAE3PfLL9FPJv43t1TvipOXQjE/3PvM
Gjc9vhOyGLvijcTbaVyneaXg/WzZ41WGeUvEHQMafzqzf7GG8BgVAnlU4G+ey58M
aBBTH00H1JHpLGFOtTTlb3Pr0enONaZ5mMPv2DEc3hD9pBjIuUlxzDLEoY/PYO8o
2G3DaZVYhl8xsao6cEfVxhi171QwMa3gX79G/NcEmiMC1eJB6dl/jUdnDXy2DA29
2Nld1UxsuWpJyd5/BxXFOkU/zSrIIOjY7NqIe2R8ligysRI/5EMkd+QGX0z3RJ5j
7obpPwgC+Yax2NRotWFC7N6Ut2R8SEj/1GuCA9PGi3E9mOVPJl8zDbdH2ypR/05i
NDmi/mCLgb4ocifS5GfSTgipBJ00irQDs33qzQTVPxndcSlAckn+TPmBihAGC2I0
boivOegyqYJ1K88MV+DOVC7XXyC0kodC1IVaf55kqNC+0EYVqTNn++UR5pgIwE6F
rtkhKuCRy67jWjd83NXesTqBjlNRfjM7JDPZ+S94Rs5Uk8HrEewuLdCPjFcVaKHm
drq7C43C5W0/LEK3/VHuZu8Cwr5fl7zGlrR3+iui35PKSzw9kIQlTXQwlDcqf1dU
9D4z9J/KsFN/SojzqFqtD9KLDIvSgMd6iX0Z+1LI0vDzrHs0cwVom2GM/uZq9ITv
jjHWlScKYEhQUXomLQSIfmIAQDT5qFub5/bjoDCcJrl0Z8Ww23NlFCFKKAXom1Wy
I9aDIzTUxXakVvQ4FS0Dj0N9NrL25kqn/FnjrgUdGkEfYnglfAzk+kN5L4FVxcLk
`protect END_PROTECTED
