`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YZloC85GUYgHRl+YzFLxGmhrQSnCK6j+3geANHOBI5NzibEu5LER1vSLNMtPR+bu
HUzDhg6VRcx4ZC0nl0PTf8IYHWvo41Z12BSRSrZgESmEs4VaU5vJ1KMg1IkW2GVB
ovXXXEFWiTqNPbi61eGWiUgO2TKNjE4wjLW6+ENUndqOKt3QBxTfUM3YkAsH821b
KLj3f9mqf3qXYZVceVDkqibiA0r7ztRPIyT4bzIfqwSW/+pNR9S0OV2KDJAz/kKf
1Bd2rDB184+21s0cIX4TSXskFUJGg0H22KMRysBrBnUSHD5nuCM7Iqm8L5bIPg7H
b5IcKGocLBNzQt0P9BuE64k/yZAliNLbxpYDoTp3Cn63zueFngZlJsHrKNGWANa8
lXJk3i6+AKYT/HT42XhBdLCgUeYgBEy70JrBy1n9KjYduBGFfxL8FhgvWY5kgMWg
QL15xLyfqGCTyPgkdkKH6d3Rn59X0aOS0ym2O35IAMviZd5OqZlUY8CpsOIwqNfr
iZ6M9tz3c1N3qOgizKmHMKZ7uOu4VMJ8/9dt52ThX/JOw01SfXhyGHGFLi9AxGhT
ePzXZPO/QTDEXBtzy2FJe9GyQqjkXYr+9H7yJEM7/fz/CcswKRQTfWE2McgKlC/d
E8dNAvk1uTqVxyia6Ni2w3x3Itzak/svGscr/CFVAPdL6AqTl9zcjnw+w1hcgIW5
JcrCzEZfdNjryjVE/LcEX82xF/y5kK5IgJneLGro/uRRzg7HESLBr0r2+g+xnktn
HJ4fQKH5pAYtt37kkE/zvhv/vFPNPOstqePCYUK8IIGW5NNW08r+XGcg+ifTGgZn
LOOk8DLPliSFPm6NslJngptmHH5yqkjBfjeeivHXmM71brPC7p5oFhextRbdgRnF
DcD2SPPg6vtonxgRQJU3CnyMMgq+xjr5bjYz0rjrhxnNQAHZyLDJ4CTaDcyeInhG
TQSLIGDNkFcPONlvi4mNgR8WvFCkQjp6HejEmyWsDlGivyZpm/BT3EK0GESssdUw
YLoNFH5lg0wn9b3WFVzig9TVeNR0HAmerq60ZPEHJVEXbVde+Mgunj+yErXKlRm8
qrEpFP8vy2VvhtQynq3t0SKoQvwpcEtJHUafQGcq5KAaao8d4ysj1Dwl2Hg4R1G0
rkFL0eov3bNw1Wqort4NuKJCIT48zAqNRTd5DTHt9KaYWh3M3Az/hyrDR4KXLZbk
S2X5bzmWx+qdt78UCph1TG+tFQDVULy/S4QqUNE0iMQaJ5+TkuBE1XoPIx7KP7yZ
6Laivic/CCfLVsp8/zprFmokiz0JvLihBFKz7B2O8RaRdE0XCkx2GAxVtROGQE7M
55fwnV//8SAw9kAAXrnt8TrlbI+gkh4p8q82Zfw281oKeEP7TP+yph5/plVTdHdc
hZvynMHuFWoDdBwotvR7DQe/EP5bzQ3ts8VzZr26GwbF3vq0V6mv+0j+imwk02Uq
+XdvMqm6K8I9JFIK1/Jlsc7JYypj0zh25EehVvARS99Nmrebwu+Pg84D5bOVuFzC
HEkEx0kQ3Ugi04CTqfVzLYxuL+TAQiUqx3TpT6hzlLYxMroKGaygpdiL91UpNokz
ETQ0C3CImqdOX/N11tBwtFkM7ZXEloExwmTNc+OfPVlstXs+ZTcfx6WbIuxnd2DZ
HLlppNssdJggUgoav87oTUZsvRZOvIbwCLIaqljvddrNQZdj7aiUIF2R2ExytDQs
rKiL7ucjNNY6SfmXu7ilJVj4xEYvKtvQZY36TYZWS1lS1TcCdUmoK0hVL6ixdV7+
xzDrHLGer2FGkxZSXDecJ0elmvFwjDu4JtM9ygE5u6xcxRSsT259YVmfvs/wyxRA
nPUgxYZyw/A2BeNCUg611a8S+JWmwMJmhKCZMN0FJHOS8DzzInb125vMl6GLV+Tj
PEe99PtmFdwtWSxkMrmRwU7x6X9N81cYQbM9enQAD2OvBYY/Kh76zdyuXJzhclxL
6EKLbogAhmfVxkOwSuOhBKYjT5I9vAnbfvMtcNwNhMcBc6217VZbIqXkIARifllI
vCdF4g85m6jVie6UU9qe6iURAGuoNZt4Sgi/0Oh4WzW3hFQ0rDOlFcZ+YwZ8dyog
wcR0B6ZN60iWW1vci8vcU2UQviISQW+enH2eUWEVK8Ctk6A4Y2qjKsi9dA9AS13W
15xHlSjfnY80dAJNcH4AIeWCe5IbEgZs1SVYc1IakdlCC4j5hrULVOxTG8rC1YCW
HZFNerdNqG24ewMgzbw6NmBWUp5QiN8zCosjCfT1dXN4Sy0z2L5wpOlyJfeql2P1
2gbyKJ97DGzpZtvTrRe0JfF3SQD30xdraTocs30HJ5YHKr55c2fLkJlzfBb11zkP
vKqNES0uAuoJcj3tiE4pt2TXiwz2rraSRbCCLqJ4r2+bgtRSbwCEYnMFZyqcBST/
wzgdATp4w7oZykdxv91YqnJ6ywiLShxhmFdZqiZAlqwbo03Nv/E9bAZ9vrBtBVEX
UExxjwzUGQQYo+NmFl3TJcN8N1fj5eNAb6dG9wRPR+7HOMyfI5xhJUZHit/ODzh/
Kbvh9aPq/hLs+3iypxjJX+XvjPqjXNh05aRGiBYeVecolV2/php9D5HUjPgL7mj9
Rnuqg6z/KvU5c5EpU+LOGKtG2xjM/Z6Q2EjbmceU6JWnviENB3gRXwVulUBaypNQ
KCJp//XUceQ7ijbqn+mEzoa5GB05bJv8aYBIIxWPPpSweddgvzUTYk0gvjZ8o7qi
hzuMkylG0LeahURNH5c/ZyOY5ylotk/1xJsLgFygxbA1M4JknlZn8I4KLObJ295f
BO6x5dkhcZ1IgHwlG7y2AAOUUVXJd1gOB0q/DWZcBYohclgMj5Te3Xmq7RFH6L89
JcVafEn72mjEQ0eZFiXtKQ3ri84pSFZ6ZGXuGRp7G4AxypmpS+m0lKvPLroHL9gX
pRRsrakTz+RefSWRLtnfZPrN10SAQACGM2RRgcr6Q7I4OuiXjBlNUhH8lohlZgSc
J46/P0kBZ0ypX/ug+6QXD02kegL9nO36BphxUc7Wwn3YzQvXtBVc4HKzHywcuQNe
fn+RYHc8DnYw07cbhrf7mY+7l/Mbd2sZP6I16yi6xe0lU7dNnCWi5eT4Hhwy88YF
Q9k2/6QYCBsicfDhn52xiL9Ko084CE6N/J13q8ZRHwVPBffvYI1NyCUtRmS5f/Nw
6EATHp8eJDtTb8AXq2Y91up1OxWoQwu/0Zi/v9zA8/BXAJtB6Gk6exFcvYfrRRLS
i46VHAZBvt0Rw8+j+a2KXSRx6OcCSkQKlFG2gglsuqREZiTqaFJG/SAhVOuN9qRZ
2g7u4Zbd7sH069ckd8YdFTP4lufQvybi84Hjw8ftvPYhluBhkFzRjCVXIBnc7Vik
AstSM7indef4D2R79Lc49KcDIb7RlkIT0ytsxH2ep4psgx/V0vrd7nqyAW0/mew9
l00zxFU/eFX3yAwtXlecOK3ZQJFWtQeK7rhZ/FZ/K48VncUb0aK6vK8fZ3OIvS1J
ARotff4Hxkf808qdYk4G6N8kGQIpFZ9tbzZXMvipHVsj9YtyXpWjaG+L1p+6PZjP
4Z4uE2h/cuvo9rZPxxE4UHB/YbUw3Uwqp0XZCZuPpBucemQyzDYtMFcZK76fyIl8
kpNnpn6ALFcXcrsAE9oZvJqZMVFJS9XYMLVYjzj3i7vtFSgKHq3wrhLlNSTuGkaD
YCaUQfCIxnnMkVR/RRpZFjDJs/8aTq9sbzJ5DJUy/BOewo0x4TnC0FdQGViJsant
rbGbthjvWj4LzLR1tlCF6mfSuWXLxcm5ib4PB9Y7P0Mbhr3gVJ4QCJziS9ccrAXV
sjtTSUBnDQes4zUy9/IEPmKpmH6jbn1lSiS5M5SUiJcQRrSOxmqIv2jBIDfBQ8GN
85PvX40VXs/XIZBxw1y9k44mssu79HrQ9OzADtUCLOzJJYNXt3ERMr7P4+Zdge6t
EywVFHiZ4uqjchp+wVY8F6wvuLQJ7M2mZ4tuQSCmsyU4SmFv6eCQ8bDYuqLnVIZB
dfAFbCrft9JNKFyzqMSLFEES9sFu9CiG817BUbrCw4pDma97WAe0j7ZWsv4/NsZe
vXwbllMniaYWvNmgOX1If9vj4wgWjHIv09pzcoAjVYHsXx2vEa/gs5x7+jc9tvm5
0us34mZ6laomABHtdG9xOYjL0pssg5szBd5usIDk6Lg5qKdniCHNKkevrKjJ78JJ
vxuzAO6SbZwvkQUEL1WquOA4jPFuLBMAfDI0B0XBg+Zye3zAO7MiF2YtY4XiA21m
xLa3pz+z9gup2dJJFItpAZabtwTr8YZFGdFV83O1N29RqY2v4Tk/ppKtKMBZl88C
OGc29nV2Rcnez4+/ShasqUjtgEj5SbcOYcwMoJWs4qt2SV0DwQyKJs/8X4SYTje8
BGuf09oF0HLxqsPWfDVL6Uy2a+G6waneqLlMfQSd5imHCQJZEAefwfYRbvGFAVSD
6PauQSpiF5BOza3ZSObL/pn1M82u9KqSVH+I0OYG+XRJ1Dhl9x3G+GvbbI4P2360
x0XUV/BwsphtGpqf7+BCf6pdkO03y0ID484+wogITAH2R3GwqZYZ9c88VF9UpBsq
AkI1UoZx3D6nIhitEmVzqW6028pHhgO1xN3SNupCRKYC7U0vqA60YzZXVb76w1zx
NGrdX1DeyV43Vm3NzsBPwfQJoGZY89JXDTfR3Ax4qFuVVc6S8kzJdVfTubI3PXxX
BLp6JnDv8wmFkK/K9ZFN/SzcjWFsiChtgyaZduOEag3mCojsinSiOkclewwYq69M
UeCqFUngt3SIFi1qcjKajKwAPNlUgce7ZT2B3yv4+cEQm5j2Rx32Dn/iLItQXRst
oEYNUSt/2lHN5Yvlg5lIgtslR/NsKrNHHPeIVZyiZtxrOWZL/dfIZx2x/V24OSO0
xVEdEnXXvWOFGWrAhHOTw9b5zJ6IfjYgAR5oqeSQ8NflXz47NETOpM+diaUE0YjU
h2Pf5XHLizA3ESI6zJmZGPijNTnci4DMARXlPTLN1uu6gIKNxQJvD30bqpm6F0MY
Vsmkrf6k6xDjpMlxHpThGCKoN3a33M7kDRL2H/XXW/TLetPpHjc+RyT47MVjVgaJ
HWczCAe5G+e151Wjp/jf9klgjIJQo/t2WRfixMpUq73diW+/UirHsMSlCySC+sBc
i4lawKrGkJEnejDRgM6psptEOsLRkBDW26OTJ35enRt5tDHclXMLqOff+kksRnIs
g8r6zxGIIyJUFirJKhuouWVqSuVzcCsXXgGinl+5cyYxh7BtkvVAW9UCUWMdw+ql
JuQgVuDs+fZQ9V0IZkr3aB26t9XnYBvfOpT1ZHtw4LFJoqW9H+EnXDxHzH5kUqyu
uOXXswUEYKaS4Yz6N6kIJwHMJbO8J72KwuCuRgBDrkBaw1tN2wInGZZRqVTKNs0s
YgJO6DBqmohuQawQE4nVrjZ0WwSJkO+vjJSkEXIehPhpT/PuQ0J9Q+p+g+iITTPn
ZPkkADjPjmPRF0TtNDuAXBKFcULA1hFhteyVh2KUVA1zIcBxoJFqenmEkL/PNR4p
4nr+4QU9EP+PPgklWCYLrcQC0P8scCjfa1iqOR9RpcfclgjqrdJQBb47tPxLIDO2
C1cxRmGkwwn+ijUvwG5kvVya12eFhzk/aUSLuDrXTwWWFO2H0Op991dvMGxx1Bdi
k3FxfhLHGMWi1hDgNAD3cVoidWp62EYHLQHmyICMB8nYwix5UcbB7U6TubN5OizQ
Z0UqInFKTmSPF2Z5F71/415A5nRJsP8kuD90hYhOucklohykCsyCki8ouxKvfWwr
23D9R+2CeppBA4WkK1PKvjG1SYmg3R4ZCjL0y1bFnCyXQkyalau+ZR0pNlmvkUAX
HiUrE19/k+KdZiIyWEtGGDY8egZ0x5rphJYNdY4gYyxxlmYg8sqC+H5HTFRQlEVQ
BnyLHx0y2cyYD6jO2krL9MzuVwNmXEzqoWGtrNjn14zD+UW6TaVkY1YhAFttxqwC
RJ2Erut5NZVeOO1FEb3wE8kPiCRQr+qGEyAlPOHs1WKjiyXpqvyMygb9mPd5JUX+
7ZEGduNmxIVDA24BFv4gZjGTNOidctVi3DpBGGGbqXIIhvSiBRpTRdiTew4utzzQ
Ee1nt1vd1z0ljbLFzN2ubgnH23RUvUmgVAWsSYqrivMxO4cT/9pIL6ejuoD9dDMk
8uO2B2dD4nR4Z+4s+YSP/PBbeE6r/H6qko9g9IQpUFCvXu1WGdQIpG0IKMYTSBYe
ClchjiHhbNRQaOg2vtvzS+twSdXilmlOA9+pR8iB9+K+XJWw5Ni2AfL2TTHCiAm5
LEFZnczMhkna7DZ6KWymf1A7aWp6EgZIxUnyglXWJK45Ps0ovh2tmBzFl044qD77
FLUnfpNDPi1FEv4xM/hI9cnQH1aYyiVbKFYl3sqsDQ0S6pEjJLVSIuCAOH5xwnYH
vGMGxjSJVB2kTW5FcMPeKy23lBmdQgkFf6Jc6klo5s0f/OLWu5GQluYspKyx6QU1
kpa1EJNFiyo6BES7P9P6RcE2oqmgvSLsRMloAVKV79sGUZAB5a3b2bfSJOWevBKV
NpOeqLi21v47CZNRm9OWXdsasU4wfYFAoIishFUHnmfyTl3J8YjWQUJqi9exxNX4
UIxkCQ3c3X36nf40KyEng30ZPxxJrX4PxpBFgNFIVxQPVa8SmUj6KW6Xog/h5Nf7
fhmgU5Ik8s9abKoqbVQZHI6GbhPA/8iGMmvN5uDxglnWPCD0U6VQ84veLKnxt88O
QvaKCWdN28szuEhfq5INTvzfjjA95r4jVM2ZoXYiSaRyosfPs6/amZ1t+JZbxrUD
PxEtoppJP0XUfTpbmBYLuV9Ufs7m+5ZNfhZBLjsHHB5Ysv7Os3DZar3DOTCbTDuY
uk4xGwchnerAHDjXyMbzo+BCg41dMDXIZxQJhPrROTmqd7wP8kRyJci9O9bL5awA
l/IzQx3czk9yo4VFhXHs//1Ij0x4FQCwIgArPNK2zm622Q31ii9lLq89GWT5DFZi
c47qEZcA4l9G8EWwl08ifV3Eq9xPen9LEXgZ0slqRkE9wcUIOeieydwxsI9+dk/i
nOYJ8DLq1S6OL8Ox/aSl4Hi/eD9ZOi4w2OWTUG5sB6i7G+LidjY03IYDGcnpkHdH
BVupR4SFX1V9gF8fTrkuWbq4BT8YZVK4ZsjAwTtfqw5lGZYWXg9GLPn8Y9CmdmD1
mczgmpHbfndKO54A88lH133XunyBbmB0hgd07cpx/Gal7HKpv6DCSb+1uIe9gXVC
yI4KxllGShSum+VSs82LmH7jQccDfw+KhXhZgouDAW19tUMqH38X1qDObsFmHmaS
19Q/O06A/mKJe+IRpWSjMMyQEcdUaDQCAr6nEYGKmlYBibfvhQDQLb1Fo2oNnw0d
CTva/Gpo6iQRvDCanVXM9gI1hMWGMY0tIwZhp1z/TDyGVEq24bOsomTuY5o2isX4
eGTJs3ytfzBP9gSSkfKeWWkV+20B8MIJBopHH5mW7R9/7pJ/kbjnNX5Z5Mw3+hGJ
bF2iYFUK//3GKjmoEAR/kgc+PyP+C1eJzWKIiYZ74ULAsF3Dw710fz5do4feSkOs
r3s1KzU9UAkfTPTul8ycGS6gMJOSMr/0HokPb4lG50yJBONSLzvKJSjRxwH4dw2Z
pIL+RDJAm1DfgtzTd+uSBU9t3XOt2M5tEDQbj/tKy0v+3ZTE6szsP0jTSGbGlb5B
xgDbcootWqRg8jRdjg3KeEHawbvJam74Jcepun61Q76ZmZNnZwQB4966v4dyIwIm
3dDnrb2QhHoWu+X4mNFF8oiWTi1WruYCOFVHlp4vWiQIXzubnVRcGvr6DylHm/Ji
H3zHCcAyBcfc0pxbtjjdlM0sPwPtQUKzqB17BMHOVWWqNFeqHWt7CSCzn8VvebYI
l192aA5tn6LX6On0wsbL8iyKGCCjEKgo/x4/bNmX6ezTtm/bvN70dByvixF707Za
U+clKucHUsLica6QODLDiPlOs6r0Un6l/LdLPcWQpQ3w/fxvcvVhy7N8PBwFI0fb
Cu625j9BxiVy5Yn8QSJQAOFEY5qYeBhUiT/w8AHHCC3FuIHqtrSqSQ/J43x+17rm
8lA+KoIuUvhyaNdgBfMgjSMbcE5qCJ9sgf7sD0JUgf8qg4oqiEvIfG+Al7ZO1Zdy
2Ddj86SzQn+eCyAnDhYo7TsExMVn4OaMZ2g4fl8Hl2i0JUkXVezcYQht7T68CAwA
cygIc7Qre3yWy3z2lxHIZyiJ6IIS6f5Gleh/nPmRAvkgwUqB8QnjlgW5Yph6c6Xl
FduU369ZELc23tOyF+AzlaJAWMihF8g8I1qm0oGF2ZPv+pnI8Qp4cXZdup7YQRlq
ykVNJf2womOyOg4ZUb5O02TtO9blRhNB6K5awW4EnpZVqmah8KWPF8oQ+kqvdw8m
uHG4B9qb9Cz55RlI2bSHPUeHAmMiN25zqpA08JjBK0GoCwI42DZ+nfLot8FytvLW
KaiFlHU5tqxxRBXpxasIqQGrxn6BaSeTC4gIDHiUdNEcuvqXVEXqnvKNyig/udCF
cA2gUIekpPjAOxm+tPNqZzYsNClvR6vuISx79aYqiJ4/aKZ8+eT3aEg5Zc1ZLo2k
R8NlH6fVJAndY3BpeYIZPdLi18VtBjUHikp1XaeEKRJXBrZI2W5Q3OnH15iWei4U
I0aqPccJjOqkLYXI6ZeBV08p7C9NxK2Ep7GcORddir+ynS1RsACGs2daLCDVSysu
jSJVvYfM/Nn7Qd9CnApOT7JEQBZ1aQB3k5asKsCTt8q0RzRHs8M8xnp0c1zRoSgn
X5kV+WXN/pc8UY3aYMh4EawZYrHwiOuxl9hECQoUdHERTYx9rrK689+MeKMLV0Uc
+RL7dylxYsRbThMFYsTBocSLbr/XgKa56bO/EUwSDaO+A5HmFTRGKs4AhzC3AAwQ
vfoJU6rCsmOSutdZchZV1kqyXNF3mbNFUtW8BN2lYAxk+gZdXPTMeb/FkbjEpi+v
C8jG7W7w6x0O+NZgyqtRv8HrFbUil1n0PmQBEjoFuHBpB8aT5uyndYNEkXnbM9Ve
VQPPVkA9qrPJDHy5X4yj86h+DAOi3tcQyvOpzb28EQIyMssxqEVTRW2kk9hsrwhd
RJmkyu1SUTsXahka67Y1ArE9cT9Lsi9vMH8p9CrSqjBe+QRxhvcsGvV3lbzVNbJK
Idc05Zyq/GTGCs5FjrFqU9YcyY680fdpLTwd2IPxONVYLH/GV6JV2EqoQG83nMu5
YTc8NkH7rwyAaJGoCyZ9Gr5hTMytHZFGPzxLPGdlwQwqei1BwX7dRCbI4Wao6p10
g6PmSTgxl/gfI/SE4HzZVjPKClXzebVBUU6aZqk2K4XKDK+OxV7NE4R+VCkO61hY
Vh7HMjd8DRvbd0X5Z1byrAcxcEs41lc6z1jsvnOGDk2CmZp4UdjmwZUJmbDL+qde
ncY0yZ+NSL/SkFF/OT/5B347NryflWEZBfYszo56wgDaSpCD4tyYK4/1DNmX3O16
Knd9muUKMJFHwfXLsLfeeGPBcQWeA+J2ESEKhw47F/aJk69O7Rip9AmUSyaE24xs
Aq6sJrvfzUoy4NBJgU8YVQcddAwl7Q9LMRwGj5priAe2BfQf//RBXQvVYQkXAKPH
ORXrPbkurYfj9y33f77cGNOV0bvSdxkPQYADZ0p22dStIbkViLbl2S+0b94AYS0j
ORszvEIAjdQPa03aUC4WX+upHiZSAYPPsmuCtLDVJiGmTqRoHOhyievYcvic3Y0j
85GKrwng3wvkU/fDUOVMntFobR1R1hCa+E4y7uw8U+BAMiUw7/nykqirCAGkTZyp
nPxPK+HY/Q5uxIJqRJprkhOQwrIKlX4OyT/lMKtHsrye5gJtGQwe9NpnwRGPN6qA
wOQTvOQwOFMhnJ/FlpnXjZbn8iO03OvYv1MJCeJDsDrYyjdFRnKGfNtIIZc3mNP1
pGV+Zt5tUROnxC1H3FzfgMGFBj+NSn/aCS5li7kldw7bnjK0tyBD6E3IIpoEQjbQ
Z/NTAkTB9YVnbNvsOmXHhuL8ideY+NApKNRnf0AvLBPrJZr3Ic65rpqM96KVLL0G
CpfsVPugm8i2iLZ5ElkL0YxDF27k8VWQuoPq1G2602oGOpLv4gG7Ih3O1gM5lWtx
WK6Wr6U0hjtmU/meETS0/S1jT0MAieV8iew5AI42zr12mdlpZJKH7JS44HEhGnoT
tdh7CJZcP6lh1+4M8WDzysUdRzyA0Kdrh7RI/IMb5ZaXn0vQU3qR0O2TAmcOwMNB
Fk6jV9biWzDFh8qtponFLo/LQProlF81GTFqMTz80vXG2iD6gE3i4ewJ2VPuZmbM
lvDkcmoW3vuHuUAIpVQrWwLYYxh13HRUS1SirijgleEXWuQC3TDi+L1wkkxkeBHO
TpuMAjuUAA85mXmt4eaH/2vVwpCsW4HMnmHJ6FHHUHFKVdSzkPrKqbUqjcwhfTc7
7mPR8CaApc7UBxeTriJEFyVjVQJ/G/DjtYyNA707fy2VhhYdVV/Wi+cni1oKWZ/1
MKc7tpdrALJw8ou+C/PtUmUberHEucDs+73h482hYhHOJ+yZ3WSRsAt3qPC0MZ6c
edmwIZ9CMhGrQh0d+sBCqAHqJweIGpyXnYIRZpFYdBmHsqdoDPSQnjPeIjLe0Fsk
UO1D4zmn7P2LRzUVj+OVZ2l3AIHzONpVCLbL6m1uOxBU7qCV4ENflgInsuHQHzwr
u+ijJSy9tjGV6o847N/ZGAWtgP98FrXxsEG5Hx+ZmIQwsJtdK79dIrY847OyuKLg
HsxnQzqH5VIvfLr+tir426odG7mFcIVeuMgYAWwcyohSyHfWu6TE1UOxlVZSiR+X
Oj9XRoYU98VRMEk8oYFH6jPlEAqVsX0yROVUPPvgbek+TDLxDYawo2636Tpjuqyr
pFf7D2WG8sZzVQzJH+pd8VRvyMuuC3+dbEPKxF380ABytVJax5Ro/OtJzg3cbZfL
/ZgRRyzYLqAlfqqrrPXeKmSGDV83zQ579lV7qDfauZUbjPKvjot4nwFdj9i3ycWo
oOQ/nJCsiSkLY3HnV4PhCrGRUdiCxR6d6IZ5qDz/Kh0mdfrMA0tKZVvSscsbCXAA
KyDOP85WB3kA5cFgjEF7yn5EPlLp1IREcWRV3iGlYfDlP4Lc7NyUifdrJKsLazIW
Epe+as1343zZMlcNSimF8Yky6fYOSUdkeIFtO8f02yLGCcB/phvNkIeDEfOJ30Rg
IZI/qt+cO5NxOwl/Xd9WTk+B9uUHtA4T/f8tYiHQDapjy5SPYG3q0NbghMwNq4Ou
KFnhJclTopA1gGeeCHjv5PLw5OC35YINBaD1NfqtWY9p4X/gUCkcukVxjSpptmXT
ARFtLMzCPGu5psM6+WYPX5GmF/6XAX8+ONQJjUvrPoY3le1Oiij8uRFkIsyHzWak
l0xuArpLOS2GGvXd+o9Loef1KjPEmAwCgXZR93J8pKtX2MFxDT4EOjGxX9lefPLs
qkVp+8ejpb/GJvrjqFFS3j9wHhjJgiIiievAnlbPVidiDnyPoxip0sCFZ3NGYqCq
Oe/ov62jUgMcYBEDoCHLUGT1qpbrWJ1ZpFDMfxgWg2zEljNyIjmdc6eqoDCTU9Pl
UYSrDRv/HQzqnkz3tAsXP2g1PEGMdWirf4AqdtOhvHFuPy7bBJs24TrIjoNEqQuf
af3vOOgD/9Ueg49mxWrhwfP91Wkrrn2+AZes35IoXH4MPU2DrVCUoJyxqA6EoZzz
VyCxmu6uMmNmLX1Gyamg9zax031YBu/monG89ggwzglcUxGvBhm8MqHECnLWKcIE
rfwOGPS9Rh4YrCjzKLnxjyXNFOh+P3/83ttQikoOLs3/XUZbO+YJzXz0vwQuL87h
vZyWdKYKN+0FJvTRo/+iWr3N/oFy480Hx+RDWnHOAt6OOOCDTeOVV++rhhgynvne
ZGvgEJOkJ84kzhbAsbOvzZsupG44+DBEuEn0ZXO9JqG0L+GZ+LOuDFjl0iM2Af+D
4r+IY9zyl9T4ixF64EPsTZ9iqR23a4veK7hy0sFdCjYF75OWDbafMRNaeTTq7NJQ
bS/VD+qpveR68j4fwxCmLaKmZpJndxYMI2u/P2sWqu/uOW1e9V/iPCJRW/1y3DjX
jcS2KRRh8XHrRunVIqHIJPEijxbyfSstq3+SakZZ8+ilJ2AJAAR979Q2NRwM9lNv
9Gd9qXBGZPBvS19cfouUJyKPygwMrgD1yTlqcGDRfH/uSQVcjRXrTjpqZlqtBFdJ
+7DOfbpBjhiawfwAG2PUE5IZOHi/5lSvEcKYNa16AojGuVZu0EMKcD92+reC8DgD
e7r0kUfylfgGq6l2B8sCTcX8zRgZYhg0ZKfcSop1zfzaog6gkkmh5atLMtle/HMf
Vc6WSypcul5VsMCzFOdSX+emFm9MI5IKZm1Bz9pKHogCrz0CMd90zrqnvo9vwa9j
lafjogzfoEElltLxoyjw1WFgYkTdnxha61R3+88dy8M9Z2vt1mga7NsAMm6RU0VS
ZeDI1/5W4uEngbUI1zBnijCpXVuhSw8isXdBYL+vqI9/Q6NF8ZMZUrShvxP9Cmql
KKfKbojfei8M5jYDJhybbgVAb8W/x1zhvGWCPE8HvPDKtqFcfkmhcKmvr5oz7Kdm
HDWXjmTqTRo5w6oMT6yaP8T/8b9yBXNopnE6IQSCakcsM47+wTBgwt3IxSFEucH5
pmwPNbtIcJz1kluYCbs3Vhk9lzwguuZk4pTYxiWJaqswly/246uYRcsyVWp7YbON
syVz9ToHI/+kPv6/k2hrv297Lz59R8m9Q8TLL1XtWi+GoP3Vni8yicjzo8I7L/bG
KUnO7wU7SnYEc81/9lnd1dO51OTyRmFGiZvYesEhakRJPialFs8Idn5YDPWkTDsk
y4NV47pl/ryMXLL8J+wm+VXonlrTvOXiCguNED3+Ra3vLoxU5x7jlgeQqc4+umsf
M7u6Msfg8DPxeIWBsGGF3jw13Vt5R9CWaEDz6/jTtp6iUG0YS5dHWXR1+PXFuFcJ
KH9/G00axpu7evxGWD4fQm1QMF6V4Nyw/lBLbY0scVbq0ZqFrJOyit8OuSet9EKx
hg9XQf5ZPb5fyU8x35KIE4rOWWERLuU+TX/px2usLhVsR6IaS7PuXt3YF9fM01bg
tihkoViZCsH05TN/SCoMSXSOXEQEfD6QKowzYcuFh7g2WMA0LBpkg0/xClpTI8bq
HDqRixS0+CAPtiFNL95mPLEXGs/1hUiEO73if1lFJeCj5zz80aLHP+v+nFUr4hI7
jKklrQ/+qLnj6ZM7HNqRCp44xwH1ZNAXIu4ux7mOxn0SsFfuOjWHf88MWfGOhUmk
dxiahWxD4yKs6PbkicdgFGJRykzaNdpmPN5t0tOyroghDOOCOoiqE+bNZcpLpnBr
7MlbBECZswL5yNViFf9juZ7lJAgd2PnQFw6Tf4et4ud7UCqOBB9wIboecq2egRqy
R2RLT2k7KHItk3332XjqW06nxhVQdjePNJjc3lZ/hSeCOQwEZFf/L91mpxdC82BN
CeIU2t9i6LKiN79j6CAT+m83QYaDtahaZrjYmTW7VZfXSMDFsXoYvpkKYcDmdsxt
1biD76MFxh6c+yVYqSVP11dSEaiiyuKROrPAeAjB2YGDvQAYv4ZKxrLPBPM4AQH9
dw/Wk/94Y9YnasyV5UBrfHY+0eOdYGaxrmBBX4LVKutG+76E8v6sE/P/sIcr2WQn
3ns3w6HkyUC9uJtleSkBkvBzOHEtf0/qBcithg7tKBhW1FJKUKaUOKVWCqtJQ9Qb
d6kEGRn9TaQQQmqVhTSt1ULxHdtm8orglTAjqBZy+ll/aJvZZuLdje8jGhHlXvB/
98obl46SfZ2QOFbLyULQTwkBqkRL4nIzcBE8Xli30jgutWgKgTcDe7iPejP9G4GZ
ZuTHmdVLxoQzrBLMTlSvORAi4KfOUABUIc62ISjlT0lFjcTc+1G08GAriLrt+yai
MJHyfDR43EhX5G59jHCDqYJHImZILJAhKE4mv26rRXiiCScoZSH2OTkqKamjNVdj
NNU17Zq/K7IA+4znAe2FRkCbDx1P5y7oe4UHlIFvZ6mMVm87VyJFoXqFMXQxA2Gc
hvqZ+h1ekzFJAStTNYzsSLffKj0r2deKf69uBNF0a/uzgq2pdkE3jjzhWfru39NV
xbig8irgzAWyNQnB44S9aOWmkPqfQ9jA9I2Lv6VLraK5eSfPYFQ1JZA6/KKyJVN5
VW0sCDdR3CLZHn3LHIc/VlXXScjMVgjriABnLyB6yYfZFReCF0xM235kN46m3mBM
bMy5NJZ/iZTTTny1qn7MmpVJMYVnRig08xslaaDAypIFJYz18rErjPJDXtiOBgzs
rz/jVfSSQ5AcmBAFk0X9QkYftwemyQ2diVC155IZkzEhxwaUsK3Qr9lE1H1DuT+N
35pl3epHAevXABz/xAGuu70526MSgWLjjbXPY3rKPh0IzharLdalQjefT9bfz9OP
K0mx+Xkmycw2wodtHZ5ohzYQOofwy7uj6zlh6cjF2UzwNqtA/406QB8t/ZLWWsOh
+0X45bCOplkGI15ngoo9FBrmvolra+GfWoTKdV+z8Ji1lXKJatMOhzmGIE0RRCrL
bOw419RWPrP6PyzjTDNUJUr5XviGMzUTh7ZZM/SNiylTLt4oHI1BKq40Pkdr4WT+
owY7BqVRdocx3iMtqdUfd636NH3QSwe5+k2yuuKDNDmbxAosQt3X5WWGWllgRvbk
iNcRcMDbkhZI5520v0erYaDmLIAHoipok3GP7gxa2YAPN97yFhvhbBgLmRFKtV0o
OUtvWUKFo9ec6MhgQjCQtXPENsd/I+ZeHSgpKFfRvGoLnkwfJs3ACmvywOvhCOCg
0RFDKCOGujPUb82Mm0GNBawZNMX9Z0lmTB6wfndD2/FgKaPLFCszMTUl+yduHafm
QO61gqzXUPl8c17WiWSHJxVSuwhG9Ebdk68wM3JHoz8Uhd7PkOA8Rr28WSAmTwFH
mFLOVf9AeXsQ3Xfs9rSbxs4xFAdQUNZqmmnmSWljk+NnA1BHyZVFscw1b/hl5opJ
DhxFAsldzi1BlV6Wa8KDrp9QYBiXXFAbbo5WTAGEEoIJCvPh/GnZSbkNSzV/aGzk
3N0LSRoBxa50o1j+pFX4jybotK4zVGSvns6dLDyFRYhnkgQhzt1t9SvtULwcJKsv
eWR/tImglRLeK6ND0L6myyYKK4WKpEWM3cmAgCIz0AxwUcGhX12krLxbpU1e3UiM
75Jml2A1n21cKW5b4i1m0BlV/WjOASt/6L3NKhpevJoOTog9BnaW4wqr8rSSL8uK
HkI9HsPWcy1cvRmPtxc+vUAlL2ylvzQYWhKm9KnAiKcxgA4yHRLmM0l9K8cFBCtl
r6ezcyC2HNi6FQuX4T4zA8UkQMODoN2s7mABLNfMTYRIFBNDNrfYrH0OlN6tfMfG
Wij7kjqABUlz8ssPeBuxLEDJ4TPBQZQJaUzFTzc7YupLr/6VhqZHoiGQ8Bh8yhIo
wN3Rk2OZG+LU24eWAA0BUbHEc3IIxqudHgUaL2S2yeCbWjGr0cQHajfayek9nw6B
8iAmwhzzeKtdkQPeupr470r7yg3EJDlyRwTf90WjrI/8sijkqd99+VUjTMkL2Fsl
3z5++6biwSOmyaSimvNgUp4yQM8Vj2bE+p6lvVK1zOq0FqC+MXN2ltB5+xISgK4T
8Il9XkjU2h8kogbxv+MPR0nFyG2qoajPHzwIixeVXsHXIUq74y80wSiLwA3e0yo1
+ji/xuvjKXdFWGevhA5gyXKwPhxTbbIohjdqD4FG9Pxcr1AHf8fbVRFaIF4pmq4b
Lf218PuJxuxuP7D+lKbt2amLqXe2mDPan6vYxXJJp3gXeen1SF/N/RQlh7c/V/8g
loTKqDaeIxFQzP2ab3xPobT9w9w/zyyL7f+QuWRnambnejBb700yWD8vciUQJ457
2RGlozK3q9eYqHzgIFInq8iA0ifdxDT2+rQ8c5gXJcEj3CLsWj2TVw25m2Q0OvBo
d5NO3VOD8i253lIVMVIrpWhCGtHraut6wbQ7dk/m/xe5cRlNkNpwEccOJm2WijWk
opnOmW2ovOpVnJuRu7TxTQWmJe2K3qRAShmNjPXGZ3Hs04Mw5cuHScpEna0cIthU
GN99Qgmtog2U4+DfiqR1t08vwQ7fBQhynOqIOGIlvR/rq+gDcAzZOKU0qM30hOJ/
qWnCFMQJ3HgyCxpR5LRLcwQA81cY/ZLHM39FiSQ/estavmBuc5wfQXbjsA3hg6sX
VABjJjEROvBSf9ApH6AobULCrj9eON6oG2/LPwpDxqLfqzDVfPlNmsJo741N7LZw
u8wPpPh4WSJ0JHV3tjyoPOiAIEFLglIg7ImLe0s+ExIZDwv8fAS1CbQAX8AZWy7Z
kwd2jQ1zH0q+/L+Pd1rM5VE+0Rh7bCMALMF9eGpo3TNLy7dBBXKcU4bNEKGehNAR
6r+dfgKTmKki6CJemqnk5KjEnuiYpVuMOsPc8fTsnuhY2FrH6VDew39IdZKJ4SW9
sIjTX4/Ej+52ks/hR2vjOKTzfwj9fnxg7UMmdTJ2V6XNjXK5ly1iKM2Ho8PE2748
Z32H2m/XZOxtTBrvjEgxYzmAcEjmtt33pp7nzw2lzPFPQKaq79BIRvhdFRbRo6oZ
q6gtTr46Dm5sl7oaDv9z6cQe6TC+pvoBeGuqMIYIc1ZkmOaptCLTD4JN3WJWkFqZ
Vubv1BqCzAg4aLenpWGNCT0HDcZ9PDFgUgkRvwsPT+KX2Kc/ND3haiLCMtnEQ/GK
GPleIc59aApfzK19JpHfz4KWpVi1dykVbNJ+LL7wQhkjlfKYuYAnCd0gbVb3uq49
3fzYEdOBrgZlQTYeDMqoXkuD8T8t7pDX/waM3WtGDqiDWY0nSeBRGBebctTkPZm6
VHoJVecGbjpoNW5kjl6rI5jHOcKP6Ue+gl2gm89KIpQKuXek+/7XivsolRYZ51zL
RuqnvGE58N0z2Ngga/k4+9UH0N3hN6PUQBJ9/jWVpZjdCctFch187hh9GDFbJapv
B0QI2F8BLVT5kY8CTOvtkLtZN66Dp99XXVqZqOty2YpDbwiyPXfmKBEOfbpm9oIS
XSs/S6SilE1YCUaRz86aTJ73DyPSTjWTU5GY77NAqKaTItULMC82RzcEL4Tz3yBs
IVcA8OJ20xNWGxU5TJDGRlPqJXDwlDx5hJTNzVggGFEZYBJeLx/l6882U1TjEjdS
BZxC71rp/a/JtDsOH4Egb+7gBvLRl3OOSMc1pwnQ9S2hkyuYtBSzNgRdR6cLidcb
8BoJArlnjyDvJ2z789nivTqbv6Ough/qpLDjfrD0EaNAXcu0h+BhYm6BqymFia+M
/1SyIt914KOjP6rPHZwRNwVVnmMHknVroO5GROtH7X3L8ul4f6pqWAxT4c1YFg61
lG/zYOyasMbw+lXk3dnH+wk0vbrP3rJH2fQXPhdzt4+ysL24i3CtNdoqM4p60Ah8
mkAYMZOvPHnZD1sr0CdYF9chHfePG4UemYQ2UUjxRGIi/puG1u+R8zPEU0rm+s2z
S4E/NXVZNhHmmSPgoj5MCtH3ZxDbyAAVViWmb8BjsBnTtFBNDbmEdsFEB7oLclvP
ljZtbxCyUNKItsvjdE/phNoa8J3lm+x7Byuj8BQMy1b4Z/WS9eAlmoa2rZDUWaYX
dx4Tcy6hfoKZYqVmEvlAo0fkOpW22KEHtScYNh76WnELh37GmCnN/f3Jlomhz+uN
LmvWUB7ytbSLH/cLNcNe44ml+7lfWJGatyfuGdgdhzLEq+8tIgKKRup5HFS26Xkz
g1OL7h+rbuX6HkItWS8e8/QwHKkeDuPNdMiDjxlCc1MHMbfE9AQcUQUYYoPOAvsM
NbfYSUm3xq2H0jg7nuPqAoQYGAUJxIIDoL4bG9IxqJ5/loyBtbOcIZdmJ19rKVIH
IZ53Wz2umMH/3iIHTiG8oa/oxNyvQNw+SrqnB/t9FS+qUyjqP6UwdDdjgHWyejql
CxPX0B//m9R3Cw2Nt1tKdwZYsM2CZoO2H/EMmVEn0yj9ZcKeN4X81quzAksMZyo/
DtCZyksIy1roJKuCuZM6Sv69mVRTXzZ6E/Gxn+fJRbZqqHkDOfApKtfKzT0e+HUT
JoYdipIyFLJBMQmihowoMUwNdPvsNKe2KZ89VvIdWpU3+Lrw0JZCWX7KDf1Mf9zU
2guLQffTXqigOOPU5t1L2MaheDEAKc3OHOSzM0Oxi21L/uRx09FQlVBV4MqzU3yW
fcLkKEfEXBvV8k6jNUt4P1hMesV2bexkG+0utYaSds35bwnBg/4Oxi4vjQv7S2qe
lVerecx+ezxACWZ1Xa0mu+Jbx/CDwPfIqbYeAHqnYtuwQXcC0iVOxBZfPZGT089x
5avR8YdC41+Ul1+fGquX10rz8EEj+JUn/I88QouaTbeNK6KjaAg4k8swhcxwkax/
4iZjKb3X4ChMZCE0/MUq5zF/HDYweePM63QBS4Q+MR4hKXBxlNurcDpPeJ7gugQP
/bfNCzOAjTB+TBVSvqvzEb9iJIvRBtAMfTbruP/XWXkmzHpke3EGl++dAJpDmnHd
3t4SbGhyaCkzaLRW8vdv+ipfqgMIt0a+wfK9/doKouwjRoT7yYISPxxPSSEMm+ts
7NqHyNAbHFv2nh2ueF9w3U9sR+P/IxA0ZEFBpVB0qOzBvAEGi8QbzswjFDffAIZs
GEG9f3Ut3XEAQFPAFMs6lttiKW8f5p0m/Ae8fzcmCH/21XTCJ9Kl5x5DXtkMNqWq
VlDYTgnUyxhhfGWrUJaybLfn4Jv6QntWJELuvdpN8w7UbmC3UYVcDNdSoLgqeXTz
hwtcRzNO9nifLKIkvpdB9qBRjUcpQJbrtlXQ4XfEcRVh4rl8QRVy+KX0J4nD8Z3d
te/U854qa70sgWTw5JMM6Rz4SGvmcrarJrlTBIxvFfLxkzCrO3TGkEmFTlHFxFtF
y29hJ+kOuq8NAIfLG6OmYHwRi6ooX5HZQBaYmBinvpL1Hm7SbuJLb+L/IQ32bH/D
NkrMqCpr9p9mC85bllkS1z9FFCsUCbzt0emIZfh6daU+cvX4CR2wD4704YACtUh9
G4Nds/lghBnlbgsIrZNCWIPbS24Py2MLrmHLdPbcphs7Cpx1wRUbZp1K/kf0n82d
w36vXzrW4HgF+Q+Z/tqVUQP+Zxx2liqEf8YMiTA5kbJYXAGmJfJJXjdCEcgvi2Ct
gsRNXmq0esYyDgxIlSeewWq0GV9i+IehHhm92vkPWCaHMrYiNyLa+67qGMYenuL1
ThaLUP1o1gZdF2AeHHdgKNG+PblBCPcphcFr9tndDw5zqjTZS+T3FIO3a/kOrhKN
GLQ041sQUu3Dkf968gA8HXL1dqObDMIfc2/xhFaUD9W577FtqBCnPEVsJn8Fx70Q
aO9TrlVAYbhHxAJFwZG7mY9PafcEhLXbPNZ2zqurK2bhMzIt1tEBtHD7m0cyQgdl
R8vVjAkVPqnVdPLvS/DZolG6HOBaYrZWnoJ8y/RT7lS52ooWa57gbYIFE7ualvHq
+JoW5GTxO5meF31l6oSLERsIywpeOGxaUW0r4hgxaqfqUbRps2XfV29DRweCS8yH
TtcDLNsM5o5bdcn81Zb9YrpCo9IP/+LGc2UDtFoebRbtQ+wSWIGNzfGitbfxwuW7
mUp/w9XY5mzJvwIhLbz2dXKXs4ze3sV3XtcZVUari0ouLTa4U2qwpltzacked6st
Rv+3w0lX78Yrt6GmZikh4Ix2vlgj3qDUHCT1soskuAeYCaADJFSgP7DpaFaWnkmB
kefbemvqgGl/wuLSH9H6g9ucUtm+9wH+Q8W7OD0xK/ekgvw7niLvjvKiumXkiWST
+p/Y5pPkqiAVQz/WWbJr2XXbnuu615LeAwxpaC1OfrcdexDdhHqBTkpR32tF0ops
p+f52cM04SbVmN2raZXUp7T2iSQeMEsP/N1ZYcTpv58PL2VC0sfWISw+7Rn+7faU
nCN2FMFUW8uLr7+y0UP0riM+wRunN7U6J3Ds3TXVSXDP2lQYl4dw1rxCS2F884mw
/FXtrWbyGlC6fY+vb3uIbV7GqNg8VLwOTgttigpX384Bqs2f5rr0ib+WAfakC72V
dm4y9+tUdHmIwHlHAH6BC7q8LglFcOC+vyVUbGZrj+lETK1ccB5DrtMp9FMx/pO6
t4wjWMTUmlNIvd/tu4vATPjLY/7tAcuXpFPDYpBYmYKa4/FcTK5Dv+PLDIQ8XEW0
68mphg7GqLVhy7LalHEzexSDSB2vSZRK0A8psXas6S2xtSnLvONTkfe+kfj2cBq7
iJXhxjfOiDKiD29G/Xncb9DeGUg+1itPdxBiYtUp4UOQ5kdAUMQp9OM9ODrmBZW5
TM/3dUZoCjYPLVPUnNPFZ+PxFW20aqGyIKtL8l++i9BQq0cIbhupEk55p/HyBUa3
zvwlr/LS+KomqN/15MyuGvBAfB3GfomVjLREQrgPCvprc/xpH+dvuVcE40tmsTIk
67lVyyjirengOlCeTtf3OcKYwZr1ps9MF/WeE6OZ3jyNUW/z+iZNBOKRrrzzWoHk
z32UguXxiEjyfX+LASqiwsCYwJIhdFdZNDYqoSzFeaHmX65waYfVAmLXP0aYThmP
JvrOCnfKl3Qg/Ji/hgiiWxasOfpD7zBhpi7gdVIH+8QbWlCBnd5rEpyHTxY/Kevz
Sa1AuTb3vjj1CxO20qkkpaO2kYpVIl8aoNfBe26oiCxRZsyGiP8PK9vFMp6MEysd
boE4m6ul+tIew56JzFSG5NPyeZygUYcrPop1rSyC9IWZ78v/7GqZVk3zsPzS1mI6
kZKkQdhib5YRA3BZjTKLJo1edx1QTatjmKO9QZvVn7uYn4QhSYaSf2xPD2T+8d7N
MFVCfcaTMVuXXB/n4rVVAbmR1n9JLxkqxj9lKQTMq1yrvm+mgFUrWYcYfE4lsjql
LxXarTWxgDmrumC20t9n78q9YB/N7Vl4XpUQNvTIe3FD5l1rZ07OapD/v4rqFIJV
nH480T/houLmtzCzbaEF/2xwvKR7AUYggz6+enNVzj1e/9gDMHD2wyaE0jZS0Zma
yxaUXM0qgoZpKp+21mZSjv9/R/tWX9X2kdXgYNoKkaiWjAacuhFd3LaVUCu+7t/w
W7ZkYMF74ySb966jhP6K8EifkOsaO787jtdFlr+Q5RbQOLWx1FhzcqK5hPZTJJpT
y6R1pnt+PUnJxJy11M8WesDshqab9s7GAy4+BHXl2TXbTglom6DiSnU3eUm4Ybe/
apMTSmpbxnJzhSai1MSj++eNU1k0h477JKx+Y9McQkhCW8yXY5AS+SP4zQaOXR+R
dBst1m0LOOwriDPtb7UuITDb0H771X8MLAoiqBH2V2+cyxpeF8gKJSDJ4YKEH5WW
Wbrj82bW4wAjY4VSl4HrEhQdRLhgE5W+UyCgtjsh5ohcwsaabsKorsCt0iLlsHwz
4Yk3C5MV3gaz6B0spSOPp+Rcic5vFgoVFPFsL1IKo6XCj9+PHDYBeybTpOX0ElsG
CW5TM+RnDot3RHzWibA4g2Yb/d02FzH9JLaU4SD0eDzLOG2QTy6f6b1aYh3UC9GF
/ilY8iM1Q1gjyskApaijAdX7KMJ7eK1f0ICWMHXNd9zjSjOXC4AxDuGjPlzZyvYJ
EZLSIDnBTZK5AMKNiBSr1Wk9KSTyOg8zDHRG9E4jyIaxvL9S7iJ4lXuVv4DvdttJ
RTzqbsn+dYXyFp7zI/ScZZgoTL4HXhYHXy1/A0cAHQiUMuF5Tx9OVVaKgz5tvage
HJ3aPTkNmxAOFyxFZvDQShDcV/Aq9FH2BhgsAwUC5bFFiwv81yriNNVcCdZnB97z
qMFHTFkd8HWQBCYmkNS0P2GioCYpWo/abIPzoLp2R7KIC/KAfLI3yz/j2CsG0dIk
NATqebCuGP75MGngRd4Il9W+zAFBzQa5wT4QAB+YyFsO18FzybK2wtu+FVSOf5Jz
CLiyRsaWN2AXZwkuu0FT/eWs5z3QVRqLKKyzT1yg4ef8tBnmH03R5cvqBCFcDf5h
Ogc1pu9PIaTG8EecbO9L8pqZS5i5G9uI81dfFoYhtMMPteUkyf1ttG1RVNPcPrlC
JAbrgfiJA7WIzt7rKp/buZN/JccyVFjLCuRbskg5VQaPSP5qiGkx7ZCkxtBSg9IB
6KHXZSutrvaxReqhsR57CmkVxuUC2ochIeDeu0Wo7MdEYeP8f/suBZLCQzwStffY
fLY4Pb10M1zzhyf7zSq4DONpN8rn6cRVh6UBLABukVVFbxXG+zT9HASqJLqtmwWh
dKr9U1lVcIVZucKox4MoV/sKpaYHziOdi1bQlFDKPVSadVQlwkiHF5W8xIVOJNlH
P1F62T954nAjbPOdqg5x5oH+wwMGv4iT2ycM8FgvPENivTjKU5bnajC2sOvIX3Zb
qISCLx5gQnO15mkW5wPbunvweRAvLLhq3YXQhKn4IrbUqX/bIJXa15tMzOv6JHjL
1CHkaJ4ElIu7WlqMQRvpkfS1UFBgHewoLWzhXXJtS6d+vsO7TtbncWZrH8RV+VfD
yH88VLeKwIexqBdNZAjFOZHVEpEp4/x7NvfoLKvaVt7ufJo18jvl4D6ibR7Zi29A
L+5ZBMv7MUBTh5+1OPQVwGLJFs5z73S4SpzWrqqmo6ntgkwOVx8QhBanhxAyfYbd
AMpg3pn5JpHj/ID9cytRuz1C3ZuNu5XyPFhReh4XKikVNB5P9lDLNTwkLuBq3fIW
tN5EsLnl6up86TU6QZYnRVl089OLFSdfXfJfcJ7PnUJMLQ4HEyLupzssaGbZdBqW
yrX5dmAQImgkCJlG7nPEC2+Tj2utN/BTo2zBGzR3OzRt/Hr2hnWK5YVXddqfZ4M9
CdilvXXJ5JllbedxWlwL9fXiGXkYWA+acABdevVWCRd+NIEnC2o2xE+TU3jsXSgq
I7bb878/pIyMOmLZ18+EQwvmPPGZBRVw64hU0NPQPVuodFzoaBohvEGODvOlUBzu
SH5zlbo8YVhZErodzCmYpVZ4mbJEqrKFXgpNyiHhTxrzUuSQ0W0oCOurrOcwWLxk
WVuYrnYwtEErfsV1JToW6kKYDj9dSFu1HWJ6lLEBzC1aHe52ceilq/SuXR67lGGW
Gqar/ARKdo0MQ0rhFQbVN223LxWOkX/O6rZro8rYcn38sgW/HxfrJLZT8atPHu5F
9+mdBzhpcuND8hj5jvEnBFCn0N0GplJUs6oRn6zWR1I9ofiPGbQ1M1Jkup+jVhvf
xevos8N/cxSXJFxB3McY9Q5e5SpTDAUcxC7SJiJTSRWQs6UECelK+1CpJtKxni8v
aLS4kcq39oOqyvYuim9gmyrGwwSKjmFRBkuV4yOgGY5h8U3q3YHDmqUKy4ugz4zo
p8n2N0hfPcnbtLh8aOg6q5uQGVL5Xe8k0aGID+rtFdrdDYy7hF0XYs29dkZKR0b0
CHoNbcHmHsXbMww4A/R4VzXla3JkQYj/Ddzj91cOFQhzeCZ2v9LbI1aqiqE5M6kc
4R3lGl9sCv+FUSazjHS/LDyeMnta5zlqVpseR9KsBRIp+S6i1F9+UihkGRjdcUWu
06r74doof0UROot2MjUKqqmX39WjiW2hA4+jEjj9JtOnX4mIoR0KsxsIX0zcJs2e
l3HC+oawFc3DOQowSwKSKf4+QYgAiypVQzHEigmC33F8LlXGP/aS710kqM3UMR5/
AboVAPnxXpwLz8ArDt+/3rAltbqmihZyCp4ySlE81sQZTxn+vuQuVsTloGHdnvpE
EOntIGJEJGAH+jNN6HqwXLpI0iNcaaWwdhN6s/rmFvRIRCnwFCus/+xr0CaQ70T1
sagr8C+/WNB0h2FndUev+EBSfI4+EzJhkRS7VKoBPQmBe1cHbPxMGwreG141nbaK
3mpaf9Uiarr+GGKSd+JvT5b6iXBYkpemH2dUf1p38D2KE5tmE1Y6d4mxkPavaYxO
9wMnJKdR1xhnERRCFGl9/AYeOnEu4tamXsVcmr2WKYSKveemBE9+cFPhNuJ5OAIA
WbDf2LUR/9Xzk8+eCt0qSBFMX2qymir9SByDKwerqnES/6OpFpcEpzfms4KxVpFZ
JfwoLglWrJCteapsfk3yUyCYcZ9quNKR6C4EB1xMP7B9izuaGwG3FRCVSa69zKbI
W46QgkajPQ8S/vnTNIIkvi22j/IrP/fEyRkl/CXsFtYn94Upb0inR04IRLMmWRTg
vyUzjQtMY9M205JrjNOA8cWDaTfRnW38cBeBwIbl8ecJzaV+NwPTxJjVn2iEolnI
XhCkbZZJP6VxM7L5JBlxcud0d21PLb1h0Cul7Vnamc+V56FHviYzg94qf1N3KxCr
JlEaoPLUOL81fJmU3iIqGu6zZsBkJd8LPthaSD6D5C2hFRP1QZ2mU0RN3XWDjhJA
ZHGnT0KQQ67jIEqqw+bcEuzh2ATbmD6qY7/I00jDfq+OHBwQpfmjeTv5hA4yFVf3
6cu6j6YpsRMssO+dDqgbEOzOW4EXyCEHd7px18v3rhsEZBbFLrKDk37Yp6jcavq7
nkk6AFhJnzzNV57oXPrBdIqtme2+E6dABO2FmV6yYEFUOrWWWfcgUMD8dHMNXAIq
BFArd9/V3l7p2/1nOsV/S5+nmdNqUmW3ZcOL8tgTeR/4vyU4tmxfTXRSYO4+Og/D
Q/v+4MIwgwOVAEkE5C+YdiGKT+EdtzbQ/CxZOLZSwb2otOL1WwVTilEyEvnYWCS5
1pGFyuiXRGQe57xPGQSMPws2srmOCPVKGJSMvmDVdja+11CpYn2lAFQgs0ANrzIS
6O+HDUrq0r84IL0ODcTiGIT0/9wMeprKuz6ZU1tWKglCjbAct/uWFpALRAfmnRCH
5sQaSOMQAMw2w349b4rlBkpkHHp1mjfchltRftHvTVaftPXfaG4mRkiC60xO0WAR
hbK88Lq5njF1LhMs6Nz2KASkuUwnt24BFK6mS4KKRU+FsLau/dyxlmJ1917Qtsgw
EM/vVsizKiZRIA0H4LDJRuTrAfzYMzsKTr22oUhpfYHyG0M8frAf0ik2XGNVq4Qj
4A4GlSa0vsdF3xhAVEipCbyT5cw7RC1iigMDnTAQNntLZTsXy6Woxr/1o+hrn1XD
ZyJZ/fMtKjVltwnc0ZwPaVyyGXfqnrtMhrZO2OH5e3hEAZLTJNqoCqTtypdTmN5p
g5OLVlKMIrQJba6dI/6a0NtQr3oiS1/biI2kaH+UmPlyyk8v2nsXPi71OLVU6lwV
y2c+5f7u3qP7f+/j/bZ3KTy18L9ykxD3ubCh7DgeOdhTG7lkEPmpAqfuSUDveSwf
nZHetHnWKYNrDDrspf3xGvvazpHbcVaZTFAWmoc0Qun9LX5s4DRBn+Pw086nicnB
voJdLNfgFf4kzoeNIxynoQNATlZjM5GZczrdbC2FIZIcl4dyVym+LyqL2AFQnrLr
UojofnPo/y1JwaOtSCPTtsUgWWQgEBeVtn1A1p/4DRo3eQW+oDiz1BAwwNYGj7lL
R0O5JOrQ9aSdQHdG3ACUxbTUoII27VJlzoO0sQO4b+8DgmL/kYDHM/0LVnS7/8tR
wkInYgnXLgdsPj4++OcfJPToXiCv5t5lkIbx+zAECePXEacWSDZdYP+5MpRK1Dw5
cY/zfnoCc8RDa7lf08AARNV+KBlhr7tY4+yzYaopFrZq3RtePl3vIBCyzk88jNUp
wHq43GrFMOgHgW0IKJx8e8FubizbvVYcUlEaZ0TjmDrWs2kmcPC8PUtaDLuR/2cA
+8Asd7myGWDXIw+42Zub2YUSX5eytMPhkggmM10vYTR+HnYtSN2+YHGQs7qjHSLE
jjc1yQV5Dqf52MybRnENhCwITX+CT0xCEHpUM2DsHH8Lo0+mHAWynOON78IfxxzY
rldMZK9AcJenXAOBHTe9LmcMAEBa8eM6jmEAvbYqgkey2kzQdC8eHDz/UsHaZrHd
WHjv1XxIJ5zqdgBq93W3RE7y9819ig/yk5E+H+Kysh7PNpBUn7E2JbJeCxR32EUB
9bTjjgMmilFcdQPBpBKZ9slesMcdWjcdvCO8sI8bMs7qbvm5/403E9zfcQiT64Bb
J8JweEprpqeZuRMHokERN/SPYmpMMzIUlbc/GZz7AEtxyUBgBib8CyNitv8JnR2E
Zw7pkoR8ouJaw1JS+a3YyYpe8wSSDxU0CQ4PoLbrLiP6OVTD3EgFGxGJ4L3HETdZ
VQEaKz3wIhMd/IoGmGLKs8yw3PInqv27Qs0dc5b11T//GhBQySLqmT78bR0vGpvb
FKNaNAPQjxbZLWjQueHQfTnFN7ip2uWBJAQCW+gAqF8lYY09779PUxxrA9L75lpa
/XdGnz3V3T2+l+kRlvp60nn2PB0EAk+6jwWKO0rWBxf04UhTtLbP33i7UUXcnw1/
FvXCRNPpo0agX1vb7y7CoZn3+pYLrsS4LHk8LW4xdpfYZBcDRMxbKKdoxUMSqO4X
KamQtstZdDd9C4F8GjsOsc0tx4R7uGXY6OGXXGowMpecnbRJIcHts5pMDiBZ4j3f
LYsmhxVTOEnWY1uITxkRwXydJhUsQphRXMU32LM34Ax1PsYqwjZwANeKre5aMUYK
ZE3k2xpmrA7HmIbtEJpfevekQaMNyaDL2Oev6UZVgCz0urc9QnnCl7AHyNpOohcA
hPrjh0gj/OpJr1MOoGQ3vlZ+10vcg0NBiiIex4b/F/2aAiCTQu+zkd5m5nBk9twP
3n6j4nIgRkCpG1xSkcfxIQs7rkCzVzBl4qtVCixOyefK4oGtAAc22RJz7Mf5ZMpS
IyXuagY/gCvqe+T8ss6nZezJTs8sf3BSC0apFa4kNzGjBw6xKWzgFelEAH17fIiL
zhCbeTFJFK75q//sQnVX4se6uziIasI1tRt87h5FA0c83/qQ5xpm7JGEwCgpWcas
bAK/N2u81GJISvRWYBTFd5oo9wczX4ptoenyqy77QfuYnObXWkRJc0FBRscgEjs/
eAiLDASHgCOAOvZ6ocy5JwTRyg5fD/1TxRUOdCN2pOHpEwOHtLPBhN+6NKjr8SH4
+cogMpdJ7R31rTxZ5FTBWWxtS8x43OvmAqgfp6ML5TXccpPAgkHh7STswJXl3wph
6nmbZdiMtRJfod7cEymLxozu7tk0dMFLwEU8PUQetR7mncMfHgXBzinSw1t2Ebmb
1fLReG2wA9j7cJqBiRV4/FlUR7qFggkhgro+RSe0fA6GtleEJa3rRU9RmGaDQCI+
pUN64Dmtk/f5jNp309gXeNRmTJ69nKwL3p33m4djW6aALV4pNJHbkjpvTLnVrk4S
06adHDQlDpcP2rbRfK9yc7mZxribCHuopnCiTfxSecVbVWKa2Vfp5vOdovnEZWrQ
qPKL/ZYgaGwaVRY1TqZwgI0fDhbLE7ZD0cET7ru7NkWF/MNiJu9eTGxdRuTOmyTf
v9pOACpMogR06a18rS/IVqXfrzZ4h0MZDdeZzOXKOPuKRWONJ535Lt5AmQB/xNp4
jI6dtHt8obKubsahY/sw75S0npX10d95fnMlBMmZVNYCD2nuWuYwTRKD/LJOiE7Q
XH1eksJO19jXMpDgCaeJxOdcaahJV07NuvPuzqRfBh1cykDPkC24GPtHkQaDyfiO
AgHk0Bub82YppwP0YlwnP8YG5Lv74FBXowxPb0OVhcMfmoQAsBCReFEArt+Qt+xq
IzAPFnDUjz8BOfLqLLX0uZAYTczbaWzLGpiOh+3Hf7Oq1hevcW/slwSLFh1ODPCn
7p7tjRYB1xap40k2mEnwRXw7k6hNAUjffHp1TV8c38uj9+QAP7xR+zbaf7OzzCGk
z/UFjyiXGdVqhhS0Il7u8NU89oOtjn8rFwt6G/1Skx6doaLclJKxW01mVHRVk7yp
/b9ERJFV9HPcTEjS74RWHI/bvknX5TsnfuncwQII+H8Dm5LzCNqBsZRamog8JD53
8PMnYoTxifpVaOIsDW3aYraAbW+2g25qlMNwHi38eFwsrTjM/RYwmnwML9MqwF0G
B6ZQl1nji9ic6hX0WZz2UNMMNX0LfjG0FKwXsx59QS1UeS15hSult3XfiXsxc6X/
v5axfFPWlEJ3UsZQa6Jyu89p0SDQEIYAmsEOSQ7Y6DTthd17MQjL2D0w+al86E9+
zB2tJJMR62LggYBwzjA54XUPblHwirg3ufiue8lUzuQ6d1KdQ9Bh91b/e2mJN4j/
JUVui3UFJoYBQyehHZrClyUVdjxbi0U3s+6JdVCwfP0SmyRMIxAOfOhLR78wU/62
suN6JU1YOJPv+1CB7F6syECjyB5wfbEOZ20+pXNFzuKViikjT3wZc0Fu93Ef67XX
JM/Kd5dLY7PiFeDESxAe7hmB4TWPmETQfCRl+2R4gfS7DqrT42rfQXcGows0Mgdt
pZh/hZ29Ex8uAnz/0aGXX79HXOhqKflzER1MOHK1XQ+kmRW8JLDzCNBuj1pBlufl
71PKC/fK4B4R7y+wBhSL7G06kfKldmPMO1uRaHpJneQ4Fk+5q5oXNJ3wO+xAjBRi
hkeIOFpnosLwiJk6z2DLVCWawE94jz6g2Gc0paJQ5dxEdrigvhIY3REkhKc+OJo2
wastO6WciH5l0fGt0rufNML+QR/TM++/tTXleqTJs8INO48Q4fB11CM3sww4NxkP
Hffuj3Fy7EzjxyifuoE0IyoWhhdv0wn1pVmi152bZAWCE0ymJjjEAb/99KRwxPpW
yCYqAJvPxC2Ev4ApND1HhbpWNYZhhWgYcoMr10GMY17nMY90j3cJ+wyGB6M9qiXp
MyK7H2yftrt2ydsUEwI90OkAv6kxA0n+FlrXYsoo/5CJ0Hq/q/U4VaJPwaI7DrYj
fe/7YalnQ+i8CaEn27nRR2xP1dsalDjjiapz01+PQKfXJAKVDhzjNoOEnX+JbITx
X2z4aDvYGB2b8L1rllesnXGBrnVrWpQUXTkkV4KJwyK8xoI4zpl8c6qD4GChsU3a
I3vci4dN2ZrKG5RuAXduUz7pa074SK+87sMgMUUj3nazpP21qasUNGz53agL1cVS
zGTUX3e6R4barBnlJHoj2ToC00eUqLQarsZyDwHLmOOH3FUY/J59OXAMnp2upmIW
18pIp053LL11XuuV84yqOV0KnQZ1g1NlDhS6oOCoF27NURGwrMhn9teAhXH1kQns
3tPVN+PGACYX2RUEYyxc1AzmElX0TMQZGy0FjLqxol0JdBJl+aKcaoM57JOje1py
ZKgy5DLV5LX1wA1g3KM6FdcrW+Xh6pn76bIg1P7NkbtatoS5IE3H3UdpT7fJpjsE
MW+WnEtR0ErWUnv++QJa7M2GAV8bL8ZXLKAZTnVqYqh898UBj3mlwRoZfuj1SGyN
LrNr9TsyoE62iyxy0lHOsh4JHWuF5d9cy5YD54UqROWV4n96IQOoSsuFUmUmHBRW
9JZzEH6QKurST+t94hKppnDNf04kX1x8KhTF1/fQt53Jgb8QxQNeUV91BkGl0H2T
B+kx3/4IW30oQ1vvnkF48JhzaEqwRjYnyBix89l2IGKWoZwR65FGxxG6sIPN1tyq
QkfI4GbFehI4r70f9eXfYdh1eAtYmnGoKJInWRO6rgqQwOfwfSWCRWRiS2ZGNwoA
qzlufaFlstZb/YouVkJUam0MHi6gQ0uw+aNUi4UeV/PMt0WjA0DlDsZ5iqUoViLG
xX/HUqQc3FkiY86F7xSZYlpzbgmNl9iK8CGq0XXX365UKN8IFeu5/48bmpnfJVbk
D69Djsmab4x1w92zE1zPEDUY0p8vT2WbYt+YFCGXlaEol8MXS+Z+bJIqJTvpWvsq
Xq2/Bn6W0nvUrgUkLiNANuH+aG5baofQL9LDWXC/xhMQhet34qhpDU6bienuSyvO
ZuqQuXScrR5EZRFo4WS/EvhDkpoDDwLAnObacxDm37NacEXh5pg8ifGN6xjTcUbr
pHizkqzsXJ3JlrH9IChIh78XvSYUpcWrktIvgg95JJ3DP4JhK5EWBPGeVBkjDybj
HROJlVKohqKUoomIE5lSCr21gZ8AIh/zOGfdSpoEVGsjjY17CEMiqSRaWxKWdn4u
hYknOd82bngoK60NeoMcnMksmCfsTs4G9pCReUBy1W9GHzAnsE4M6dE5GRwMUeCM
rjbUPivSQQuSubRFQY3dhRJhcjIAj7hKTe5bv4bFoKjvChRKfpGmrESEA3NV7h99
/WcG97DZpv4kE7dZ+2y/+8Zuq1MbD96zCA2b8Wu0CtahENpVGjB3E1h5lrdMi1WA
25odWUw5XxsKScbufyZkFZzNJdOyXLkdWge2MX1OMT+OZ7cDPRRBWWxTS6+cSEG7
qdvPIIIeb9j2VVuuSdU1AUkGJL+OB+6Aa0fkurJGLoPFyn96IEQOoGNsZlU/EPlV
MUA90RCyjFy0in+4c0UUSF0XyLX8esqC8Itisf4emRkTowCJCtqFNnHeoXOnfbVY
Q65nudxeA4t7Pkv/9ZPSzCOSCbYADThfsIKqWmV2LND/kPMXz262nOFtYwefiKrW
OaK8s/Qvl112EdpQpOV+szAl7fjgV9Kyq4s7chM7QO4WCskqHbkbGTja2QdtzVZd
XFD++xIaXI/uRNn6B8oUoYNxzO2kPno7tI/q/w4xEO+76NXZqrK7u/Scq7sUbr5f
ml/hp3SWW6op5HbAQAm9Jp2rUaMdf0r5ubfsw+p1thloP0MXiY8Dl8+I7mFD6pEQ
rDpLi+AA0K6hctQPAbJb0T505UzW1FYGyirm2uoQrY489zN5VrFXIRn28nh/0qPG
y81t3yZr+Y0bp6AY6RUJwRjx8rd4pIRfpJPpPxUqvR0jZsBgXOpwXDqZePgmf+Jo
TEZaFS4NTFXTxqbnM80Ks0nLVQPqYjldAR1bFGX1QxlpIXfhtP5AQeGgjZi4rDj6
LSE/miHpT5v2zIK/gWTmzJ+S6mf/o6UzuP5Xosc/OpC1YBXkigOJ8Rz+RYYi5VBx
bPxbjXYprYPXe22CftdkpRABcUd8l1uU+809/iqfiIl37LPYQ0mlLoifUQVV3fXH
WpZF2avE1W9jM/1w0jFhI65gh5Axv3y6MvdnvS09Dvwxy9CgjSB4lMThjC//R4ri
huEb0Sc2Fo7zpHW3JCiAWLI92YtLr7OekbWdMfitVszJgE1HTnDX12AcSZsERF+v
D5badNo1WNQW7SeZf2upc174TDiotzXSbsnJvlKVaC/Gqwxvstl9SkRcrvGNlWY4
2zjmsrSZ7G5+Id34peoJUrFxTCDIGT0MLTy6VKuygUy8VQFMqcrI2ofHD3mQGSyo
YfwvTVOXjbg7YDq1059Mh85VRcdMTbRnqDcy5QLYNuLNBKJzY+fIglIqMnpdyZvE
1yyxohzsnZ7nS+IXHb4H7Y+M+yXg439+tPozLSGiTNPVwmoIfSj9yLl6wBkcJmtV
RPj3V82plzL5yNdAeFRPUZcnkGvGUYRZiZA3oL3xajskPAg2lcxbCIHg3CL8ISH7
xUrYPnS/pwcOvDHoGPDlkqAi6CKwQkI3+784xYOeDi7HRE1OB1VsDj6KTW4cIP2s
DyONSxOK5CaD8xNR6iCoAaLSr5FXERYb7p9IGDS5o4AQ5Cyhwg/9T6OUxNfHCkoq
btQPaKlQqKcm5GIvNnIqhJ+09YKP30/7koJWMqsuOAjDb+0t+ajsTva3Bq3exm6j
Dg/rfXJ9dJ1VhKhsZrqMiln9lb3i5Z1dKKPjEacKN/p9M1YuTtlDVBRAjBg9APa7
xmlwJ9rjTSR3yNX9WvfhZetYhSaFnJUmoFf7P7ibNjBTF92VVfD0b8PVpZB3moA3
dRTpCACmcfxjpKal52MfelgpKzKDtS45IC6kdBR9HTcQZzMV/EZVPIXckg39WvU0
5xDYo6lA40QUzmL+4yggfjwI14yjLmDdUti8GJhDcVKe6uUtLlwICEYXoTHiTQOZ
F+3bHJWe6KPQhN51cCLHOFb8KZjwmneI215RUb+JBPIaJ+V/bl9LdEU4rkP1sltF
jiniRJ+FuxCpRw/uOefgzoMNELYVusUX3r/IsCVvRPcZeFUamD7Ux2ad8BVB5iBZ
Jn4f/o6DbB6rW7WDx2GQM4FgcvIXInvg1+hpgCxxD5G+HchI2d9mLYJbl32HSqD6
LaLwVugM+APlHbudgp7vUEe1JUoGlMlm/u7r3TT3yMqoedgQPwtkJyOEgGVzrZ4p
r82eS1GHN9JnFXzPXZ3tMD2rNcecLuxSE2gOWGIn2fSCkWIt4o0jdBIYdHPp4Qqs
ymjqYfTR0On+bHRHQyTt79dQFOqcyKoU5TmrX0kE3lh8usP14u/hiv5+Zr/l85QR
NlnSaG8F8AGjW/VzCSFJG4CNAr9MXQQVfmNwVXym2KXyBXRPclTwF1s5Z7cuZ7eJ
9QzZSgS8TOZzv4YndLQVFv7Nmz2som3L6+9iiZ2vLCaf9OKge+C6mcDTO9eufVTY
x1KOgyunPvstXE3B7bIbvfZQbgMysT1vFakLpoEBrcet1ZeN3roVyfDkYDmXW9lj
SSWpCwA8E0AgNHoogIxYG2Kg5l90WxsoU3y7RoMCzg3ZNZL+u62HxQEvvhP8bsWM
SeVIL6eIl/VUNCOExvKsQf5/WZi6KnWeQol91IicOTDsBhRCkLlAnNOl3Y4KHv39
O8yXhoOO4oflrhzMTNjGuNUo5MJAIl3+xJGlQseJmxtfsE4nMXwsOZ+W/NE3c15r
XVlMJyZifdBidK6sHxT3ViSKNaulgICYpMNTVcvTpmt3ZeEF7N/aEe0cDVqD7hx1
cduiQFT6FRC+nlakixzoKbL+re1ayGsxVE7PVGzihEDmgJXObaKBVl7t0PNfECpi
5MIQl3PjA8BTf3421qXOl9M6YRedEf8mqsmNAOHif40IDcs0ELeRJSEBF4B1xIjP
Hjnm8E92s3HNm9bU0B3LAPD5VIJ17FCEk64bllg3cbi7en0QZ18LiwA1IHOL/OTV
M2w1DVv5XFwfezsLgmKVON3/0n4t7szpAzwcDc7NqR+PBD1bnUo6S0YYH4YXx0lC
lB9GffKOzcdItmoM+KOa+T+kOxY56nu+iXkxfEb1fEXl61hVNOiTsfvf+yNZrKh3
nJq0NFsVURexj+s/SgDbKxWsZvqy6E2Rc/q8IHtQwovTheOB2rVaKpj9+GIglgkS
JmGqXhWsZkikKyhVk2HKsx69i1H3zLBJe3BZcvErXFYE0IE63ZQAyO72FHri7c0l
GszmR6Jz+8E9HuMym6ff6RNZTFSJDyUnqzRk6UuRiw2HEnulhZ8vkgzGyFt/wCz8
Fb9w5ygfjAlzmtLhRV9oFE0kQsFcxT856K8+SYOaND4I+1gjw3huc/RZPCUZobdk
hty0ta7hdVXCG1wXCfMtBYxAhnj71RDbo0EjM6jsubu476g+v1gs9f/0bIIT/25R
cFHlq6vK6JTqBogfvi6DNutYHxG9DCcz+vIKGmU4wJVdTAcAJ1xjLuygLWaemHum
SqaRRZiC+HyvDBwp8whfeP+pfM0WCXcgmq8vv4Ghqy6FSuu02ZC2igK/wD7tmumY
JXjS+wiNhFDIvrwQIUWl/s/yREHe2DFa7plCbZO2y2suqEimsK+8IY4rSAyCmHAs
0t7gv6MmxajH0yeC3yDuPykYxczhH6rJvW31eXRJAHYkunfJlRiNAhMFI09J1xb+
zMcVZmwHjA0tOvgB/MQZNgYJTenRZOilIWmoa+Z6kRBi7+wY6L1tQzp15sV3Rg0P
/hEzyXRvtSqLNyEZgZ27RY+IcQtcs/jwGFOWjJC3qC8desBbnLU8Zw9S6qtm6Azl
DACDQELfxZYPPGxGupzo/l4Za17lYaqrAWy/dQudUGQD3z4D3KUMbTXKk+UltQeK
0ieuPwJnZt1UpLMmDiDojuYT5hv4IsN1VC4pTXIRw9zsbTwlNJ/WReJqzyvG27PG
fLKmovDABUWVcjxzsBmvHEOqvAyvvn8SYlgBJTf6+I3TZTeqR1BQIEMy78sTTFAK
8G1o2XtLSy9sLbeUpnBVMG1JoPv9obULESedkATCNnJQUtb23pPv4ZTW0oXcT0ej
aRqa3ERCzYM2eTg078V4aaYoJJBWgxRk8bupd75ERUfIntMXoGg3UcWh8dpnCWiz
Jvf/2jk5B61JPhJDxrAYc88+KuVD98qwFPeJ6H5N6C34fbxSz3OnJPLDmboaC3Ah
i+Z/cPNoMphq0iTgnwfPix0nw7ENbrRBSNMh9If27lG8PZHtJ0Aq+jMmoR/euFH3
uluWywh4u3TTD1mLNJ0QCwSqae8b/kWb4T+pRb5JXGJLNpv2ka5AhNU2movvnmd9
qAkOJYkl9GGr1OZC7mB3trsUOIoMksh+oLSNgb3nlUh7LlBu/P6xFHC1/Q/UdVoS
UpP/wprUQ3oRGA0Vcb478tqnupdhuFJis/uOBStpuXAFeLrS0Q4pZGpzCzN7nN4E
i5G2VT1bUSF3FiLwQiGcKO1r+MrYPyp/vOJZvij0tNOEbouMzx6bprdoLTEDzC3T
IkB4yeJwGw17rhY+WKgn3EXd91iuQ+xQtfA8D71EW4qK/hu5DPPtnpUqp7d+BwR2
1+S0ATuSPQYSjVJNFckTsQK7Dc7ovrfqTNWXPO+xELwblAvlI7ttBKO4bBM0rRvo
B1s4JRLWSvoE4OzmNMQtwv8eMrsCxxjmtVlBAey04SJohm9HUsqD5Dg71z8e9Xw2
monuSmNatcuzi5CYMDQgrqJuEkNwoXzo4wGHZUSxWk5T3takRdQxjNVhSIxtvdPQ
mKIhOqhl/1MOsHzVhjeuHP3MAQOF7h4AMx9Ogl08ovQdc7UP861DZS/ZTLFq+9v3
BaXx3+YfK3oqsNlXeUqgn+LKnKyWwT2xv7YhDaRhP2DTTqDF3087xv5+S86Tmszi
VqtUrurxMeeCtLQFtrRD99RQXseG5Quvsx+7JBLjBi7bzJYlMEYyeKJqjB/jAU1w
RAJU/jK/waZar7mc4asHvebliuehdV+3eKgANY24gtysO8+Ti9hNkLfsys/19rmO
XkPHfggFcDx/+7uF2DYW7VsOjjhxjF8PcM0MYS8rx8LscBXhcfqQpa+vJyithbin
jIWhAspG1UBRbTOrQ1GKVEh2tb2YbHODvhmhGgdzRICypsHvdXKrf5xtmP4BLpU+
wnziJ8ko3l2onkGslpVtDMO1xpFlwGOKT2D1gPvcZGktZsRhtlX6IIlwUC5Vqmw4
pzLH1CbCQEEX3bYOxbwtd851OfP6oCOGp5Ai0vC5HaPrDm+fIXYmBJK2zEvvGYGf
+g5xtxmLvqGSp+ltNB6D2MWnTo6fjypqBDPjTtYUx2k1zpy8Me1Bl6kXorXOo4Ed
QNBAkAghZxhiaB+7dZeVBBountG3AtfdWc9FsYn70oUO4vginZZL9n40VtfQwbSa
NtJz7QZio45r9LBTDq37IXU+0+14KQ90FNvKv5FGp7MgsW9sev/i1JuAHyupUiib
h9PKnfMXmuMXYxXV3e8Qz34XP2ZXh7uhOx6qnakgGeAOi0tqVS7z72tGZY6Fl3bA
kuQnTW2dDDWETyRnHOu9+8P+m8q0AE9SafyMIktlsXqhzJijtYTBCkvoamOXnqu0
/8Qtn2r6mcg3PzWx6yUaByyazaRJ2DqWQoIuemKq5m/r/RwrI+66OhlMiC9WvHpG
rMPLurZhQqMHQ8rIcZcZOJq2WWOSIOEgVWyijm/ztuQJTf2MyusdZtjzicMJPtXH
XuZL6zTMD1qr/qIiu9HuDn8fEqOGvcRcefWjrMzbK61I/8tI/HgRVFyNry71jt95
9aomKHMqD7RM3dbQvm1mz8JXKvhPFp4D9TZZmEnyB8m/InWLjJjOfeL4psdtlrHw
oqI5jlE0zErcz2Sj/71t+cSPVwDwn4GT9S41snR1UhyLFbvCiuR7AvFVla8bnrNv
m92B3xaLY6z36fsJWA1zYii3vLPxtqVWD35qe4EwCRDh1pANpMik4PttqTB0+E5Q
BfCUOezgifMGZ3+v7Mk7ybNmVc+zalgWDaH0+RNl9YSJsf93uirqxKj7uyRCltb+
azAeHUL5DMxviDbK2BtraqzeGp9t9SuPWzLP+cHo3RZnAvzDsYPs87IljX3b8T/t
DmDPa65R/IcIMQvjLep90tbzEfAs7c5oqZD8lHCeOgMYRgR/JWg0CM/nL4opAH34
n63dXgOQFsUGhbDCNqrra/+JjRnTRaQ//Ld+qm6SmlbR1GwOddT8zJ+XaNpaEqR/
rlXJ/stdFpQUoI8j4mho/3/73q27qYD3uIg/lRSdYMB8BfQtyHuKNUEtCzK/xX37
+WSt4cgWEa7CQMPt6JaKavAvOAT5GsNa96PJpVB1fm+400BweazfPBH0+TWs1bzj
xq+VIzRv74cSf6CThIiHlXLh3dU+bAdzHgSUgXOmA1Te9JMsGj+iFGVsPodLus2I
9r1UaTc0ehTzFds4kfSxhgTktuTjvGuIydDSffv52wRwwL93Eiwr9toOfcSxTlV+
gsM4T1vIUMcy0Qe+5lIzlPotv+ZykY4Trc2OhnGI14SBzky7VZPTYLTRZGEbudza
fHdoQbFUDREC/i2/mrKLWAPNOW0volw3xrkPkHjqwHqnoqLshK1qU1xdwLio2St4
xpmNLs6HQ6f/Tl8ZIaxFsurXy6XxVePRq/cu8zYIikvABqRW/X8aH1sRnAf301xT
C/PKzOnXRjqoPCukV5MpWVJ8NRiXCRONeAWu8XVsTXo+d/fNP+t2erTWV69C/SrG
sstEgm6G0Y8okSQAHGVFE+clh85uu6AVa51yTvF3JgWE50TmBaDVDFsR1f4Xnv5x
xeUH5Tkb/F1lNjKvR2QQSFuJbxVJkFt4g9vZ/5Xa4bY2WyFfuR72MmkJLa85zREK
jCq5JqbpIIVoYusbBhbturAe7b4jHmBtybWnKPQRjAIDAJbnriXq3Fm1fNB8us1Q
MR7FLJflnhLlw52ianrFDg/mLCHqZMkEO0GPT+BmHQ0zg+G1moK2v/4lX5qDRUmn
PYCzVoZR3XamwKSF5gYTVXNeoSpunPvsktPgC5AhyeFaNpOhZNPDRLpYQkjvQlJb
Tq8iVSPnrd/dpRB4tHMilfr+r0sRWkPnZ3iDQlnt0anwu7142O5flX8xf8NHZJXF
oYy7QxMUlSmDhhXCFEZJ00Jec6grIdOKrx3ccQYCrhdQ8pNyQyzLivvEmnyCaNCK
IyTgW7bYkji/6pKVtwlzI73Sx/aImEbyoR7Z5LPhTPSiKOncam+6+u4OxqA0yvRu
IuDERYYAwo6/OhTp2P9ziQ5iHeS149xarQ0Mhe2kkow5JRK0cgZo8Z4PVl98NY82
zEAxrb+jp2ZsxMbpOSaV4/nGdeGEcCO9FQ1IFdbv2Bw5T1Cl6ESjf9sYC6STeLte
EEDiDX4XBy4NLDPWQ6k9z4nDTq37ls5xIKjFg8xdPYzI2X8Tu3X70tjM+EGLauak
q7eJ5bPLsDdCXM5BpIAfGEBv60lPOuqBSmJ79KiJj2I8JPaaOUKLLVLc2H0TruRp
D7dhBtNQ45a4H7kEqUvBeuZ42zlgC1lVlI//xpwW+2hXPyDj+WiN81lU252xPvdV
vUOmII85y0vGuLVtqESAm48o7lo+m/OvQnVm7O6TSTHoVtHIzJrjF6RoN/jD+79j
nIHDnW2BWtw54Ef/EL0f73vvqJ/Asu2hcSTJUVw4FxJA+pKSeugX+plpuL82St5P
Rg4qwWB3QKZt8sblFj7Rkl/cp1nd9ms2325OJG4Xv7fgwKEoqfcAzwT8H2Tv5cjg
J+E5Uwk964zmV2BIDbkyVg9ZrHK/KIt5NRg2yaCGLYL+j2loO84wZdpExhU5/ihJ
o1/8D405vOCAXh71WNJzILw8nWhbQJXgzlhvNfIfY1WGRJLzCX2/TKeYM+c4uPel
tCmZWuWLi4AF9Pvt0rJ0fOthSojiGlN44SoUSOFg3+B4pqg6x8yedvaj4xiKT/T4
+/6LR3B5H19+WJAWsrMExGQh3P0hH+PDqll0weRRAWmXP0eXyJouzNogK5qqz/9X
GMd39RhfecV4QZF0IHWWqyRx2zxGgBG174R2CiirjNqxdDXhckJqTouC5yxjlN6d
kl1jb700IZe89tq7EZHIRIhwDQ5Ptqcb1/z4hF8JrXbh8zk6PN0u3J8dfbbU5zQX
dbrVb3qctDy/M9zNV3etPqoysyVm5Czz4XogrAQpR6iZ0iS6ZDFcUHWXG9JdxByE
jh9T9eIRzuCm/MprbHBvnbMLkwKOkXMQXch6iKiomFdke8Ohl0YzinxwqqrnG+Y0
sBNw/2Lah1257TQ3oytSmVMGFDIrwlqecfh0y1gKWZNoGf4t5M+gdEz3ShfU72Wx
JrEv2DbB+tYvlRhsbP3oomcbFnJ//0oHoV9vLEJxJjY6dFLQ2jBb1GQIszlNMupr
FGjRZ+qjMnlBTaVIYNnZDrVPdKyeBGwX59vhzogDK2sAax/mfsVBWK6DkrnR1SrC
xSmwlA/oBrJco3tSpIXffPOracSv73wkXqICF4swNGUwSe7VmX6U1xu1zZnMcoJR
ImDuReBabLWpMUnF7HnQ6TRNb0hGcJ6zgi+o5IpH2NZWEd1HJ2RpMVRvf8vjD544
qJ9uwyxBHtYxKPyNhNzyC62tvMI1UP8N5ZybU8JONm0QUcLZYLEXKxdlXreU6Pd7
tIazzdS36hLwI8sW4bo8Bb3ZdUBUHUlDgO2wRmR1AaIVhgh859lasn7YWG2El2jq
kON8l7DAUlL1KNJiRzwQooDxQ8Fuen6fF5dcjveAfoGJxY36ucGZ4VgDc+HTEDi3
eSlwsSAtk9TjjPG/eZ8P3hoOWg3iORlVaKYxPQpK4eEsSIMecJ6c6t7JFGDvTH4q
PayNq0LJBZhpXMo6woTt8kAgLdeuTM/wSogu7/m1FxKynSAJImSdBch+LZ+gScvH
SOApqnt5iFa/hH69HckmmhcBTSwB5O0IXEWSiXWISI6lWVLNSxvH/OfQ4hDVXBdP
keZ/vK9fuaSmLYvI6K0gVRatSJqCVX+Ubu25n6DQhq27tLXl2CKpyKR2Y94Ar0mw
XwxKMrA/rLbWH9TOWzXcK6nksJ1rZr4DSe6/I4SbqebW4ZqQtMFtOkM3HLKex1+Z
4H0OORuWzlBRtN/S3efnmRQyJVD9R5U4xFMJXHzJgc1qeCxHNcwIXPvxmKuC7Yg1
ALjivTGSPeJ47FIyjTqi8WBKYf+ntIX8O49K6xvQKPdNIieW0FzLmcjbL92MWPuP
jpk015mwgHKXb/9UJ0VHq1IndQ+gglxgqdZbtlM95wILp7uA7JMNgutOgpiCkQdi
+U0i/pebos9b3yFZhlUE7KnGLG5cAocv4nNIXF58ytK1xF9YUYeOi0xm4JBeEEmX
QVeQiDhIrpIgA61+M/XxBIJMK61xBtg5N8czmTdi195KenZHv10CD62nv9BGVavB
HBgJwKkL/eZ4Xj6LpJzeHKaPUTjfMKCZHs9upPrlVwhOnYJExyBkHQ49I8DpZbeY
KYtsL//xbJRxp/JSiEdPEwEc0oFFuoe96QlezI9HIz/EFoi0zJWgvEzUNG/x3ykW
ecg4s8eoMrt9SydEaqfI7lF5ZFj7UQzKXz75sHkUfL2whoAcLMqd9DGKIM90orsj
z9JxY031mhXqiXQnd7iGq16iX3vyzvOZ3Au9zqqwdETyzp4ED+eURViYF/1aqKje
vT27vuDqxABOS4JL90ChhVPk2kVQSacD/Z/8IKTVP6NeSDEFHj1Pzwu6zmR2PibY
LXxJxxZeCUxGRddQsVWxYmR6CP+bOebT1/zXbHo8cQSsxmDhPSErad9c2RwA9vyj
oyPWf6WJo2LGnist668YrSg/OVMJtLUEzF2A2dxsR1rtU0QSUX26FsmtOw3V93hm
m/IfTGrPG7gLXstyfgPSoU8ZU/uOhv14xBAWzywFXz4nfX479YOhienAKEFXCblG
+eDXrpzlDfLASWUyATKoukKGhIXnz29CVgwCMKRbcKQj1eih/qVv4AtOiJaAYJou
o6Bx7cWcKn933gL6EEbbvTMjSFrRFns+hSahlJTuawQZjp0bKjtVMc9WTQSwlySF
kR5tpLU0hGFAgcLm7qnMQlE7li6gx1BYh8Mdk6pPr7Sx+//eZ71tJVXhYM061bBU
ZlNzoRj2de22dQMFMy0Xi8UgHSKNJxu6Di/SI3qFgOqH928+T7nc/PfeJa1B2TxS
cjB6YNJhH7L+I40M3Oz8wpYmUeYkdHLZeb8kgHQFnJTJ5VbN/dyDHjoDNztzw2XV
klDkAVk6b/ey6b3NGkbX1hpMbJUcTtgvIY7exCVO0pLzaitBH4t+BjvkOULOKl/0
B0kOJpAaAiSeWIWh48JdS6fGeh3xa7TH35kk9GNdxN9NJ+pekHiIa4fT0YTCsJc5
vx2+Yyb7K3dnSUdZLiYueFChUFc8h8QZF6MFGIdRXH2g1KvaRxYOFhQCYtRwulYI
P5h7WaIl1skk2ahgIgrD2C6USrlTskf7vC+5ZJJoG/163aEua/AUHlPRKglwGY99
L5g6Tmtn+L4NZhK2c4VQUUqVtdfnze8sTShW+YybjesdwiQgpdLXAnpxJYcMlagh
kTlX2uu8beT0z7Ut+dUUrR3j/cXeKrW31RYwwFksTA5r4sDnBOiKtBNMFHNoOEZ6
SHXRa5XhWsQPGzLPgSMJ3Jsl+vlUBU9vsohmbLBTsxzwMhPtgc+GHpLyuleaF5LF
f3H1g37NuXK2GiY0+4fpnBb+C0w/NVGXE8Dk/kge0IboFbJtzUANkkjcODSFb+cW
bGUu8iTkgSaZtgR71cWWRD9d6PDOvNdFMwBsZz7dBrpKQimSmsnE8J1HWPi3TrZv
a9JeR0c/A8Yi5mjOXIyoizufbvOjP0R6nRQMocYZtQhvrriwTK+2OAU8EwDmNpIs
C6HIeG/oKxkLKDyd+sydenNjLmPXqhoKvFhCERBu+igFq6368neAcM9MqwSTBCSz
vVFPZvwD+7Yo1A7t0XOP52KeSGcdqLSNkXEI/LIYfZQ1xFQhkI+kL5a9kgERIPhs
lziTLrSAkQY8uqGFgvUGYZQWRHvb6vPLBElGVKAbVA6bTrMWUAOvlk6mhl/kMPcp
NKqsaDSR+iO8vwAxfKtnFE6D8UGB2f1kcxuy/tMeGIpKWRMZTwhDq83BY1d30APz
Dti3xbfRcx8A7HhzhVM7dvU+sR6U7TLcIbyH/iHUDst+gdJ4ysxntswhdoOOU+bk
a5YyMg+OGLGPHSV2Vd+2xergv2Zq9CwJpxUwLJYQ3uYz35H6nnd0oiY4rJI+9gA8
yEvQba83ywE+3/vwQ9+aBEkroQ0UKJQCUydVO2ueLUh+q25PjebpRDYfURQw0DDd
aJb86NneRQrGX3KIH+Imllqf2PUd8jdIYq9npquCPtie8f4cpZc4jOAc790L7vtu
N24zhQAzrHX8jbJ4KcjhE3bKjnGhEKyajF/hhlyB6WQeRrenQsJI+Tyb3hhvIHq+
kkU38kXFFCVjZ16oLQz3r+cZ5IffYo/XxLPil9WJ/B6kocbjEpffT87e6Op6m53G
YNSwpC2kkjmh3Rt5+x9lSfK3fKpVAUaiDbWC5FhZUfirDpF0LVL181XqjpA96Q/i
f3F3umfatgs6ZAW9pEVxM7vr1SUB/cwYm19TCb+b3CMnR2tYuQNIrKVr/WseRhTY
3GCMIc9g3TFBJk/JalBjQLv+W7BXY3U7/3qMT7Vr+yP45tADdAjXqjKlW57OJo2q
t9/2OAK9N5+8tDfDGeUwEegrsRsNHAF7gXnn2R/fNsMTEkCL22whdmpEEc2zfxgo
GgGJzoPasvkKGEvxdRLpA0/s/WDLGgZ0vt+Wwv25uRaEKpwy1j2mOjmxg70CbL39
ZiebkPXIxOO6Wt7ZbcMtQAqD5QMgW7L5Qvq8CvdWSJ4qXaZ/4LYlV3YcBQ7En26d
OsNa2hG6MayQx+AceGDZMLZtAvuvGLRlslOXNsPjpnOkFGTQxfq12GBhVaMy5R3t
ahdX3VeqHnB1FYnUy0GUjQAm5AYdMnNZ+M3sXuZTnqQh9wTSTI55Z+YdMXuHXewt
ALCc9pbOCp95zl4tTJr3e9mYJsMDAV0l7jQqPtSoar9BQxYwFMWGTW4pIZRlzHNW
gBXqi2n+2HRPSyVceibPeWyS6S5R9coEuelPdY2QHpq4BAr8EAp096e/Qjn9NCCv
41NJUa1FbdPxdTAJjUWB+kTi8Wn1vCIAxuVAST30cGrQfBCdNHvVPfem8LCmvKlv
R7NybsNdwJuzy/vzGMDx7twTMOU6y5wE5KxtXSG8ov7uwpjvabeBdfQ080A5VUe2
QNvFNGQX8WZJgbfbZ3PlbuUvlObEUqAjHyRUp5hsxNTQJTSkV3L8jkhtieymiQPu
S6Nsd7BtpE50Ju9lvKkf8+vyXL6gQ5PaWxAJhccRPkorsmFz3Y4fU2th62g+dC00
y5Dg0n9cFtFk/lxl8Hc1U87snrTziK0OuuzbMWmuMXjoTc1tBEbzw6EdN4g800t8
8IqxoeQCZ1FI57ByZF+f5bKCCF2KA0vcqlTKsttP9xMR8TfaYJGybjfSHT3ZdMwC
xPcGGdnUB2bavUJhrx6dhkLckM/wbOEo6b2DkjBMFlR7KLBX5/Dj9u7aZxKAJPY/
5jkC34D87ieRYCcB9viQYpYkCinv6PxlBRwFQXB2vPjpkKdGwQN9HRQmRD34Hi+R
u3zibYUe26IE8c7sbOrf9XofFKQ9AQW22bfQAfvYU7JBB74Jcs7gvkrVmklKnxku
582zA/0Vk7iBtHDUE6NUQyl1azwKL+wvat0Txpjm9NtJ0m6ZHIwxzPUWMoJb0EFt
gZkofHQBErtx+hR8FqOAILQyt10OkC+TN5TDkdWfBV5oizJIqqZnq3O3PARJAUMX
8V3YDwicjXZaT+x/H6P2b0Yn2nz10fpnsqERT6kb5Bh2vDu1G8sr5TcKhrQRwyg3
H23NK5wuId4xrTuKrZksivAznD8KQcDcnSTKUj0KJ/inwT6tPzMBbHpsG9tjnDcH
Cw1v0BJxZucwiNoJfyj9p++rDr+dn1Scjh2I7WeUl5ObbxAp8+GrmNAcdhK/kEnm
6Q/mf8XbswSytIQ/K9sPlPrkX+gybsW5MKlYvTqd/dSKp4ZjCmw03wtNjxg3B0gB
cbT4iamiwVKKRTmHgiKjQHC8TdSPknquLfw7refXvpOsucS5muDQPvpTDqkk/mhx
9GAwp5iz1tPF/rSx9mDL3G9jkfmn8wWrvjIvSuJKsEXcRlDkNcnlraRU32wtE3pc
AwRdSdDipaL4ui3yxi5nqA9sO6ZzzK7blOWSpit9CrFBFJbALoHMwhUrhS3krBDg
gvJB0Agff4UhTGM89KxyELdL87sgZ5Fnm0Ya2xAv1MHrKFdZQ61h+PuYJqTWAUBb
SxlxeFoZ0YPFZbyhtiXFIIeNSr0TgmD8p6ifSJCzyi5bvFc6HWxyqEtsUL7M2rWP
X3tLY6k+HJyZOCTQVpHkrHL8V2i1jfhfaNqBppeffGwsjwVjmxIgAUKRuLN2Wyir
1me0VbdzcxTJoFg6vurKDMFTzH2lJ8U04+4alYQc+4yXvNQA9A3Qa9JG4PphTTzP
ghVnsZbdD8+1JyJrZoE/mFzH+EjOCXnyE9WWOrScKmMvUGvjF0PXqg1q5Hi6P6OD
Y44/M+GyYyeiFFp+mLjaPrN2dkAASG49vaGKXQEv5dOx9G2CSJY83erP9m/QPm1J
y0EW7EPQEAHe18XgG94fJsVbkGu1ym1kt7EvzF8sI5F/Xo9eWMZV0SpPqQLwEM2T
Nt/I6tebe6zCzs3DiWx9G99conRewpNx5t/7qZJmkvAjCjXZ/hfV9IQ3DlAbUYv6
bJF2fKnbDn8EYaOI63SsF3igE+VsmbMVbYnTlMvhsnF9LAQi72sgsLel9Z6d1Yyp
LP0kYu5Ay2xF+K6w3W90MM0UF9WEkarF4PQKOdvtzzRkp4hjZjuNofOhIDZV/j6s
6otR0R7gSAbfrcMgXHvpAb4gDsL8nJSQWoyy2B0IoS3u09RAKyr63m3aCB6AeKPK
OBbE+r4wseIaUcZ/lID6gvkFBG9Qz1UxCwW8thFDwD/qkZaXMvkYH9nSilzNck07
oNYtYKW6Hp/FWplrC7PKFpHpL820PXCfqSV5IOictk2Xi/dUvVTmn9PgQcR7+Nbq
kNh/Qs6On++mcVXDWRaalkReb1jtTJeYvCloxAH7nKfxUU9NHc39/oBp+bD+0yZv
Jvyy7lvBT2FgEqN6fYsXBJG/Bhs/kkdP5YK9Xfcc9im95oB+MCgjr6Bq1XvFtJw1
1bUxmyQYZEgOlN/2I0g4H3oewsovFpNy8AEV+hNrVt1Q01wA372TOrQj/vbt3lxw
iBBdeQdrvYehe/rRP67mAxsE4k6NUT3a37iFdUP4aL02nOyLktKdmu6r+KMsyn/8
/lX6d7un9BzvVgic5YrR/A4U/gPrWT1Lu/97dfx3DY45sfpaOIo8Yny6pvaMQpWV
a1r1y8+6fajdOdYMSQpc7Tg0rnNqLWdjmM8RJR1YsMnEcRTK3cpz59MjeKP0KAAd
OTNFmrdD7O/ul+/vtEOT8+AmdKtNOsOxaTJ+ueL63L7ptyJH8Yh9jqB1pKRSsDmG
fYSAPkTzvij9n5Toh7LTuGV9X/3wwrPqI6vPk3u7mOnATvZSaY4e3CVS+ogrzhwS
gIUA5G2IAol4iVAaChKm3jpe9OiYZ6ag+y/dIpGdHLVAtvbK9lcCsKnU4BA+goMU
fk05rOKumuxTNMWhsUwyXvPyiUBGJrSGPyZJlCMAI1UL7Bg9BHFx5lvihsMLFFsM
xnLjl9eXy+nP7E8ymngabpnldZTam1k4I7L22fuq2s0Ynj1BSPRQcF2/GsWt4z1p
6EbR8LwnKOXGN9V9C0pswr4nsAn92oei9YwJwHbm08K4UgGF7HRBrtXxUxSs+Ea6
rEoP/kLBXuIzLgF1dLoAyCe/D6CygW468LEKb98j8c+3I5ZyFhY0ioih4oV1msVc
aUPnN+zADoJuN4EKHHXX4Hv5m3D0qdsEiC639liGQaX1MLiZ3nrx2v9pi+PxWgCf
hqztjeK7idcQZL9c+mnmTrlXQfNbH/+hm+sXYb6EDxkSPNsRIhLuiEPNOoseKAWR
3wxO+6L4n098hm1533wMKuayUe820HSckgQNgq6uMYdVwMNA/0Vj1b2OmN1fKNED
cdrWGsPDOcbxw6E6iHxzdBgQFXPMM94xXb77ho2mWquN2Zul5wdO8JDZ4T5fpWft
jCqSNRRMiibxloIW85W0W3g3ZwXFV+QsYteFiylol8fcYN2cehz6V/iFz23Bf3un
AmvA2st/zSIs4ax39T4fMD9Niab2AKuLZUOOa9ntwrIkr91lSpn7/fSw1WpsEf2Z
bY4VQYYEzQuM8L8VR6XCw/UKAd8uLmveeZauCFopDvpiXtirUI4JLjeKp/0JIooH
O81GF5mYEsOfk2+iXA0GEOIzYgGHU9ucqQ89XemWaimQazDEwcy+fcvzt4BdtthC
WMfp9mBmN2OoJign8gTFPVgkWhtEfgvlGxcQmGj9raVS6ymzlHkQSjifAj17WhI/
hjwtIYi/whkdSr+K4pk/cMCXFEmOFehZfT/MLfeNQjfiFBq6bsPTPGQonqbAAeWo
1EPeUgM42PLzxcPv6k8OCDEgKld6h+EusVc+MyUeNF+SGZeTjcb7bzs61CYELlu/
DBhRBQHnrtfNPdvnDAiyjqYdpQXwGXTeLhUlPbECtcpwK+sR94GgTey8IWx3txhM
nmlkkdo8qlvxTlAXnskWcHtBN+nAx3G5AqYCaVy46GMs/zdY7TMM9ObGXzXxLZSh
WcW6sAxwv2jkPCs81oYvYvVG+oShO7BBYtUyFE1cZVCpPQDbPKvbbX7qrZYpDls+
SMBacw6OxKKuej4h+3tNmY32GJAq4oPvBS6710vMtE2GzlQv0VmzxFsbob8crKX5
ZIoG9fUyF8DRlS1lJQh0nz/Rr1oQzDNpR8BBW+etSQE5VLdWoNXwsE6tvtTYUeBK
mmAyt2t6S9p5u+qzaVU7lxWQEDyy+5YMF9kDrP8Tmw3UngMxVx67JXHizL+6f8uT
ysTjGwM8qvhlxvTUHqgiF2+7Scqcrh83Si7h2YCox6yguQJz7RvGgJYk0yRz4hRa
mRAkJeyUFFETgoCtsuCcyifsr3ufj8I3uJqwxRvTJiaRn1P7/nEl3kauFasvIawH
IxHmbQkbSBbysB8x1jnZFyHpsmJUKhV7c0hl/Z+wUkKRsfRclvl0SHmhuZIS0amf
TYNRx1K1VcUvIRWpwX3Or1cKcMCggWfO8G9OWi5ChhYRh/J9oZZdYF0kd/ACaZXM
UL2is+puDoYpAoWDAWZMbOvjLS6MnoYfMTxRcRyp0aAKIyFFJoOywXYkCCjqKF/Q
vHLmiCDctwWjNdHLVONPhySXJ0XaqklBvqygkfVvqi8D89qN8bi521pSQoYERSgI
tXcLN7NZI2oHIHCeAa/fXkM73FhDDI4+CiFiK8bdPPBIcpJPZZOuiRRAf62IMV4O
52oMSte8k+YIo+GF/zWHmM3lZMaHpNBSAdXrDrSzVI2HJMz3Fd/UzLpDrixI6uQ2
fEL7PW0LXUG+b9Fbh4SNlWlLqt/BqTvqnp9vQZRiIctfAGYyfKpCj/CJflWz+Hc2
5YSGucPchZA1JUb1Qcj/+fRklmZEvSWOzL83Q5sTutUAm250Wd5Ao9KTxLBTGsOl
1b1TD9wuCoHf5yvub6+0HbPo8sxi1mjx6+4xScknrb0nNxKkOdA8ziURgI9DLQwV
mIe7kgNGU3BgZDQImqigEqok3YmNZkDHXo2adJ7Vjyxrl6SL8BnDGvX71yrM+n9y
PvN1VuHP7faVMLXSd0biKkuM8dVxLYkWb9UPV3xzTE7d0aafcYVttxgx4uD8laZ3
abZeRBjFJ1MfDeRJyCreLEp8GzlZSH6FbiK3sqxa70WhTP1eR3kNlEAMi1LztXty
CvUFrO114V6/gpxnIh8LMxfN6McNiUTOj7PIHTjcZF+6LqgSXFiPTyaBI8/lgKo3
4+yUUdI2gPVW1ZPYR22csPKdYuXX0nRaoOjPRa2cillnrJw/4Ygde5PH/bUvPXLl
fis3QdZoxUcmuOrjU68D1qcTuvA5Ecw8h9djrar8tejKeFKaPRxMzV6xB3bt2WuT
t53wAL+DdyGJBPokRcnz3x3Lg6gAfXVKgtab52y47XPfXt9Cssfx8uQ7ab0HTsmx
tMU/OO1fYyNFAJL3Awai6Gta57uSkBVu5i2W17EIQTVM/9PqwN3dCY4kdDRKUOxM
MDHmI2+UwprBLEH8t93iQC2pLfcLUIWxgJUW8I3FT1MvEx7gInh59AjSumUG7Gr+
tEWjGEDNYHBi83og2CsLcXJmLbvyQN5/A0DiiQ5cpi1cap9IzLuPZ5aTKdI9gPw4
YAeAcBN6Dd7K8l0Dszr6viGrauYyUgaygMluqyeflLSaRPcsDLqAqtWiL7D8IGz1
euebeFvLf1NJ1ItR9dBx1s2vZrIQ/fXkaHUu4+AGCP/wdhD6r+F7+pjkMfysRvTJ
nTBn6KLZJhoadzCAlRO0H+a91I6gum88WP1mjjdSXyv+KzmzdTLhB9fsr3IPEFLm
XvPUHCcgl8A7wuH0eJ3yFOUqozSOROrmz4ehdPMBYDssp+r+zp+B5N8ECj9mK2WF
nTdFhIiby+et0oMFD6tvQDOJ+l68H5LTmnsoG+Ef19AxWTdpwX94yy2lY8nfIg8G
SHGtZKbMK9Jl8bGW6fJoQbNy0dtczoBKqaP43EDYndymVGDGpBOLA7DGug9AfVI5
LgkFb36BuX9U3v2Ze9JB+fTYKDPepeu3LgIzTS4shtml2EY4hkgcwKE2/Fq2E2+O
fwlDUwoP9rBLlypvM3110nww7uKsWP90LnpTb4+vej4qEFHpHysgszlAQpOSH3hm
tu2aEpOQwAe9UumUHzZCuSjssIPtUYwrytSg63l1tc0H0i4wK/wUFJJPPzsGXjaA
Fuxfe6zQ2YpptqyLx8icy9cviWHZkbDRwoR7O5Yhr5UXdsrlS8PdGzN1Rb4qXL/x
DwxF1pgkxcOeXqDR0Kt2rQbjU2SXUCPzr7NoDgLQYVbsxysH7eEKa7B14N2uKIqo
9LVbTe3QLYZD9+13yvuhUOBtuCBivmrfwVIOYKEK2Qul6JN1d8JIWzVbcL9Y+wID
n9pc1QHbD4GaB9NppVK6ylGtC+tEvSEmjed2KIpBAla/iwvc8W1EHjyXdp1I9GO8
LJcM6YiC/Yz/vKFCELtp+/rs4lLRqAFS1j/WjWlfnHZogZbh5ETXf3NyrwmMmjOm
zWtVuSyzMhLvamZxkqK/owWvwbXzAfSv27afIqQORX4gY+tkCkIVBfwX778biLnX
HOVDOyMGA5i5ALaOdft8aA3UTeR+ElaR1eL9EcDlDQY1jpvUul94sdOPSrvmFilU
+eedSNugMhjVIcFd3pKeO5XxzknwyNJ7O9Hky+yv3UEvHlQQVzlSr8d9yrsalCkU
yDt/CEd45bLsSLuvItUAAHpdUJ0ETkNuthpupgikb2ZAXiblQ74QJasPE4SAeGYE
tDg6pWSWSIaBmCR/PhhNlu5qpUYfN7OZNRA6KIe6acvBfonDAEj8yvxJkYWn/cF6
hrTOGRQPBWgdXQ2PRsOIeWbnNHOPNOCz7VONZm+bkjAzWHehODLxyNLlCL9Jy7My
GhgqGQlc8kddW0168NZTCuk8ejEMgMzaJ/dZsVIlQaQupgz3GwJtpmzDlfA4NgAe
+2QClLpiYm/U//TKxf2KXFJ4IJFf/poNV9gotIO3TMAh3t9HXtcwOWANYhe/Hyxa
Vt3Te3SXyIkXs0VgB4KHMIZuQDpRaSdbTXV35g7ztGnElhWNxToKx0Pvr2ypfDja
VJFZHbf5QqzEsjqgdWHym22FuXbdox0MOr8hzz17teQl0jl3wiQJ63DhqGbYvRFp
5srcEErYSx3zEPR9LyR0AwDUSw5xr1v9pj7MIgn1b6W8m561T40QrnwqHwa4JGW4
+D6saWEkt3603rOO5pFkNYEDtgEH7M/2NOXxK72SHiAPjT2jIjh7aCNn4oaW1IeC
phq4WGvCrgDcaxzF1xDj5lI2XZXPHy7w+LKBrwfsekMQeUCFYkbQErDD93bpopSJ
Zl5L8fjkeJfIs9j1GvbJmPq3ln7qGUXbaoWPtWfrc5wodsqf2JPTpOMYNroeC2Pw
2fFTzfPxvQelPlf9sRtOdtgJG+mR889IseTH965IpELUO1QLis7yqZx5nN/zcmHW
gkRPaJBovV4PWBhKwVbivp/cnbfFrtmvMbTiR4MWNoGqAiqOYeNlU98S7KcejnXM
Bhx+cSAg1kW52xH/f0BtVwigKlpEE9zH45HvpZRRmNyax3XVDLCtKxT3Kn8PukXR
FtMOIyxAjRQrChnFFXEAYmMzDe0cP/PfNK47utctD8q25/TngvfyI9bNHWgTWzJa
Wx4xlIByUdGmOhOsBbE1LsaPadIGwZA8bS2Cy1WPqR7EL7maJNFvXc02UxYkNFWt
vFZq3cda5kThG79kWRNXtyCV3oRnM+opDxOiFqLRXlCmfhS2ZLGll7OaHQxuaiwq
BmW4Xlaja6UbjLrVOcier0dPjQiZHJuy2gSv825RK+W61Gs3/CtC0lwFbX71IMRY
rdMzEcBAiA+BsKZfjPqT0oXos/88zm+SNGCXnE2XhoSMBmE4i2+Zz6JMUg6WnTIn
zzAe1bKs5A2PT08/Y57/KydMT4MqU8KBty6ctLO8HzTv+IY4VKiF2wiuEtZxiAIW
qPnTD8N76Aan0qLmnbNJBeC2mmb36gNQNgG7l1mwKqOj5qTMB4gbxeoXjHX0Clwp
cUjUzXU+EW4QNM41+S+kFwnGKjsw4vjXF1B43d7kMGjRX/1NRRl1wNnw1tgEwOf8
BEkL80T3xkX8WgBMcGilEm/v+/nVMxV3HEfIRhnrQiKyBFp6+L9lKdydXeOX4J8q
dVSKEZqwTkYSu6/HEIRH9jtEQciajeOlwdL64TWJgOj/5lANcbhLDkfzCTLUb8pM
71gbwxatVWxxn0zFqG2PfL74NgXznH4+fGSMqNH+YZ1xnfeu0WDgb5I0KWFNjLBb
+uyIGxQgw52C9PlXoKsYt71bOYlrQ/fC3kl6uXVNj1x+1uS61c4ZdUHUyoetVZ8j
DvbBVMR5RJ+3yI9Za9kUBbxkj/Tkkus+69/BwPXgAtfQbhqACGSuf2TwpMhYFn/k
ObwSRtuPlW2jDUZFrL2+w0NC9ZzKaPhUBb64j9pZ3NWZ/+UhLOUTZpaPq7y+qktQ
zQktvhigqb5i5vdKfy+NZIR3rwcKfYdTLZUjyH5RyvgsjLz4fb8x2PKAEiUwOyRw
LUaIlyrQvKHDjUKOTNw/mS3AVOtiHfZNKiaX1KMExXeQ1sGf4EsmqtFJdJzHPoc5
1GHJzU8WVIPNsv30OeKbW8UWRhTkTSO9/ezu7vKaS34RJkrjX26SGFbUc95IGhBo
TCW28kYv9oaL5p23mz0VRuhxVJn+VSyBV3NHd9ACWFCGmcqYhTFPzZd4CgOOSij+
gKq4YuNtjeI46gpP53haLq/qQI2RR6L95n7fdPWAF5v96dScOFcXe6cdL3zhSPd9
Up4MswzsOAojGB7N9c4SLdDrHWr/GWBLSW2J3aOtchEsR7L3jVai/U1d0dwA3NcG
EaaIM94fm6+CdTV2LBFUGd53O6P2nMP10vWlPfXp5wQtKtSWLzuGA3GgJx94jp9m
RBxR0MUPf4WDWyIpvkssPjZsPbxVAjILYitHVR6TWNC3BBZg46ZnqHvxv0qyqrwG
o0sAa5Pnemzv5YSVASwBZHKvk5rpqtGduCnGy6i+gyEVymUEd5v373Kgb2Ce9/Lg
Tzs2nbwtp9EPr8r+k8XezAWncSD7+PovLNF5iudQFdSOR6ZipLZx4DZlBZY9H1pR
beL6fEwCP36snE/Bxg3nHw5Gv9x1TXXseJ0W4u21RB8FpM9FkhckRdAop6XidEVS
LQ9V13EcKUAdDJ/B1xYSPbcUYoblzXh/15GjBuA59iL/9QlaorSOOOfrz2ifyKN6
hsB+fU5+wejbMhNlO6ZXzPjohVYbo+w8ndFyc2alPa27Yortd+nH2i/VAyPCF2kP
uRE+TwF66ummv7TD12DlkqDz87IwDChITG71y7/soSAQolMHrT6g36XD6/lcZQvv
Z+R2CNwEG1SJ9+TEjZBhP5lshZNl+9oMQpSftu8iyAwB7NWPeV/RnUMvA21XhRLs
wpjZcy5o+t1HPG/qjQUfSyz3WbSHUs6tV5wmp0yzfxAmwOFJRSU3MZvWpUAL+Ggn
o/FzF3QkSXRGDXozyU5AUkeJDWf1fJ+8SJFblzVnr4VL8HK2ZYuAxNK+XKVbDOV4
F9rDhMAM4o5SxfR3ZG03Ieo1ALcf3LqK0HIfMbuOiMicIZhyRLdn4mVfqhlWlcEV
qS+Fz7ZAtUjZ3vgirhtQdeXLniy0kInzQjGv6dMIdYECluqQCIF+MloLNM92Vy2f
UGliI10KoGn78vn8tzDI/WM60XUfNF3w9mXIBZqtY95q6J6sJUlKLN7NfsH1Bsqa
S45BTn+wczF/QJxrFBYSLX+/ISkF8SCmWzjqeG80Dn8slbINcJeeyrB58yFcy7T9
uQ7U3QK3lcMatNo5TuuVD/zTw3pZrpcGJTj+jbmfZYa3ouIQKzU5j4zlCUPFVYAi
vioyx1qeliNDHmPdJjKW/1F5cF9r2hqiMKLf7ILt9GFhcr4KlwEOCGLu1z/L1537
HnSAfvQaZCld4QKcNCg7cYqpvqMOlKh9VmJvpsXm8nO+ijkoKLpacJaMt8+1L9Ho
Gr9+2fdEdk2mLzG9M06vmRt9UxZR1cCpVLkEIE5RjUbL2MXySnzpDFwqrGQYwarx
0Oo1s2vVdwwhp6gIh2Hgtk3YlEoBsWYGbc7EFgX0HcGh5MxpUORgxGx8xFtkGcJ0
yX1Pcvz7LunHfH6u61LewrscJSZk/Aa8YNQ/TJqwR+/JDjMNeevDNdKnFRc44UuR
5aHMp5UZdZOj6SNogRWKUufm05ZPBFSwscifkCi25jR3IRQ220mOsII1Tf8cbzRR
LvgyYEx6mbyB03GoAj5hSLuNUEJu9e7DF0kuGz2uRz48W/QNKhV8o7jJy1IiicgY
n5pTiLCIKKsQ5JwvGy/4NA6NpRBFxIL7eGzN8pDKZn51zhYl5HDNOe/WJV9kaRGJ
HolGadxB9M4oX+VkEuHATFxJ5+YQAWyU0ifwCKeAFA1kP2z/l7TypIyslY6VTI2A
/s4z+RwDEJ6+RlEe2Xn8knB6qizNGmGMiOhGZa7Ne5NG4etYfZZ2/XEKl4oSluFH
tdiiN7l4S/aTJH+uN0GZ7KFjnERzwabloEE8VD5l+aK4fPghyooiBysQVR1Lo5jl
SmZHs9F0udXRJ6VudvlP2eoUJVZd3Vg9eImev4DERUSK2v4RW3gMvqPcsU60TprP
Oit5tKBsw97OrrO45sqHh0EluQJHvIrzruKIApwsywj4ZDo8/IQoXPzLpyZl2yh2
OjeshLKCEtt/lNDmtMzSY8T6MvFvatvD6a0RiZkFx+PYpNA3efnziD+v/0XMZ1vU
jQEcwBXXGZV5bghfWbn/NyQ4Z5xgQ+40jyCUFV80vJz45nFMAOuoS1dcLDN2x0EH
rRuore98ZcHGAnvhglsiv3mFcKs66m9JRQwoWXu2VdJptUrKQxhlKmnh98io7HZE
1Jl0wdrVL9y+93o3oSsowtLUTeaM5CNr5/8fRW6r/9occB3RHu3pVgAR2AeFEI0y
EiBoGHl6SibFDmHNaGQMgMR/SfaCkHjmsLVSqn1O3aljAvtgMSBlElGcdL51Zc5V
IV/Z9OOchNk+/KcbY2ZsHNvpXfVl4mt3P+q7Gf071L4eTU+nQDHLsnrYV1usiE3W
EHG3B3LpCNt96H4UuG95ALVFB3V3ySq9m8u4ax48bGMZMR0iNF+5rctqmnqD7te8
qON86pcz99uQf+Tfy4uyNM+cuNeg03Gpr0zvWtKKadxIe+As9RotikatJD3cDHxg
HY/7ysColyT08p9Yj2pzkgHckvzT2djheufQRaK6l1PwSuSu3lN8Q+5iGG1FxSwu
kJhoXO/0XoCLUgulaA3RADSeKEN+1Sk35YQU6dbEuXu1cUDdiHsmgnefPYdUQJjH
tKxDaaoXszoWFGorNxYOZ5jiiS+lftl+5Cc5DAGGGOACUcsJX258rgd9Fs6b+iOW
JefK5R07x6A0eNoJZTtPcFiKEP1yEU/ajTjwcDWkcJ/vDY3t8GOHKmqzmF+fL0Hf
PDN+EdmA1Sb1/umcTUPsNYXlAsPMvfptLqY9Z9pq6UkTUDk/cEbxpHnMK8W4mdpX
9gbHdmnp4i0jX61JuBTb/wG86Grq9MU5kN/tmsN7z8v8kAYjk65VPDtE7wamTeGU
SVvV3PDSp+lwa8GSCGG9rupfWtUSNptSwTNbidjqzasgTljL1g4cH0t9xuc5K4+I
5dYHe1mSo1fXOv0Kvp1oBxJll+p5IpcFezkB31hvyPY+vF3/3jRDRcCI2ymV67XF
2LM2FzltR4Jhe0ngnoBU0PU8wa8fFwZGIcRsPwiq28Migb2T3aP8OXKwn1lReFNs
MP3xi1qWGQGD7KXCiHRW9m7S1EUzfEgXmc7+8cN5zhq5mlSKhgid2+UxF6JWkO7i
K5kmuwa4RWxaCo2DNxtCgpAZ55lYDD2zMCoGPQ+n11U8HBhw2XE8lKWXA3SREDry
YJvh50Nawz6grkUdlgOEskMAXntAULBnvFseUi8yWCRjBL1QkVWAAE97P9wMJLpS
3PsCGpDF8iMpjzY6xxHsFPv0OmrwbSSzoO4L6HNefRnadmUEDzAS0Cf0z3ZMvCpO
YoECeLxwXVj3irGwiRB2qHYx/Wg8dWM4yPEgohFzTKGxXJSOJU3IvSp4Hxps0tbw
ors2h7bauFCxarg1vidhJgei4QaIMFHVXfqdAcrUwKuMY89x9F7oIGKHgNB916H5
uf/Wo4D6v0cix1DHrIOu+EKP1e2UDSoT2rPyOny+C5ruCcOA+qn5gEM/xBAR9Jr4
wy4n6rdOk+B45Cao4kswCmlohi8oEajfOT8a8Xwb0G/Ecvj/g7yboRVC5+ac83yI
ifIyo+p9wIA/G34mUX4lB4XYSVFBeWGDwC7wbnNmK1GF/3sEQym+Ei848fQjspsM
5Gney65IjmotJHHj2GJhNlLunbCWuOFm5DYZfBD8kkkLcqNXIMZIjX9NNSHYLMVC
DBIb0ClRnF95AOVpSBGdqJxPr6fmtg/4Y1p92IF79uD93GhgcxRwXLJMrNYwQ482
a4QgyzV/ip8G/vwfv+p16IYwrwVTIkVnFd7ofEqzcaSf+NZELoxZeUkeqKUnYFyU
yY0z9vzLxCDHFk2TNbuYdYqkPW2XWU4QCauJ+eR7yBmZULy5rw/9HmjoR0FvtNCf
VpcGQq7VZyqM5oS7/hXwRfLvzenKtBxn050mFVXnI+zkK2MmIYJOXHmDMw0uqatG
DEzHsMnxCxc6iGUezfXtLOo8GOUBhOiokKJbRhkXhcLz+DyO64SS205OYN0d5Prd
8EmeCwTIFXtSHReCdiuXXTcNckj998bbvAQ6Df/+l1HhkJOLklcbZ9HuW+8jdTJp
3iGXfRihfvkPML+qUxCFXqMfugwMKbki3PSWtUikmcQB9mwpwxePPnifK2RfDDvX
pRKP/11lMPUHLK5LoBUJHAqYi7IqyEO+6pYi4o4xWfUiVqbhmTZ7zctnHM0YK3km
PPtfynoYTJMAGaJgkxGm6jUlInZWllUra/vNqSBFkhYClxwhQ4Vx2e9zpywLOyUg
o+SlS2b/A/+IBJki3HslHOybNNmeI5fKTouH1vUR5cIHkw0GF2QA7f2OqvEyDSbZ
hKEZ86Z3Ueb+eK+wx1SI8oZO+Neg1c65DxeBSpBO+mH1Rm7uskUNBICBQ0gF7ZaP
Nd2MXCzE0//ZW5ECpm9J2JKMqpGNNvX8jYfVjWmBreilwUekwpnPsMUOMjUErNr2
JdikSgoEY7q11Egb/8uXQW+/+hKjYKMC8ZzwjKPD1ttjdYbaS1AVv9BWk8ZqEraI
5FeACaXpwppiYHaqWb4rRKDppt4HSP80IeivGENOx9cG/W5ldcCN3g7P/iFq7wi4
2IafEwVv3p+0/PE8pcdHSx8PxFAWGH48whxCkd/Pl7s69zixuwHyX4xzZZNo5gsL
8CVcTUJEtPwEBXokb/lc3RhK2lHJ0HjAJHrAENK01uNlR6vHDUSfXsApoZtQl4uw
tmaBUg83gaWVP1Mm1yuUFEPEYgb/1dbwPD+/9EG8G7OUu7sNJKLFltIEj3au2xDE
aYD3LWMZrcGDvD3UoAHY4sPhZFMPae0q9cYEd+yZhOEcRnKH8aslwjS1KhRDjH2P
N+pi5NyCgaBjrXxkJEorZ24NyNKd4RMIYPuKIzGZvUdazu8g8SA0bzwtdt4V3ax/
Yk0FTiAJerOaerOMA9UI/L/msxDb8liRo+R1bHHi3XvZ5PkoXxKYpTekr6RL5uXP
TrIiAVCzM3lJPahqwYqSq5sQyAXhjO01++SxvSucemC81jHLIKzZ/FnSSpnlabvB
3h3X9cgaKXEJktczDK/Psgb7PnNkS0djc7YrQX6Qz/vDpaW+Cyiy4eIEk2FUTf6f
hD0pktSffjqG4eGxzKmZVyC3VdW0ax6j4Yavj2bNOYtpV+E2evinV8kZuwhxktVi
SjXPrlf95T31QvFpjaACptW+AbU6hqc/d8Unm7fJq7AtIdzhuEDYqPPH04JPnu0M
PB857n0kfCtB3eLn7uZI+E4FUEIaKzeFr5kdVa7b6PgM2yqJTweQR0ikygB0s5qM
HSMQa1ViTOXYotx1PnTCz4xpEPwqzEmbaT2uzk/eWtdmWxxbOSraVPzjjvtQixYx
zfWtynEbFXf6NRQqhFA0zXn8ZK3mAJSujTGnlTPXs5gDHRhLpvCxhiNnINuNEA5+
dlHxHF9OT+DiZVU65e+z5eqNu3/er9vJPf2gETBmIvsjcAQcmBMHLpZrehSZIwvi
W3ACzkSivO2hyx0jrXhuzb4VXiG9P6U2jHAsbmbqtmZ5nftakgRLuZvE9DhxfMoa
D7BZj2ajPuhJjWP7PetavS80fxLOHIEN907WWQMlJDboYZBX2sZho5vFYTW1Oh0J
nuq6qRgfN4aYj2TN388NSqcNleIowIiwWJ9zcUNo2zHCxvhGKugkN16LatPe2DGV
FL811jTUKkq39uT3Af1Wp4QYeCS/iYu0xLmkwLEW1eXkNB6HN9C6xfswRJqVXhU1
1uyMTeyw1Opz3zgdlomVDoMg0c4QFPO7OjhujIhq5JiYvw9oFHj+GoVt4xBaD/Hw
iTLSsLuQMpf74UGQcj8565iRlo/GuCAFPO3Ta3Hk9JFIu3+FDEEMBwlpLVD1hbuW
rzVu4lwkcFAzBfB81WkKlVY1vFKMOmQNb3ZK8fPPTpH/lKjqBrooDaxSSvpPkosa
vKqB70Hed0Q2kzJtP7NgXFFw63FPMtzHUShFK+aUAr6BDUrmPromX5U25kBwe/DP
/5KLkR/YtVlL63xvsT9wWGAUHwKXPoMczLHB95Z9U199iV3xb/4MqINBj5NVwx10
5/dOvHbPJkDdPjnGExtZ8N0ktRUtNNlneptmnn8/9yyE3iq1r5VC7183oSyDXDq0
8AGz2jQDSIOJBKrrwmanO1nn2w1ZyNg08Prxxs2kgmy6/+7prbBWTwP90utKljWO
W51dCR9wFGZZJkjxRVRbifr9FWK5QqBkJVOLIfxW+d0uQLniMRYDcIYG3Vlc9kBe
h0YVVNH7waGJ2JdkdcXJeXm4jPjbeGAi5nYe+q9YNBw9gCF0Hcwr1msodgwLkNhH
Y7OQariBSecpt0Ys002pTGShVlhBz09BIJ/ojaJZf1aFU1j3/Zb7igUzhhUQ8Xbw
gB8OtC7RMDbriXWaJE9lQeNY032anmIN8YhQI4RFvaY7o+SbSB41YjGsJhATpRjS
OvE1qSv+HlSFnVbItKVevi2xbfjdSrmX9Q/zNpNhTWbjWMTBU4EnpywzS4CF3Rll
uLp3D74Kz+RmFZ+LxgBYKn0eKTGVUUHT4G99nTd6sAHQsBVzOGnCuNEHuLMw56OC
VQqYoO5DJCMtXsa+4VNaIIcuOr1FStoF6qb2L5P++ZqpydFnO1yr8Zeq/thBcElo
clXEDLbC2Xx/WZd2RRXwREcfemYFYWD0k7a4OqhLB8SbvCklPghviudyFrSE/Yw/
tv42kWTLf3Qtl3suWqxOCYLtwJ26P9WUluo0RAv8zaVHTNqjGG/bcor1XInRwelR
D5ndoMcHYAXxW7nVIzY1sMh2PdbM5kFkscxwgDoq6Fju/CsWrf0hgPc5bSy9jSvX
zcbCjAkfztg++7bEVwO89YCeesP00+viooYTVTVen+umqzEkuy5u7yexD22HOQHH
mmjHs/vES5l5AjHF8+DWEk8n289ixjygmgOCe2d4Oubhn7LFWr2NgWkPE7mh23Ix
x8bRtsgjHuAvYiiy/rgPNi2MXCUhHP3rkUDY52AcwFbbUxI7CGcVZne+bh37JI8z
yZUjgFrwbSauWiSUci/3HWZww3ybSXGRojaTWHSnERKYAtQu9RSd6gG1I2lsa0lQ
WhaABHXrjHOzBLy/7I88hy7LP+ZsVwvZ+Y5/JIlR3GdlVoxgFiBvmeZ0a+pUAIVJ
yAf2qfzi6YSYo3VPeQcZkcXpVKcnc3fZJ+UdrVGFGteQjivf08mhYwrYk9h6D3q0
zT+qeL9QEQLnbJBz0umrQtBrPlRMnCBgNZTAXJ3slYSLe7Uyd6YOEUUQUluLSCIe
f3qMBKxXRWuAMt6U4gUNPK1JgXtccijHP5YUbhSBeX5ueY39bh50FF/6IL+EXiiw
2ls49ka+XOahAhajhxwjph6JaCU59YqSIeOwS5+jBQb7xWcPlYHChbPQNwczVdy1
G+7zKyZWikesGYd8IUzQ5MTShBErfW3IAqEbhCCYGVeBTZuiPjLWZANXBkfgwDtm
Drj3DT0vzctuXJnxqmGnwJ4ZngBJIlz/Pe3Z12rPgfrdjv0V/R+FQF92dmMMzVC5
n9GCY1cDNCQBRVlPEoimTZRcO+5/TiRj3Fn9cvvlz7XkuBd5SuCQkZqRw2WA6+78
U2TB1Uz/1P+IeDnc9fmCTu4H5MFBRQ1x0G5NdQZdrKuaueQBw5DpmAadrpauUGi8
pveGvpdVZGhf1W8wMTIzhjVPJIR3ytuaU9qpoNZeDuh3GTdoP76XPLGJyxKk17h/
XwNPDFg5Oo/3Ld4r1M0i4jqIcrMpKYg41ohxkC4vlNxMCNua+Ow1UxIenXYJFgov
cmroL4xmHzMI4w6e+rIFAJb8Iqm3wwTzuQkjlyh6ugh6gRKzsm2UccuAweK/KmMm
rzBAx7Pfupe8/3ln4Wvw0rY569HE9p1F5TCSzCiiMPGc3arhCIS6VBmpvU11LwhC
dG3eMoZ//Jh9eGB3vdBX3kbYEjYW4a+MxNQJEJHqIghYAl/qPV8lbPkoz0Fae/V5
N2hpDH+TO6IOrhEziBN8vD9LIdeN8YRsAGHbBOrejff2mam115AH65kPJ/V7oPWP
pvS12PR0Vvi5Wnw2hTE4hU150XVz2cQMp0vUbdLce5QzTexGFZ8EJr5rsd3dWtKn
ZnCioF5hqQRJd5plVy+GIogSl94QB+XXyyMNykyrnGuBInehONIeipqp9ixHu9YU
jecVpMglebOPuj/gH2MHimRLlqwAF0VMNukgSGm9Ni+WfBwCCrzDxKsMXZQdnHTh
gDR6usvI1smvGgZ65yRZccqNhlsm0k9Cv8FT7x6XPLLeWAm8cR15HgDsKznR/BiY
EZxcJBDW4VHWKdMXr6BzMk4xgP+xnTA9VA3MNYjFW1Mnp2fWW8WGTWVjjNVOwCBq
i/aaEbB8TBd2bGraT8ua4rL6aD4M998M594AncSQYxlRgVEj8QocANtsWfB9euJu
ARthzj/fhHLLa36lmz890Ad/dXbrQuUDR/6rlM8QGUEPQv1kh20BDXhNd57EOOb5
pvcZ+dEC4gPc4iYDtj/mEUUiJQR/qt1cYGZIvyXKHdLitZKyq+pwhY5v2kTuZSIB
JtD58hrgCziQukaG1K777YAtd8/z8w0DwaG10ejuir9mRz4prZa2WuKc2RlhJ8Bl
VeK95/ETVoN1nqSHg5UUL+0r2I06zk62GysOBiysp+P25tv9ryazaDbluR54i5Eu
RAxuTpG5UFKwPtQ1CcWACWVOxrVVqT73n+GVmisplZJTqaWWPQq2j8G19s47ocWW
E32TxM/MJDbALP4CoeZW5sDSqqWClwByLBItcIxvcwgOHwFLJb22YT0bLwyYr2ce
oYTJf5u/F6TGHh5/TdA/uZvaMnGWz4/dGNWL9ZPUQdk5pj+2fVx3u09tAUJUgwO9
XeZ1cy7ntEq7XOWnuwOt0fwEuVph+j2mH2Vc0CfXGoatg7DaVUxsKngNz1why9e7
5w14r2Pkw0M3BgXFeGXs7ArYxDsGmdMQwWzwmS67nU4FiDw5hFIX2Ry0ILOaxOJF
07NyhmEinf8HBvhMIG1nyObc2Fr2wN1NU6sGgKj55pa+py56l8V/2mHCrZaI8OL+
NQJLvkXetBtiAL+8tVuhH4LjHloR9MxFaOFONwo/+miduwxHVIuc6S0SkvscYWQm
6UqehgHcM6fmImw7f+cDsNTI4ukbqkFLx9IppAcQaBWF6tw4xwJxHOieTXtoeDj9
2SqJJI7gBLiGEPEpHe7Q6GHV7XR8WagXOQNDEfZ/gstED+ZcDNXwMEkv9x9sit2F
Jw/6ebFiywFO4RUF91rkfv4ewADB0r/I8mT+bzOCtBoHNP/ctgZjzOXO0qnn2Vw/
UrWndaPWp6y7OS4ga3hVY8Kgp8QbJ8B/uacfgy+3uCWN/OYH4CW1T/Q5p0zCsTMm
C9ryG/dYE7o6H3MHzux/a3qAFXMoR3AKa2yAHtPxhMCEup/d+4YXHIHACn5pj9P/
7fjhzfSoyGgS73Sl5hqTom2riHlyYNHs0YivFCbgPjJZqTpmSoJqCqpJE9PiQ0kG
b4z7d1Sw4chtm1j182IktcGvzkqG3Tbj6WbEGX1bsCpqs9M9Apcxzu+x+435C5rz
V6T49ICS154dfwB32uHc6WCSlhyIfVcXUvbfvB93QrQGwqnMmUyy2Q95v02u15+u
EUzfGE2wr0yW/f9n3+OUDdPmOCJf7Yzip6wPO7U2vrFjXY05+QfVA+T/9dv2sd5k
m3DxLKKzmnXWaWGWf/h5mB/J9a+8G0vH5YDvMlpd31goLvNDtSdcGI1DHpCuRS7p
BC9XuzwaOgwGvTo8bXo0oP2AOAzIb67wchOCDELPW61tLpFvYc3dD63ou2rloUiZ
vqBtXCxAo15PyMQQb7SQvYCHKfzaSc56MIheThG3FgmXRKU5J9BgUs4L3f2kHbZf
a1uN5I0ZYfTeDUd1Z1OlMfuM0NcRaC6vvxtpmltpws6n0QBm0AqIAFJs2W78ATGh
Bti5rcfQVdjRkY1XL2bCf/uDBzHJM0KsaCu1294e8ZoI89tF0D9+zPEuE+doCS/q
EMDxBsioGuxHZDOp+dfmSfHiinDk+smy9WI+RtydS/7p6/F9mDS/x85AJIL0Ewkv
YDRoTdIsojPJCwU2aCVJssVj5vI+Ac9LTQmDzTqN1U+P0cc4gnrOhMEnwbep1gQ5
eRrvFyZc+xYwh0EPIM6ajv9QwSVSgJbIQ5Qjqn8H5xS9aXxQhQ/xi0liQbLBqRj0
hULzQ0HhzULg8KYCNiSeO2mU3pmys/RuXmjYhpkMDqAzHTOdsHkl6aAcIBW7UxrE
vH76M1qDvtd2sWVo39u7w4T0X5VtVe3vorV3MWPDv0T7i06s34EtnOiLQnirvPI+
Gl7yxCPy5mPsSgMKLRwoytpbEoaJ8PJAHIM13onrrayPyWXmPcBdGDylG5SF3hXB
+VnVe9Cr3hODOSrylffmvL3NgA3u0eM+75EyqK801hHaAjpPenrOnJO1H5+nxAd5
b4YliLY4GaEO0VamxJdHj/m7WLNLLqdAxyjrzIjavMlzjz+y0SBvAYsobyWcizQl
QB7kP4Ha5E+esIFTDOnsDNn/qjx0tmXVIHi0QTb0/9scO0nZy8IhwcCALrKXPo9h
PdFAHdHWyz2P8saMWwwG0zho4OP4sRZoguXqd2yVZIwxzmVF0SBvyO4X4Zn8a51c
tYj9S3Dar7mgK9h5K6Jp9gFQJONAQPT1fWWgUSYLTihRZdv6UrQDRhJSYyQvLghB
9rFwHx66kP39a+97W5n2r3xY1Yp3bTm4xagvFk3nbHZ5ZoIr6RCnCsJpmb9NbTJN
y97aORWeO6arXkNtxvhlaD3onl30D7hpLMrHFCaMNy/Edc2O2mpajkyGBA7qFwsh
8XdA83+MEuL3ES6w3SP74110J43KzhRHa8hE1JcHF760twUmo/WhXo9zDJwbneNk
eEOvNyvo7BoXk8XUEisTV+zRhGKy+b/Z/sf9bIBDOoXN949VPI15iyEtUY1W6vs1
Ut5chLM2tf5oZ517XtxSkoDW1jeODG/TB7owZ82AbB8VGVVMEBElKUnB1icikucn
lWxu9cY5wC3JLbcT2y4Gd50tOHIvWVAC4/AjTLi0nE7OI1hJF2UzR+qmFuTFD3To
kHSSD1Jc9Eljnd5ahjZ6YA1x3+LdNi9D3nCGDzBAT9UZRux/h3ufKhW88fRsuFBt
Sx1DNKZ+SfqyLqIH4g6hCOXrtr8/Mu6wuL/s1m7PRF1dCsNEJmNas90OCZPIutrZ
Wv0FQBvr5HD4/+NexPvafifAL6EaHLgLE4EQ6i0DNpgQHP7suRSqNdPKnYwOlb/N
590eVuuKonPFaJAZAbdaytXJbXJllmPLL2dY9SNSJ9M+yMMALOCkszjM045eiXkB
UeX8V8iorQKMp+vPZJoI1xgWuYLU8al3di3liiGSoiJpxYAmSOhikK6EtYHOXepN
yYtkMLuC5mu0OMBuoqupiAKFKi0J7RFYB7mc6YllwyAd+8Pu9q7B0cVxmyBQN5hU
pIgJIsPx6tHUCYh4R37O6e1rj2d3pD+BHbWfDhBhCXatC9otF0b0lOb064pVmyw2
5aQ+bGjAx8igIPtPZm1F//vm20uleJUlT6OuK3Kt8zdJt1u+SQssGCJYhqJXWrMC
zNUEgob8y2Wpnoz7t2bV0AnSEVZx50osaiZKe7mXKsQN2ezXZjP3H2GQhIz8Qn6G
HlVnytH1VGEX3/KtQhOtiGicL7RHdAnYItNzJmMF0a7DvGSh4dJg6apOstJRTdvs
lBcDbZgWM/QDrq+uC43Ux2EfkEUh5TOtFevsxx+j7bcW/cXcXcXSOqAnetcPNmcf
Qy7cXxlb2ptDwmzzOhmFNgE4fZGBCuqHxS3qQDCPf50LE7BLitDlw6PkBYDkiK4j
xrIZ/O3MDY/WzPNOD1KeME9YHgAgcxMk5DykV0erifiHfmXrvNNq/9E78pj9QKi7
eogcqdq0PMU0DPHYG+iJYrAStRmWzTKN30Gv5HjJQMqLghpUPuEw5W3LQ9cdnUce
Ef/M5MUlTv2VUwi0mNDha2VXt1/okK2j1RgoYxvHg1dC9xvt0c8DWnmYod1kYa7y
25nGUsPSHYprSb+9C7l+efXufqWKKDTQ4ZuwxAGVQQ+XxkFjrQFgn1WKAm3Kdk/c
TLWNpiOy9kbx0AkoXTxbQwvaQAPr6DkxnpkIwN750ss60yqgIbClg27Ao1vSdA/E
pQBs4uI7EdWgxJdkF4AOz7KYEcDf0HPTAHxJ4jjefMvowD7CJTgTINt/qTcmd8X4
KGz463Q0XlkHmxBijblw/FoequObaHlMXBejs3n0748JTeoUeYg/H4F6KPATEnOD
Kk29Yc1y9bnnAMJ6wKNSZtT9lG5uahAmSfcaJ7YX2gIZLnAMmEAHgZY6QCXodjcW
qrIllnWsenhunpHV3S4zVyGdQQLbXBvQX/LD7ppUxvOGkewwI4xBZ6rggHNg6Zbm
Hbz3OwUTbtwWgtZrNUsA5ImmG68T/gSdhhWB6kZ8fXKYBaeoCWRwKi5dK32VXkx9
3ljaTAv3pKTBWqujUWDv1SjRiFPWPoIhb+ckBCGtU/dOYm8GSMU4y+4GKO9/1jC4
GAmpC0jGe3Pz88lUq1yQGEBNfftbBA5/ojrtDFZPi7ZsJJJOrI+DOTvjN66ZDld/
LIh7l6WnoA2mN9vtgGngqGfQqLsHjwZDGgErO2CgMFfd/gt3gMFa4bHZyXbTLhIE
YxgtSQWBo/szpUA7qrssEoxG95yd7qw06dJ6TrwI1dD4G8viXm2Puvt5l+8Y1Y0t
7LAnD3P203r7FfnbXCcNJIogrcEQitsQc+GZZ1X/573dCfwwejDV7RxMFcYt1dbs
zkS3wsBaYR/dqD55tGysJFUfvMJm22OCClYenD3nJSCFF3MZ7T1QxIytsWU5ZCzg
MXb6r+ETGJJn7XJ//BWt6ozCPy3xFHFfBQ3BFiZUFANMgxlQUfQzAQyFnPh8Yjnv
M0kDQfPBSC084oCiVPnL4bw7psxeSKA1gq4EExtf5Z5AEc79CdHjNoeseFUQyVeD
4yKqxf3MlF9uiHUmyRKG5//aJ83rBgtLvlWMXUhGvPmB2fvXbyIfjJjZQOpTrW72
+1jwntvFZaXSyzzbsqpl0mKvitFJVDvL3Uc8TGE50VbC4hamYq9mYuQd6F2qpAcB
cEenocsljd8OjEJ1Sh4I0S10Q5Q6ymwGXdFDQHGoFTPKr4vZ22f0rR72xOxZ+/RI
dNpTSoOjWhY06ZnEtjnWyvXlQSeJ2MqiTsrMt6VkbXOYGehOlysJjYg80UyCKw3Z
X1UwLpJ+KB6FU5QMh32FYDw9A/C9j7kh9w5xPIK4vAdUr40AdhiJZ6lOOV3u8LQK
ynaD4u+l0GTU5H2yTtFpcXXuNSr+/4Rp6Di7MV9vXzYPD5OyANqJ7MBNVOhizvkZ
UA4ZliLo4rzU74IigB4dwQjTBc5FfBXwuCyM22oTDhNd+x/wYBKO1lzeojJTnRSX
e0lwQttXJvpq6YAAYHvwI2WDer4l1amC1KRFUVOMrgpHFWYAwV3UlGcex2yim7g8
IrddXvgkmKbJfJbmyLAP665EImXqH7MsKyzmv2SGcd/71tqIbK1tNtbwmQ6N1hq9
7pI5CQroc20GfQkgIuARWtL5LzOHbj3lH1CAYehhMIvPOl1vgx7/cAtIB0CiPINW
g3lH9W42k4WwilqSCYsQ4QtQL3pQm4EoR2pm4FpY8TofvXjvLeEY5tEyrdsAbf2d
tiBfEl7+TRay0DbNesVG2iC/pNV1QQD9OIg4mrRvuq+KAucf7/0l2xGHZ7RmTmUg
PmZAv6ZZzuY2xTib7zzoY6oCb4auzEjH+dJixXqIsLP/SAVoQBiEwVvv6I3brkW9
1TsFxkPUw4jarzdGV97lj2fay6IvH48NXmhkkXydIi+AQ/JQCENxbJQnjW0mO9Kn
CTEX3Ol9mpAYg1Xkn8An7A3yPUhyrwvIC6l+h9Lx8Db5HbfoBwWEbLPVNHrzt0qF
2ICdWUUvgszO0OgAtHcW4NpxxRFrrkuBGWNbkniH2n1QWS6CC8Tp+B+WdPLwsLe/
wP14Pn0Cu0p4caeX8bp22aEleZDosCU2Pq7lwmF5GWb+cVaTUB7chqx1pOYqSPJx
be86o0sxksKkfjt1ibKrkIexO9LGK1yRuFRs8Moiux7DXUvIjiZQb8OzInv/bnis
5dzAeVOlmbfnu83ajMEGUka6yB4C5HwopPfWHkStBv3LQJ9xyjwemZVQyr/94OCc
acFnGFDBCWhVf7K9lnfd1U/A8G3Vm75e3VvYqALZNd50s+mWTgje0AuQd4fdrgU7
yeS5DgrvGEIRkMUXfAvmnI1HbtrFXz/870Gh7OtXtcUdX2Fmn3HaJBGbq9+3yqwI
B8+BPQ9pv5i0QOa2dQhSojFkdMICHV8zV8dnlMjqSPnOvpASjWXZ9eQzYUF+vNng
CX3CfJwuxUZYoVohLvxYwZ4fRQ2HkYsxkBqMfuWwrWjCkkopr41LmXj/FVSqWuSi
wvIcRiVnAzkyKDehP3J+mPXfTA99zdCSU5Zdkk5YoxwyKbQJE+NnWvSWnquFqaoM
KAJvik67BcBZ/QMArNE+DqKy9ea10Mnm1wSRBTgfToWqJr1LzPYOlr1HRt8QTg2f
rBumr+vSwYD0EaHCNGYsqor4qelvUIE8X/5UEpcNZtQdgARTtaJTVaae4u1fqizk
J3qR2UnInWiHc6wwvgvIhNIgAv3V6I0kUGuAN33mqzkaHg8/XSF7KiqSncYbOYQN
9RU3FoLlqnk11p+7flk85fFg6yp6ARYqLgG/h1pJMkZTZTynERTdtgVCAsvviJut
3qZL8TDZXXBj+GVNsYSb+F1q3FWNn/GnMLqcjYZGVN+uzAtUNuPctkwn4U6KJL/W
p3g8BaZJ4wCtK05DvUsHrrK/NiIBXQoy/hv7boX5ptEk3YRE/QDlZVYys2JQJ20N
6wzwigho05yTso0aGjuUBAhzyLU0dPmY3ze5GaA3VtkPnKqSJPBf6D+M6qBC8i2G
auWr3hvSTpXXnluNLZuz2tOOlDn8LIqUisjx/p2qxOiba6zSGi1MBSRjUiZD42F9
Dd+lwdiRMeKCN123ohb0PAK3ENqqZrBD9wFfm6kA7dzLYPyPyHZ2Q2BWqjX5S7tL
k+V7O6SB2YQhAJFWuo3YpnPkke2cXB/0yxhBzs9gFMv6KVof4wS5Q4R7XhfoLXUq
mX1UbxUoKkJNvtZFYa0OXy4nb4cQOiWj5o7X7IrA0uSSHVg4U3F7z/w/6EXRUW2o
M73ta31MFkVhndjw+wuKJScPpri+AHWvOyc3554wsKHbRmS1jbnxe+TARa29tWSn
OFtCXMHm64HEykEsMDiHSkWfc1p02gXsj+8HKKov7RgEQQtD9W0QRJinIYcEpgD4
naBPwYxltx9RBDFfBJraZ4lpWHqqKeNq2pmR2MBOHoOmv8r1VvEv9z5kHey5c1q/
/otWZdf4Ln43P1ClpdfOOtIXlg9jCPgdvdmR9gsuKj+tM4BPKpDKmGb1AskTdStn
VJ/U+57RLHKOO6ZwQ8/L6xlvvpN1LZT74fFvXNTGITdEbTFHEALmFNcVFN9MfLms
SmnO3QryeEpNVbiUsFryaXwjXkEG51dgv4yXUWZPNyZss3RnVYbUhP1UntgZ4rTI
IYUFP2k9YyGainqEJhQhevE1IOp4F2cNCfxbyYIvJTJTJ54lOmPfU+2ivwHUkusX
u6+10f/4iYQ7U4Rm4K15jl7fWOlWpzee6oYELB+Y9Xt210KBY237nMZbpL8JQBQz
N7l3VoAenE66l6ThS88/a3yoZE5wzg78I/cOTRoZYiCeaDBFfkka3uxhs4YGk+qo
2OsttIiB2NoQ5ONolZ3oeqYMgFbL9EfZctQQ+Y8U7x6/TOuSAnefgTGNOleyTCDt
8BVV0VkbF8DR8CsEMrOaydpcQZCakz1wse7q0vyV6X7jbc/XFONN0dGpe4PKVUS8
Jd+Bjhwc2waM8oP5GUJo/7ES7ZQfVOtDSJnx3qqXqJQK1wBBMfsLuhveILmWDQ8M
5N/fkliue56G6qmUT3aZVe8J52M/lFWNl0vrG/TNrZBAnWs+RdrnlctwqD2Ogvle
T28y4Ze6GdGHrqzsjV+wjZiAascIUlUCf8TqWKgyWLA7DgTI94f0rmc9UjLiEOhC
XOS9DT/oNXZvo8mD907S0eXhQl6aQC/uf8bVfvRQGvNipanho80ZxqMKOFMIDuVp
g3csZpCGErvxiBv2JObZuy5BdseA+kmjN1zcvY3ezzp+gXL9QigUdxNEQrkNUgyr
7WgKQt3rCah4vGjRTtY3muZV8L4dOiKVFij2h0lH/os3aQCrN7TmcFq971ZmFnxI
PfqbgK5GXK25JqmHHCq/PxnqJrqvK7pc8keRzrv2BcqCcWYDYgmMUyNoVaozAJq1
xaPrPX/1VlubqAESLjwYvFNyRoQA6COwZd6uqAasDxaWj9z9fvkJ9j8S7ugxKRod
qfV6UcI/E/RY6nmq6eaMAlgaHm02k6OzaIhlidDzt71yZJuimPu8yS7Cb7eEW2or
UtysIpY9Vhgj5NQASUA04RhJAKTgrvOoeHHGtTciM8j7NKleq0ucueIC70DA5KBE
su3KdRIoMcjqZ3x9qba+z5/WFruY8HH4FOyP12yy6vthBIprwuh2NTUduW23Tyky
eMbts82yjMBD+U4ZkFftMq7+6CxL6g6knGJzOyKrBVdmtYp1p1yAmJnl5SaXZDkG
9ZCzP4TMOWWdFoj9sSP//kIr93A1ruNk7BnPcJBEauQi8AFMFmTZzke84M6EQIkO
DUcreS40EN0ioHZ+CcRCY5WhycRBd8hc//yotUPVc8pa1RmNJqfDOama0McWkm4b
+DUNz+1W0Nd3yLHRWK0EvtJ0MDf2twa1bdFbwX9zKct0BSovFjsknjCVfjA2Sb+s
renIv6Ab0Q60F0lbig/C6aTuKLgNF1VFJVYOS41rKcLsNcxxw0MCbWQzMQZCMUA7
AEQZqxqKqyPMEKUHIpgJ/gpvA7qpSaKRJrnK/B7yNluKm8tbB3qwm3L8LKkoAiQe
CtVTm8GkzzaXdq+DjlJ027wfHQhx5VXiRZ7tXnCACprc5xT9F0Kl/uiUY9l/F/Z0
cyxCLAZnqdf/flKcyz/UY/2xQf3mF3Iph16x4Nv70tYy/s7A6wNQGqhNktKDALfI
e6MD7f8g9MeDq9rq4BwZf4LWVZDhvvMmnJG28dxyT8jg0nCc2MvXvSX2ysMcW+H3
UhcuG3nM718MLAdDGFHsTMWp+P+3hhwSuQK70epqrlShHmdNgjFRSaS5oKLPqKO2
WdtNf9JO6dkY+/oyVL/uNSqgybSTMpM8mbKd3QzBkUThIfpnALhE/sJAJIOtobOS
lkw53B1+mHnr0NKKmxXQ+QA+Nf41phN09iTAl89/iECw+TJ3+iQgj/PFa0BJGoIp
Zqd7eNZvfn8e24jnOlDy7qgRUNauk3loHavhDIsgMXmWPjjORSapDu5x9PhgWDCt
YTumRCwbkFlg+gsU/+DkksNRVCQvMuGueSzBRlUMaEGtA/2GmlWRxp6W4MN/ITcw
JSlMm2t7x+nwvbSNVfC5tPZkNf8m0jcPh39mRkGWWqpO4FPhixC0FTaKEEa03f/D
8yXiOJHVVwFLUcvrCaSvo9pp3gLHH1dVPHqYJwqdLakBMeA6lKQdcvS33Yvsip5Z
AsrqO6cqQiwzl5cJgf1xCilbob1ta2aiCrpk+bqA52zqt9ctpCeWJBogNxKgiQ9i
X3NAATtmELm2HTC4tQAlxh7gl5aBeAExlycBVXqBZMkF5jQNQNS2dw2wjFZDoef7
dtbeLFX/rBWax74fqB8lYrN30u/IUMCMEROkrOrOQj2UpMFRaxKAhwlNcRO6Emga
EuqAHpBBlZnLYJ11KoFasQ7wpgYTFrV2iRhTX3m8jiaK2SHe5RgoRNRMH3LbuzWT
5vJKT6xRhISLqA+b1HzsX9rSeCbs7IOLd+lrjMTSD0y+pAiLCjZFlj5oDWaG4PAe
94tLDE+itsXpVTU7Oft6/kcINRPBe69MUYw2qK+zDw5GQSroqPPmS5ULRbj23g10
K6dhHBjXCpowL2lGr01fHmt4rL86cEvege8SYng37fMaDsjBtpfmnynBS0plMi0+
WaBqYMo2BOkIhMtYv2MUAdHSltnVttkQX86Zt/NVEMc6gPh6RKBuc7QYkkR5HdU3
OcrDV/QUEOTtzqfNuQlDmnCStzGfyQVN1d04dMKpsTJoO1deSIwczA3bAi23VgqO
gdlyesJfBCJG4hWPaSgmIoFjbeBc6KVIAX8+ZuZoN5cgD3ENB/WiojqKDnUImuBn
aasHf6JmYZzNZ9NkgfRCEQKkSZl1DHc5XZVRXBSaFRG32JmXaFM+IX6Omm4YMvH/
M2A7XwumU9XLjj8vw4KXsOlAGZi03x7yw8/omX622n9TgrEJU746eAfFE6bqWfGu
oizX9XsjUR1xPPb0a7wB76Sfxm5bie3CScw0GWwMn2vonlm6jxsla6Fl9WbKYscA
rgh7P0K08q52bVrOY4G7v+mxlyO82xrJ7aYfeQ+okKpnVc+CzFGfEO90TavEQ+6w
KB0Mi6prdDomKQ3si4P3NJ168V9uG2sQGk+/fyr4WfJ3eFQqG3Whw27/EBmLKxwW
IohhadCUxSskcIkJ164dI0c6rgr7AXkh0pyni0fnlFL2epzKHPUW49pkSMTyuvyN
TBcHryXyIkprTOJ4mW5tObsPFYf8VaoFCqOzpFeNV2torj9p4+QLr9ByBMa5Tao5
S1LI+0HBAai/0B1aZBl9UPmnbacvUqO/LQlY+0z8XL2ejNe1NlHvtk6V4dzrWsyV
AF78vbLh1jNRej6i3RtF97fjCQJYAU0du/F7RyMnbDjNmwauWAitUnEZ3jcJ2Hx+
fE+pMCFHJ+gw+I4T2/46DpyT9ZRc3Rnb3p/o78XuW26F1J78rcJZaOp3o07eIv/A
fuSF+GpX2m+Tvlg6lNrenUmBku7Ci1BQbvnKzi2H/463rqv8v3mbCZ33iqn2be4u
H6v+jENC5J+k/+lrmzytwCm5A5F++w5c36yaMpih8iVg8bGSsYlc7ZMeDu9eKgR3
kF01iHhBZ3fajIYxWlw/7GCK5E2enyX6wUk7xiSVH/ZuTZwCDa6qQD7mD0h2Q9AF
UpBc8t/WWRkWYgFyW7bQ11m9bX+8zP0a0tke4Xd5V5Sg4WV/8rRtDGWKC9aVZD3E
zVTAG2F1b+djmXzbfW25+tkgp4ih+5wzaT1a6dxhH9QsomT5taGlxv9r+Va2L8Si
gEhl/5I9H9sAXc6o2we8Bwe0Q5IcWQdZsnhVTwoqtyAicXnFDks38PeoMZWXwM/Y
7CNc/VuHPx4gb1StF+Mdsa+6yHgFZM/lj22Q0YyFti9blOMKC5TeaH9+5683ew4u
X14uODbsYZgKo1aDUaPmzZYBG0mrKFqr2mej1uQCDeg+C02A7dHYZ8ri+z7H+3H1
/YjIMJRHKx/gxHiLXVVCjkGIEPCN7vbnQ67/K3CzTpo7wHfb74TbzEEBUiwKgvLK
gKvx+rXRGd34OD+M4N1ZXwi5ow6pSsIpsL67kBXDRmRLgGzLdfondv46hsPstyUk
7WphAUo0aS9q3gNJAyihSfEziZTKwIiJvehT25CIFpcM9ugv6tJtJXE6mibWRT3A
s6h7kD3TJYAe6bmVqwWWuDunFFS1zjAIWKgOmc8h6zD5fj01RX5tzo436mTzqAvo
h2kbtl/6GwGrkvhvJJpfi3vXw6syhB9XQ/Rb80Mi78ZEKgR64V9iAqXQJzkwohYT
NhrZmOGFVKYfDMC2NgEHqg46Vz6M7Zfd8oJRgQhA7+AuZktGxNLP7y9YIyipGAs2
enuNwTD7OES0TR4DY/btPcBuH9OWVLXHhveQ7tFtnXZGMdcRSK1JTbWZgYqtPPi2
iUeX0Dz/dnOsiqTb4CelYW+HSNFdaqWy3L6Qk+UYu9+uV/nmHKnU9ow/7H+2AxyB
oI9LI76W0OnXN6AVhwq/Y6izhlg8e1aRQjZdcFOYCRVnTvKvCp7iXmEYJBFtO49T
hdZz/FXdm2uxXAElpKnhwP+UEYJ9tJ8fAQqWKXnT5Ffgq4gktRgm+8gdE7xLQgV+
Lp0m7PPd+51g9kqxhwteZWGqoV7G/+uWhJ1aFOJw4GVOXxDNxJQzGnB7UWd0ss6z
hdnGNlMkvgQ6UmTQ9j+FF33sZ6nH9inIjTPv4y2Vxt/7DWDi3uqaIb2TsqAJcp/5
eALbUQWE/MK269OCIeprGqRyX5e18+C4uwDWJSIiVbFv818m/1kpaETX7enUCjLa
PRmLLYZHiGm8EOYStRLh/VJymGpalbvByg33j1hjX9QbPiob+VPsm2As85XRHE3A
TdIRqw0WRbjARqb+QwfHxjEvG2ZdtO1JKGVX7AUYxZif/YZTvI+uuN5bbp7F2Und
+BnGpRywpZXnBqAR1j55c/a24C69QuoWmghfB3+T7ZBeLb/mlrlVQpioKRSMinuF
RkPGPPJeVvhaGX3e9LweuaGcNg/jRP2+DvPXIozralqex5fUJmZ9S2pPIBzTl8yg
Ybh845Y6otKGly0uK1NK2m4+hPmQKEC/5gLPPhMPPuHUodxnOx/Ji+sldilDepGw
Yqs8MZkroV+zc1fsO4bs7QtTsUUU2ERbnZ6B7Z5PrMO33Ejn/su7WB5+/fX11Lf1
wEr5R6i2Tp1YWre+4OPgTeC+wZyWcH5TGXY5OJbSy7v9d9VyW9DxrF1QtCGGOUYq
HRn51JCTxXOgH67w0MQWPSspxt+dfBf3mZRhVBPzLLG2avJaTmFEHJi6OXTUnOqx
SBfH+4S6Qw0TVqTeDt2oZDziFzp6VJ2y5b0QU0kKqErOyPD2ccaMg7BtzEr4Tnf4
67BqbWnvs4taIedaSDajM0SjMtd/IL5puK8i5R73YuEdHKGdkjN/1wUe2PnfZaKJ
gXdZjq1L3UvUbHSZRnfzmN+DM9LBffPZbi/87iocppjTBnLb1kG6eHcwZjNo75ro
S3A6IGUs8VvNu8NHns+5He00MwREherhPMZ9oQfoguxHj6GheHgNsmEs8CXjRPRv
xF4AQ9RK0rq4QJgqSZw73/qrY8I556q6vTfeFtFBpOgIGTsHxtaAr2EQrgG4fOYd
xahlZ8CcZLBEksrkC6nAzBJoPdmmHkmLSXuCY2N9OfbkpM6uF4oea3ZcObXC5Aou
dtZzhWCB/Al1QQxVs4kANOfxBmaz2HE7AxCNspAXY68i2bcAyAqQlRRjphuNgs1c
9kLDnZI9C+RCbFwx7YZTeLBWNovNpbTGy7Gd01mLGpDWg6dEILrBwpJ+S4guHsEB
KO5Of8PH4ZklJpQ1VYRCZrI8XMtcPSlLDUipo1rHDZ9doh0Sy6UvBu5ZUUOwrGK5
m0QSWJChz7ZKggNLjxgdf5tQ5w5VQ51yepAh/ak7njQgRRT4jFeerb5judSV2geT
Iwm9k1/MZOTOfDTszyb9pJr3Yfl7oYxUcG3sm8bok7EKvlVCOl1STWYcXl8X8JBd
AdvGjSeJbaNjfl+fnFB6Ph7mWGXEDhcX1FR76lJIJRLL1ir87/6bbM3DKf5K2nAr
ifjqXKN6Kot6EOPzVZkjpWk8NyMX4nyY5Ge6oeYXeUrd2gpaZhqdDxBO5Pbfp6lg
bCTo5kmNHECxuhH4K+LkkUHcxQ6QG2lZOfcXuhMGbRgBwlTJOYD5jjwBYKQesInQ
8WopTfDC/Vs0mS9ALNqCFvHmu1hy/hqVxqSOwquTK2cVy8Q4XGRfGu4rZ/m4xZOO
oLpqSL6CSRJALHq5fNNnLOSokZ2C2n8VJh+TePdgDhNZYWpWZzUBa5FGvADR/837
XvhlGT6kzZ3AvQcHtL+EbLRhEz1HOAL6ThQHlPc05QX+dzSMe2oqYW/Hob7wopL7
tQrdvaBWup0CBi1HUvrf9qM3/eSPjHcaDK6fX3FasaV/XNnRBSyxnuh/tbFmUa7F
+PKw5IWlHXi0FS8FYyE2d5ejV0pM6XN3Ri1UtmJ9kRY2MLJFqR6uA9CyCT7F79GI
sm8Y860xu/gCCl+E4ZsRYekOrwYnN4o9rVv4EG1BKZqCo4IfmpHUDGH0xWGlK3w/
cxgruDmLP6cdbR0McrI/pDy8YY7tvtuSjxElFLS6iSzpIeIp1wkdUlk8N0rRnnMU
6ICTTtnw88vqLeXFlXPLzdoaOx0gWfJ4fhA4VLLopPaslWArHXfvDnN1NAxn6KjI
6l7K14Efz9261L3b3FeAj7bb/eg/2V2yLeAI78BCYY3Yl4zmQwfgdtuz13Ax9vjn
NNEcK0LnS2l4ZihVCpDuexQYdaUA/o2BlfbQdK0udS2MF3x+ZM50/kRExnug8O4w
7EcG8UPif2D7D9dgrcw+OwyvAJfwrGqyFrBDRfuJ/pVZJGk/cIICgMqZDnhXVQKj
kWz3ZJMkNsr6USm3lwU1CzgYWEHHbl/NF5LrI6IaYniSVCGmZGBPMWlo0/qz5aaD
IvEHZ25YnvelwQn+QGBW8QDncONQQlNHrABEyqkP8WW6m12iwakd4m1lxjhEpERk
Plgd06kmNc+oCvo+NTrXhFUPvJDQGGMIWiQyVZ7pNr+m7RtrRE8KwImLEXWwDIS4
tajYjd8tkYIZw9qhBKFeGu4OYAAf61k9p/Wu9kbSpWb0itozwJuAnzQ0xEakVqh/
865nKEiPzD2HGDaKTkr1ibLFDMqLgwXnycs+RS/pu3CheL61JJi8qlDmBdu0zywJ
+erSOrzhHSxp1Pzj1I7KTKfx/H9qJnK6TjL+mBfDMVCdzGwOKoQppKRWndDFVUP6
vCV09z84NVH0XraIJx/TX1/XF1zRj/LSvpzz4HrAZP6Q//aE3iVpa5QnxIXY0Abe
YfDOXdeSB5RBL5NhuL2jgr3UVixHQF2SeVf5jQm2aEOmd9XXn5t9wWQra8G/EIpD
2cc7+E1VYEJke2RPyVH8iATfWUzpEVk3kdmberfTFaHA53y2Jceh0MxZn+CULkpi
l2fvSfObF/RN6aL2sUTNK7OUBRuAz01Nt1X1A4ONF53DlJHRU5j6KGqlJ36C7R81
cHH0orCMgTkXH/2qDTzZNCEYoz83PiW95olb0ZyV8/RHZxuG/K2np5jAAYOEzGh5
uOqEfLHnooOjEzYe5sdAPnmfCYWt0zKzdasQg4OKchuzf83mALTZW6X2P4QLYKiM
YJWj9cP+wsgjvbSA2CbZDY/FeoY5bTzrgUPsUGQXFc5cdYosuWbLhJTdyHSr3+CX
depgFx3MP+nj5XilBmNfc8NS9eEnkxJL4JUcgV+dQjbLSMQJ4x8yZu1d6vFYZ9L2
vEjZXgIDwCm2CBXJaXR6GDqcRp4yNn3+bk0b1laJxgxA8nrWAi0hv1+K+3hbHNli
jgQDRVsHMEqncXff+luot+GjPMp7MCWKOPD8XXVC2MLcAJiTQ9pQrkE3ZTS6fNmh
nNZpbZLNPOJ5i58wuPCTE1UTsL3hkFcfIaKl0zetk0p9GfRIsNOydcIy2PMZHK/V
xOogiPajHqpA+bTBGft/if9XcEHkpZ1gpU3IrZg916Nmm5v2JAGGDAI6ZYoQydd9
bzVWdUaI5ZuUnH1z6vg8hf8l6biQN6op193GvWxqKJ7yPmMkvDfoB549wLWWIT6O
qmQAeXy29dtxsbPU/Y7Q0ekVXG4GTEG6S+xQqpwtX0mRxcSG3YM93NexbLXpzTTm
eCAasNfrVuTwU8K3UVx+1NXxBHiFkexM0RJcMRyiegoDDh02f+VlZ3JHYIze6UZi
Ur+xz7xrZV4s3jtcN7qL/rb4W77ZMYZ5P0CY7hgA0tlEJy3e85h/YHaHEvMzVOm2
A0nZCMll1SMkaD1AbDsC/FA3GnKa5IZmJoOqLgf/vz+BW5SHzur9PetNgQpAzxPO
HuqHFdrSMDfHNhvWzKfStzWugVTaV6DA+kHhrduqKugAthL5UN7jc+Vbs6B9yesA
GbO5NFIVR9lEmhD2IVcrfkkgFutV3x3S3REmPd+HnQzHDtWFhWW2k7MzJM9zudV9
6RzyqpbYVwK6HVq9nCpYS69kjBXAfviWjSlezZ4u6haO6Ady/OhN0cSoZfXbO0Ko
6nP0l4yvlQAmNQIAXWvgOZJ05sMx15aCyRHRAFfP9wL2nKEXbmqmlrDexqjWRy2O
mks5L1QffKJfAH20vxQJuRbmz+KEQ30ZKPZNeopzrdbBXR2UK/vaUJF3OC2FYPVB
zLiTGiVsFoEXSCIzCabUGA+QT92cFV9FDh+d2xjzpa3Lhm2z6v8oBvDxjSJaIxER
e+3s/JsDhfrqdh3TpQ0jYUmcncDJTqPcRBdQPKAUJIEMrW9dIVZWva8eQG9aCjhQ
JAf2uQC5CsbYckmuImuvmuTyjprjdTGgLE9zbP8JHHbXyUeQELn1Z7aeCr/Ki5f4
KOZY4BbqtqXrfo1rLXqwU+hAhL8G7p5twI7N6z4Nrvu9QOKBb2sEVOzghuGJx0E3
w60PwDA82CwVAOMgqsUirdBHUQJruLa1X2QKquDVFOPSfId0UhtWd8BC/jCkEkkQ
VRNjd5ch7CBfF3KNsh1bTZg2broXQZlKVxdEOlBF4dwPvDuVeKosWbqxdreflPdL
Lr99Kb/bm7YXFLbX8e5wqSuiCjUVbvoYlYbyDz2dPMGVOSEkaArqBgHS51y0onof
uojwZSCim+Q/EOuMjsSYoZtTAWxk+T519D/BfwlE3WITrkBDxWYrUzQvSI3U7Sui
9+9dK6M/yX1hsrmiFohIfoaP1SfbF5FxSOk1XS9KtQn0Yf4Ve09r8GWTOt1IvuIU
0Ss0y+cG4RzUGnDEu2RXBKnsXjzobyhWXiCNauakg4w2tcQATwPS4yDR+HWkMpWo
We5BxutbTpqt0Q4b+WqSdnqMijNWFlwWoShvKpV8QIWq8Dl8EcxZ3Q6DpXEppei9
g8IfenNwaC8CfS0868Uf6sDWQdljwM4Dg6so58o14Dp15fMG/v/csmgbxzrotuyX
G/RjwnzQrWKgpo1ReVPy34mYD0IkbyU99fWBY892Z76QhRYLUl1P2keT+YcK4I/o
80TBnOXjMA0pc0ybtG/q6DNhUhBfwsUFOMD3deuk7qiSBs/v7Hgfw2oMPQHlOiBN
kWy7eU67ZoH98srXQhTKi9PUTdf8tQTkrU1kzCjjbvdIRR0bg4b4U8nHXh9S0MWu
r22hngsNPdroTIDfZkeN4M0hBJKIomi7PeFBCQp9B1+n0OL6UWL/92rXYY8R1Eeh
6HIDgOFmfPk7myvN50IwELNqgo5ZsCFHPpRoPY9oo6jchkmjBqnkezAGiMYYv+1S
IseFF8dly+Ya+E9p86odXViICtJQJngdoxzYkDEj5sCWYZRgp0YAc0G2TIEuqNOB
CoucD5eKT0qZ8pEwZRE3s9taMUWrovmVBTr7usFP5qE0lvTpSruOYEVFEeg+jj7c
a4l9c8rYGBd/3xV7tMIlRtXR1uba1P4jyTmL+v7VbAUVpBeC3aqPUA4EZNJY2w3P
8GkweXq9tP7tqrAAKnSyOYbl5FYipAxs9akLDCint92pqcx2taoLCBIsmU8QU0xY
ldzgkOGAsJzS74YkAeG6xlSLSDtYtH5ywExhZNXPA/4TkPMuzZb5G3Om3F00mvCk
uM3CZXq1SLceQn8Vf7llp5j0cU22l1PxMGY6NNlR7DYP7rO5taDntniiBbbAL6KV
cLDPK1vQMXNXeBCTwHuokjWCk6ocAuO20lM8GkSGdQXz+ArcobKdXrztV+K5X/OL
lAQ6fpZ+8lwycwtzbOPBx+DYcVMSnNlu3/zfq468209BmB/HhnQDvcp6jt3s/Lqw
p3I/au0HNLiiVAhL1fMSI8bSkQD3XjOfMfsVHfc3ghDJz81PzUu3TAByl2DagZ8v
OzGWeW++PipDVjxd0zPJSsZpSMgw/SwV5c0DqChz0v8Mx06XEyoP++m+/PhBBgrx
r1sFrHBRLAs2B8NGjQlHrXWuYJio0gHv/JI2B/Wl1lhhu9nPg6nIFnqZRFinBSf+
t82IaFYqMutU1JKuaHTibqdFIFtVFeu5iMWmsr6lkO+/TU/8hxNDXB7hRl2ClG7n
zyN0Ib3nVRpfS8QobqhP7vxShHzTJUBoP2mca7ABvUeMoUr5mG8lBtwVwoEE/MNe
JcvAJA/KgvfQd97kdxQbCWBXKpOx3jFdz4QbjADRZ3NrEJZ90N8Z4KPemPf8BKQw
u99hK2XvVlZ2+eNVRigJlbtKjAwmrcvrD75NGZ4BPfgkua0BGECet/d7kKjCnO+O
hV8txHPVl4QzOC8uSVOVFmpfVpJJIxODuQVFPUrwQeecQmSGKQ8Co2brQwCLrDeN
hu+kE5H+Xfki7TByHVs6ETsl/KKowbV0vR1HvhhuKZAJCVc8InEwSAK02cJPHZgB
k7BZnKEyJjg2TtLNBxG+QSJ4IV3FWg86L4KfPBNgxHJ+8WatWmbqm7QU+YC933Wg
yiAdu6uHc9lwLgcLFlbF3VZEX8Qf2bmPXwnE6bEWaV9SWFdAdDeQ1G/k9cecfWpS
1UXeDNz9DPrXl7NXNpDg2p8ZXl9Et8oOhbkL/c6NUIpkwd7KbubLFmuFJZzjxp95
RlNVzn0J5DJLkSysE96ZEf62MdTC3chS/HBCJxZi6KJ64udjbie8HrKCk4tiXQSn
+gunqYZZm2hiw+KGkdCKMUvtT/wotfgmKh6wydhQx6AKreF9AO0WcWy5NGna1hYF
RiVoJTWtSTjhtZeVzQZOW1I+vp57OOTSWW+qdOpNycV/4iNWqkkXW/H6Od8FOMDZ
8yZ71Qhv+SiwlDseZVwrttqybtCkccagaEGynRXK91f1EULOB7taYkIi65/H6udH
9AuaPGyVt4JSB7JAvsC+gCnHaUWFoaFJJ7ptvtarnjI7AwZEAZjHxylcxp22mQqk
cfzBLHweKqChuf7L/E38QsBwwVOvQp+2fDEe51SoQkWNF92A6JAT/j6+fgQCldEq
LRvAFAIURu2LRFaKq3rFnyWOOLtJnLuCw3HWpqLcc2wb6Eb4b/kTIaRJznWns+Hy
UURqrqDG5SziGICXE0ybcsuqTRBUF75iqj0RVRQnIkzdWS6itfRWyt7eCvVJyvND
n0RtG/ATOcBL8c9CiY49+vUO4egKBrK5nIJURoX7M4RXkaka2IwiNA1D1TJQKX4N
Y3FLNmjf4Byk/eaIoi8K8yTrOeh7QdB6vJ02rukk3l7V8zvFmaioMyQFS4oOBIf3
Z7NYRfUHvwy/BWMl8Jx3C8DuuAzEHtmQRUJUHqrG0iPdRONiy0vFRQE9lG5k0+sh
V0lfaUssPlV8vlOXwOf0kJ/GcfEHgUdI2rLBqWU9jshXsl0vRcPJBLo1rUsgoRF6
9+ujmeuY+lOR1AVc5Ij03V44iFx6vBlpNWNeLwueAuXBYPCMam3sPzczD3aBVJN3
jdaeegdAdbgEMbATZrijXrIufeJ6HuaCDli8xR1osqKUK6kPZIhE54E/Nl0VbMD7
clUVNGXZXYgXIoYw4RCdXgSnrymWJxZ8weP/8AvWgycEzats1XZmpJfqdYKyj7o6
XCiWfWpLdjLXu4gzSw1f3IiDZu/az1oAGZsZDby5Gma7Fz1U4zEzs6MeUzCMZPtb
I1JUO5bETCYrJJejLDCDdGhXRGWhtI1XL+ouyGKjynkLvHXmBSKUw6lkPdhH7V/B
HZpcv8DZVEP1L9r+nntJwxVTKwdVUS9wjidCyWv6UqHh4m+jWcgCz5ZItlr9QGb0
haq9IYTDSDRS29K1NdXesyrx1mqJpzHwXLN3EP3wfG8W6tlinC3R8rP9zU31c3CA
oj5yMgDc6YTqzVW5cj9lQbxhTV9pjJoOhplHaZ0l7JW+HcGX8uZFUgEB8TYKl5LW
qV59YW2g0WF5YFLT6Erevqv+ugmrSkfDEoaekK+45ji6BosLJrL3lfwtlsJhEJtH
lND1qAcS4+qs11ID5hy+XLDvWTqXZKerbbyk0RDW5RK35ItJkAo8vacDtVspBqEZ
1xT2XNqSO+YvPD+YjwO1rUleCBlbCa+2kd24f/4y4DCVKRGk/Jb57ZqtTwa5s/mn
9Z6o2JE1KP/ctrZe7diyo9XTvKslBhB/iIWcxHsA26Jt++ByST0yIs+UG60+4+kw
cBAmYfdnkWu6QEvV/kOx4zVxNWoqzdBRS8l4uYJJzXeZ9UI44G7eGAorX7pyDsCv
6EaV2OU2/aWpLNYE1eC6bTCTDo5JS87f9614EFzLR6GUl092K9csS3Z0Ymd1q4T2
RGnCoyWVuTW3C9tUSI7DqzyRQE6sFojFW8Rt9y15SZ4qD4ar/Oh8C8+/KM3GfnIJ
w582nNJPdncTcR9Va8WLdpFcEcOZorESCtBOZnxIc8FSAClfDwuUtkZ32dCv0jSn
W8OCXZ/TOBl0DJIL8VNL0ZsrjWgxBSXStKxqG0NRrg4UaM0ZRCTv8K1AUlvU3j1r
dEiw/LGBrifKwbg8uko4NZpp57E1jqJWp75QevYPwhxVbHYBWSzZQv9Uc0ksRhsX
C6vXY45C99NULZ4VQ65BAf5bxH/eYa/Qb5oOohqGtvpN9hLDCziIODW2qetql9Eb
5dSQ9Y9HZAIspRsNxj4QoflJBvXnQ2sTty9x3BRqc8+jEEc4bUH3vK1GqAmGdiFn
LW/jTQOSLpE3WFPGdhLHmeFD9ZZ3AqOrTIAjuVaAkEWjX8rNyv23DmDgsJNj2O2o
utX8a7f7NymYRyTMwJvImzFZTJypLoghuZNpaRdgPT1Gh1xm2CdzPzLytxbqmVd7
hI/TDArP1J+RaFB1hW8gO/5cbHyFLTQUkevkVv3X0S+kUDx6pXKeXtyku3BEE3Fp
AUCQ0z80KuCkpTLmJBKMlIK+qdWO14XNFHsWY69yKPlGD5GcKUYWGRftOzk+IlU2
UdxpkoFt0EsRdfdMkBUC2zzdnEuK7AqfzajYV7MBSLg6EwMmky68ifRarhVkkPV9
qn7P96tj5A58OD1TSI0R0JNuiw8Ajcq3oCTZbtSSS8YwFygttqxyf/+kSe/EEo0q
pMFliYsGeS0A7zFJ2c9f+I5mMogbFdug9smXXeach0nfzTX2noHgE8LhVPw+kNBC
AUG4K1XDV0GXjlwZALeSJEaCW5ilirTgT1c+1gUxCw3+Q227FXVoBGtvDQouXrvY
ozark0cZtQ1Rg1VA0+nZ1i/DkqM8txCPp6rcdj4EyHOzNLfPwmranNkZlDMXXJWM
OKmsGJFw0S+kNVaNOOocqIDfVSP5ErlGWAoX62QI/g9R5iUoQnT/L0srkbjUkxz2
7T+jYk5+r8EljEOkD2LRP0bfuewLD7/8qC8X7OYuPXpQ7gAGO9cojb6SbugWEnCi
Hg1gAO3fqYFvD33TAsI2AxpZYNkvdKs0V3P05eGxBEDYTPP0uZNFybd44dm19vad
agcsrU9lkKxYrkAE3i6rFUBxZ1yXfmUe56pZNjNOn/9kgmOWDQghU3QGs4HB2OUD
ccTtHuiWZ9GxmGWrEJVPv0HhmB/Gyo5MIebEYdZb9z5EMNSy3fa3754y3EV41J8f
5+MVLmNGa4k7166P2DrSGrvcOoul573KGPEGQP1cEgYpIZgoo0pG4xIH8NXcj4lr
rFKzvLX76pBjLS+fNKUWu3lSlc49owPReBXtLFwSxuzK43NtphQ2jIMIyYuY5hme
mev8IkuAOdAQ0mB/pWIR8/RadFDBaDzoG6xPyEl0CdnUW77KY9VIjpqEA2Q76gX0
wJlJfST1YY31U9lrw6fwk76o1NIBNHhchEiWV7dLIyLq+FsZhblY69GI3DKTvCMK
XbXdltLmp3M32xh47lLtQXI0rSsO96S8gEwgHEHz92qtTFoNVa3yHFJg+Pt7qGzg
SXoceSDnKLk+A0RvaXPr9U4E0VaX0CLo0I28ou02AaA94R0cWjfvwp5j+T/4JuK5
P+HWC7MlkWzzzeHCTGK5MhkUHg9xpEWKbR7MU+dz4KObb1nurf9pt8KZ5ghcXBl+
r4FUl4YIQHwdunxMYXt1/C8q+aU8e59bqa63nA+7Bhm1V5WRvoZcxoWwNfNydJzv
KhRtI7xOxm3a6+DY7cXiBtyN9bg63MwADcF5IvWfiGti6Pfot9QiXKPtBLD1shPF
7wtFoRDbZagXrDC0MM7UiPOq0oQ9LslC3fpK1BFQ9+Nwhouk9usjgZt9T0bDy6gW
7ZPs8Ufg1xLgDtw7rMmHZxiTIwxMvulwuafcOuEH62pDwEXW3sHcc0/ywdUDGiL+
4t4V+sgHaAEHRKpV5ozRSEcMALjE7RUC32547rccXi3JrYRqGABEizd/8Z3aSMdT
Vkwh3yeQI9TzQAJZl7gjqv0KSc6Mk9hFvA7s8cHPflPPkE9PnGC+xT9HKvvG7pdD
OL+O/ihs5bLQjy4QI8+ddWRK5VY8apBuQbNcbwFD9ETsB52z3eI3MLzZIgldVFLK
umcZxMnrGIBDOpU1oPTjv8AxVixq/WfDDubhqIgUuX1HB8qFjGSar4AJZ3tX0iGq
Wd/kPWz6CQle5Rb7TxGHvZ4MBghqL3ciMEfqeTWLJ2bFYufo4Rqo9qX8LlAWZGCN
5A8HgyqiJMwVeFyO2YqvfOSHrEmcNknnsFfE3VNnvkGEre3LsB7cYRH5lIH2G5Y2
6JNe9djI9j/FcBj4PszXV3RLf2QzkBybms8QQhOMsA8RN4LT2mo4Ksx0z6SwiHQn
LFz1jSgxMvQj0ShynlKyuvNI0/pJFu9UYRG5aiW+hi0ornDug4DKIQ1yNNC3VbLd
iT430XShPr3cyZtOne4KrVWemqKE4sgFFj3BFbpg3qc1jOLxpUpLd4enVaNTtssz
EDfolEpv9oSAkTdCs4Fq//Z4zy6bNOoMO+WSU6jcu03/l3ARLiWxbDoSvz07a0/N
P6Owj1CiAJvRrQh+cOjImB2YygtRSgHfZZpZk0LluYoag3CWakC/Zg9ENuA1FUib
aZ6lwZaZ/PV149fVAkCT4WOO1Oc/H3kq2lw1qJeM/OJix5iMqXuU4DzYaMbiGbsk
5ueQxMiGEavmc8Vg8z8hcw75ESK9keG5a7+FkWs/wt/aQT3hqNfNj5L3/7P6SvLF
jzWwtTs+dUd/xQBgmS0P/5U161dGLejRv/HtMq22lGLWBrKXzMBZH2SqCAKHDukq
PleWZ6qDOE8UEY82Bcy3GplwZBD/kE5pJsgNMeLG3JheuCfDSaIrG9XuMNytCdkt
JzggRe7eBEoaJBc8eL3ZfcA3HMod/eMOGlWRoA+WfB+rnpkDJ6G06pteB2fi525l
bPGKvMz+jTL+I8v6IqbZqJFOZWAybf8N+/68CXh0flntvDdWN4j/QhPig38wu8v6
GlHnwsX1lDh/QHyh/9JzhBUGx+mSnMYqXLf6BmaoWbZfwidYAebaBsxkV/n65GN3
gxogCN1q5/vrztVGLaMBOp8ijKLl3LVtNrUUyxGE3pGsnL1sEfGWWk8yBm2sc/cy
xygD0jWnJ2pjKQifOFwDUEUCH8GFM1vmLsSV78fgAbrtS45i+n6YdmJ8fLKkz+Xn
tCajGprvGl69rClhKGCi+s1NYgVItaLfI7vAP03g9jzvGmOMmP+TJb1WQv6KlCk+
OSN7jGVxegwPLcGQxqkVJuNKFXVSsNpxPmUAobyT9mieUDE+cXirXIQyR/jGFjDc
bhyISaLMvzKCAzM0+Xqyhib5Obwp/Yh6h41JUn4y31YTU/njXjUUru/plLNdgOM/
pfpx46R4Cljvf3RJ+LK3cFMVC1Nd2rNHKev0xCbopAvsZJOP9EmdqmtIURFCqjRN
e3oGW/BcjDJJDeUzJIZT7s6SbnKceSxXwv/v694WnxcRxWCR3p314g+Y92hYMa4v
VTXEzEAu8ISjBL0Hpuilof+0uIpDlWReaT0IW3I3ZGYrUh52j7e7MqWdju2r/01g
UEDlNzmMVKlxTLGyqV/ZWoW7P63hY6lndCilNYoNvAvZG2/nZAbzID91wnM8TgWK
amBzRzmgasUcQrvAUfzlyV4XfWraJRcnG7tjl7M4ei72hrfXV4uW3mgayiqFWHvy
66/QElGa9KlnJ9RbX9nLICtosRSPZm5jQDo3NjOelnwADqnnaStafemSXVC3TUUe
uDEjk/2g3Jo22AYm5ZkVncj/e5nH4jlopa4vKPb+KEX/RLXz1PqEmkeiFPfOSrrw
chHXZA8wanX89jJaBwsm4I1E+mDB0Wd+CjfID0uepNj/myamjocXmGWizhpedoix
i052Pq+js4KKlA6Q/KoqZZ/PybRz9XMYgol7HO1WhMmFhg1lbNDgU+K5JNwsgxBM
WCqLSboBCGYcYjvCjNSlhJt18xN2/3Msvu9omO9xg3Rp1GUXuipX/2U9zSmq1HAn
9Pr54nnrr3nbcOaGAXuyndz8OtFbXHapomVh61WOXYqbjgBFXmW1huD+t1tcpYp1
0wsXuP6uuLDxsttULxG6AJsTXDABR/ivv3qprS2fvRys/fNejJTThjz3ezLKWbdO
vX74PPjRaAAeTq74OcBPfXuxYWA/mjlP2FCpD/Ii2pcnHetlupnqNGplit2rhqOP
s/pZtzPUBzPDCGeLmeYBNXAP2/MRoJCZTtLQ0To9nzfGjLW0TBdBMz2c8Bv8RgtL
FpLUb186kvHca9FuqO36XFYYDALgwFB9rQ0ytNCbayPkpE89av6uOHETsbUu+bUb
QjxiFkAmOvS+aE7Mx1kibGRwDYv3tpGsQxgI3KoH093rr/GhT487oOCEy8nNuJmY
rWTy41EYdh5AFvvpyjbyimdv5i4XTvEup23Dq9TUDyeTWXMY4cbc20g+mLY8E7Y9
jZuRT8xWPsIwzKMqNOUCCNRA6vkIfmWyL61xMtny4Kr2iSk0PAf9QmBm1QRV33L4
W2d7hXCAWllQQJQFBppI3AF1GLv5rAztC7hvVW6LhDWZgbcBrxwswopcDu1ZJtb3
OxOitQfYGCI+W+uT3NORaUCzlqlpIJ6vYohtijZGnN1enqU94ENY+7HgtoSnp4GM
ykZTyfILlxAv4T2i/bpYARgbsg+ep96MaFiPu2wibiABxf9znmhtxJ1+juSGcxnN
nEvOzAAZBJPUDy2FSwTCb1EbvNSHEXKo2HHlShO52dCWBdt3ty/BQG2mXYy8FC76
clU6SOIR6E/FcVAWeXHk9gWmHzbKYW4Qjkmxzfo1Vn/Dx1khuhdcxUOeE5gwEpBd
TTUG12+DUuAJeON+DkwVVwVW336A7B7RZwks3simyMLVpwQUkuCqjw8VnU+vSW6v
PkFKh97tRmFImK7QruWf0zVhhZcEnA44e7bwAYw38vRFJh7GhG5oqgyZ5K4LUSrd
q1haTLmG2hO0/zwCAMEg8e8lcY/ilQWpLBM6jC4/vi7KBdY8HwRoV60Y9FuLuIQf
PVBL2glciQSgitqfwX9mk+DiQjY6m8b0WWO7EbLy7S7kYfyEgMmlFl6XChoSo7TM
N64Mrc98n+4bhoL87mwf4GriWDXHQ5PTx3CRetpUu4UgnLJ+sUF0PRb8NJHk/BXh
4cyDnCdfp5GR/RsZeqydZRi/XS7aFyTa3H5NjP+lH9i+EbuhFyqJJk7SUBkl6yqH
8vPDoNjq7+gPHHJa3Cwi3yzmAWtViuY1L1a8tgA42Yx7ti9mIpdk2pg7t5/ZrJgm
85aODpYqeUTseEhupwlTRQnjS6LdmkatFlufUSsdKyn2DSNgIAtU1DHoQen70k/n
RZtYKTljy7s13kVN14e19m+3evtVydblIVK79CicOFsRBBzdS5y+sa2FVJTETDur
7ywLtSGdQbSBLRbXD79pgMx6gJnOrdaACGMYVrUNtF/AhLixJrX8KsIt62TFoVQU
Iav0/BdSmgGGF3eRabC2zU568FVoeMQFp3PPsY8gW3VW74C+Llx8BjzP3ZQhNRTS
4Klddk620IA70a+bU8h6NEmLnBZ5dg/MgrkLpd4hnNA5MQ5z4voPSh4paexHZqzr
HuklwY0SK7jJbZyRFLFXrVFlYXUcPAPRJrLoxBahVFn5thsJ988S/aztDKVy9Sse
0+Uh0m65ghvmU88A1erLt7yRsY8xHjz5qsRJzX4S7GY54J25kCvF+mjzjFChxWCW
3uYpBPU9LLkLnPGwKW04w2iciXxw8+IRU39gCcBir2p7stEJAfuFD82Fj/roKeBn
PsvOMVFoYV+5fXaNAlZI/7biRF1+t74oXupIt/3kp4dJlp5Mxs+DWABxH0hvfuTN
nsa8TeWo7mbCIXICCdCVW0cA6utvUKRiEy4DGbkoz/zMLVQRJrOIelX8oMRuajLj
bf2sN/zvm08YiXWnIUXV/s2WcJ4LfrNbFAfEO+oRZypG1WmuxHX1Sx6t3gXwzLJ4
WDlM81e05Mijl0acPVG3LL0aqM4OpD1HvBO8qdws6J1H5Xuylu4rGhO5EPZWFgWd
Odr3xyvAAn5nyS2FlhZJG3CY9tQ/P7NPR7BUP76K/HTrju1KUoUDIzzYi+vbg1Y4
5LD8XhGj+1GDA+7002EJmOgopoYy+EgONB4KcWRLiwUq5mSb0f5orXXiJkCCYN6C
3Uj8Ecb0pD72FvzmiagCUnKkTD4xvgZEyP1MsEt56ph1MgY9ClFkYL8CCyZP9lIq
HWDhvwisid8ax9ILUrgSdIgCFUEX3EUDhcOhrE875Z31UIJRm/m0L9f3HUZdzyQs
IOkOdACNYzJ9SYyszTpwmWW7VFuVYDFygAy0Ur1TyeJxrib6rZNloI5Fu0Dvbymi
iqO6fO5zeeSr48K62CN3kjBvLJSIGtR3hMTGeStJQsSIvrLgbbMKiVjLbwwBcW73
rl7+jK+haqblpOB2LzoTJ3kH/m63sKMWiUjTGyrHlkz1XRRDop2f3hGp29sN8NyO
Q2BHL8d9CfmhgJ/zF2pwXoj+yjHzS22E3TXObD19aYpfnqywFPSrB5OzP2lbOQVi
/r/ewpuGoYznU9Kk9j9Q8GphSMNm2ta6LuzdWsyKQhQeLZMNGO1uZrvBWLy8vKFl
F/X60kC4kiggHUaPgzu9flDOOL1raFLuZoMj3AVnnNvHWqDzfpWirg3wk2diBGLU
xiU45e2sRMO+81E1zrYgdazG2BpHCK8HZcfL+TFQGo8y7nIXgErWzw3+a+L24ZNO
zP6rr3/L8gNEn2xP5MnBlNq0VvWbjNrkWyAvq160ip0mjWCvH4dIAWUWPoXbBUU7
HXIsKMyJyYcC6rH6AC0Tg8JctN8yyuXwUd1xJQ24+E+eGbySHv/pUuqhAytM/1VS
4zGfCxBLal5ik6wZ8UX3qeGiHsO+xDbJOc7HM3BTwmu68mUvL9XOsKTFIuW2Hvnk
FvptpgBRS7JvpfzHYoVw7fnIZynwcMwhECa9AMLK+5i/Mosc8L1k88PPySzIp78w
XUhcddnKNiBoxVkr/FNzCCAD6gXbmi9gOWKUAs2/4FaSrYVI7g9snp5QGD8HGDP3
7IVlryEKD4aEGMU2/ATvtMJwkjiirmhhlphju8mUEci5C1IZGq3RHR/MIb+7dCPd
+SCHpVbji6QUsKoOoUpFIQ6pAyNM7Dkdlpe3lgzwsZ9CUvn158f/QKlobhSXj0Ub
5tsPURIXxJ0+IWgif8sLMvqm54XiKLjAbD1siXzArQFQk3AUTlIIOca6CTVLPcw7
S3vptuE6/qQFu5yS4xVzXeMQ1SWvPHi0WOvRjwqP2TsJhCuk5aWSi/DZYCdxB3xT
M/YUf4HzRtKvuOtMxD4gIg2lmBbP20rAT8PkercMNam7yLwGQde8Wa1yLzwTSelp
g8U4pfHdTqiHxgpg8osB8R2PEndDSFc26ifCoQE0ueycgmMrlwVvfqxOgLrh4zl5
sU8EQ7emS+eTWjZ9980b5iXIi32voJyhBJY6XKhW3d3qH02+GG9cnk7LHR3uL7EK
DmvYZMELAgUM9sLOex/e8oEDDErFivRjUgeOav4J5PWgYX7iOxRka0rCAn41R76z
Lq243+UidJI69ZJAeLbAFpV4tYFOCBLvSHFuNirxUSguLGAaRD2d/8/9AIRz5wZe
mju43DxSF9wtBwKHgznyEb261fulwMSQbOtU52W4eFkrkV13tgTGOm0bEiSTCBTe
//K+IgypFAAO8IXMqRZcGmiv4z12qpjY+sb5Knfh25y0p+d3OnNDkR+0wFFavbPV
1HS4AGGtLIDsFv59AJRXmvfEzbjdTNaI3uWVPLJjNoouLMKm+2SaBB+V+sQAxUqS
PVMoBcazwku8EtkWkezkSNE9/HbXYfM53UHnO7HI6BycB+3AY2NQaldIUb4ZSXIv
HPxr948LEMV9OtJxHne4KVhG8ve66F8c+CFeED+VYSoptPHTv68Nyeg2JLPVKTDs
cxtD0KriMEsHmGcGnO6fTSbRrgz/1Py/nVARjBS/1do7INgRyJUj4hhYpRAkn2kh
ezakOf1sd5rbZBILxxphCIrKj/WWfZ4TtB+DKS2f/vN7bz8EVXj/OHrh5RCwDvMJ
+otBpMgAv4wZ17hEAnyXvR/o+3XnI5GA0fOZ4Gud8I96blXzY4duQSmPQjRK2Rr8
gSzpYhQ9PyjkBOWq8ZqOj0a7xUEaJ6o7LCv6DD+bu7qtpPOmI2WeJu037fk7xA5T
Njvm2NZBXEF/mwmr33+ThHTvbjRcUNSyRvlVt8UOcYeffEhUpUZ5Zee+6bKsBIiO
TDU4qAFFcKL/mHciwyBVaIUcXArekBjAL0hld+Gfpcm1lH2P3HdLIK3854LoNh0K
25gOdtqHRsynxwdjdN6JA/11UCy+TiKeWtUjyR7WcfVZGbQETQpB/YHxubkPuQru
W92WLY8Dchs9Ybkgm20jP3UdNy6nrCAjxiqDtP8h2KSmFrJJHa87GMrO/IjL1Ssl
0+2rbG5xFIT5OV/V6v4sNqNMxCiBolDFm8Ior3x6v0ANxdWqpNRzJWJOjDpHrUSS
v2XU0BJ/Yvcgu9Fu3bFWNCKI/uJ/L1EU7/eLZ+Sm5W9DTWRdZteMPyViFuK+opM+
bt8WWTcdUw06pE/2PYLwJvDnyQrM7XS53GhSeJTJ8Y7uwx1AdIn11i+XrmQHK50X
OaI9UeJR+6afmF4w0s7Y6o8d4v7hVcYybNr3MUbiul6kzHVs8xRbF2oSc+23KjV+
jhOb1ODPXDg0qJdHxL9QdhVtuRdCjx0uLLG9tpx1yxonvqJMCirkNpOFETYTvkz2
sNxZl3JD55FzSrQyt/bSsM4gFMxrUhNGkQRSlv7a83JW9nSjqEyZwVCRHiFA3kVa
BlGxB3uquDeSqLyo2ZXZ+0j93u0ICs/OdFZ8WS+riFSpcV/q9hmZ/UgMxjyl+L52
R9A3wjjIt8BAeuzGARNglSetuTtJ+fRBEX490nrBJA6OACS0rrE39/j8wOT5IYfN
3ESCGfd/Y7jLzCGkUs7+jguSrqrv0LZ97g4Yvprg0mwIkYeqDFW3Gk+Bq32HRXGj
kFWiHBMzCKXC94hEeWIO3GcboOUefKwMHlB1clOAiYNVULWD2L7TIuVtIAb1jaUz
JGuT1toy3cwbCjvf4Tago52waBWelCfk7npFfdc19C7wjT3sdwIhk8wBwwCyLQV0
jco0k6VoTYeYYKyXALsZhQ3bX7iIfWy1ysfxmFvTRR2caQFGsOH3UjjZsks2LVZ3
uMYYGpLZdsocomaLpUJu2t1CkS5fiZ8t4Q7yWkXwReEKkHxtvT1rjl9GnnbPYkPf
pYR50rwTbjecczp2ks9OP2rqJWSsicGh3IVXRRkt/ffg0X2F/gQ5JLT7ohreG1uq
y8uQQe7eZft15pLesUubDhk1/RFpRvkvWqMUN6HFIYodxepgVz1lijvJbnKUVESO
2zkACV3asmUQF7tlVCouzKf00rKyfm1hoySmkAHKxURNOtjHKTAX4Za4xrHaUqhF
afCzbNzEcq2K0jERJyc2WiaDr+J2tH+4FyOK2y9CxoJihzOeYrxcFcJMjFknBCIZ
mbc28s8DCUC+2QB01VZJxAiGNbPOn5gpaUdVbMIRQKnGK4swzn8sobXbXC+7sQwy
ECMDkdFI47OaaLgyda8C0W4l0ibknjaPqyN4RjBzwnoshql4sKmGOkC2dva3Di1T
QarkWZLsI7nRtUP9bzoi1jzDFxkhLYp8r6zW4ZmtCyaITrtWoXjFpkumZ6uto2Gq
fYnpzYQYk72CZSgv0tUH1/oRRw7+Pop41m01yb0FDRfaOLgj6DE7mRBUzl7QBU9u
8D2N1OAaq9+kNPCLcElMM/c2LYdx0C1qP5RQjSd/xiLelZQiOh8fTpvuMVfjZqJs
RFyOHox+NOsBw6LhLXv5LH9bbH5fug6EcJkYoKt6OB2XeiRuG1vTumuHENeo6Awx
i9h3lzSqPNXiHc6LPxWbzf8C1yQGJmbdWl/M99eOUshj/wB4klvO2tYFvOg5DrF4
AQuYUgSKGaqHeuhgjFXvnEejh+nX1lEf7mV6Ro47QxQvVRAuR/LBJIWVc/tpfs4G
LXmeSrDc6BYop5r1cJxBjJQ5BWV2E/ndZv4WKRNde0Mz90XPu2vWTX8bjTOMg6Sz
Y5bFO6Sj84K9GjK0N7gmihnyeyvmigCJSUmGVD/50/9lJoBUAroAQG8jiH3JrHSh
Xt6WzeEx+9AJuJjGrazgGFKrl6+F7HAsiRqk9YAUFf8IuU96SI4oZw9sgB3V136q
UT6S2qqU7b4FiuCQHCTGbKyIfGch/rxI3MLgq2VV4c4CYYPA2U5foRDrIu2B0PId
qiDYvlJ9GqBPSF+tUYflA/NejJ/wxi7OKpnPD9eK1KYzJgf94CS+cQ69o5Zit7P9
AL/NyIQaOjm7RyWy9SuxuIyYz/kMqvFgrpopuUyhkGQcuKXlSelD2ioJ1P3Rw49L
DlQh18LN8Oro6mjs0wqadE3agJzyNtrTNLhCuV+XZHl8Eg2OxtJH2pp1GgXJRohA
hBpDt7wb7OK1VZnrEMwgHY2OHi5aEWKTD/vRKd5gvOX5/6i9mQbBRC8/nZWz1SSw
vpj/ygrsrohCGERk8LBlKI1Wcr2yZ2Uf8gL6xGippjrh+gJJW8oa6SsHv+KYs/LR
rk9VRrX7HY2L6gXZJwZBtTY0QyxHVg+5VwFqBdvTpLYjLi0ndCKqjKmezegCbV3z
AedkyUlR39s/9qR9LiKh0Uq5tLZk9U9nXy8JsZjq5Cn6dzRLfvIs1Ap+a9P+n128
Jq1GZfPsR3qZEwRLBpWkoE9mS/7ttiGhl8xRkjmot7FT+jnmRQpcDk8Hqu2iccb1
9GBciJKQPp8MYnZ+J1lsbfZxmKFZ6IMOEHbSldROhX0eHYLT2FFqQhis8b0jXRDB
h5HoyAyELHuUCrpPYhKyTkcK183LI6EsN4jx2xnb2/fAnJYtR61QYcQ8TRJfNDCx
LE5rtaLNuoWixUtZ4SaK+u/H0hW+SxTRCgczlFj5L9qe6Y/vh8V3r4o0VYM/9WZj
c99QfwsL8FaciyRL5SOY6ikdiSGYymkOtf2dra+ZLQpn1IajWklaQZODvIIFAalG
fcvEsNEDrTBbpFqc2Lox1h8XY0KaFUy/4yx1jjfA1+aYBSY4FF962N1/5ORdOPC9
WWa4CLt3bSHWO9FaAIkHXXznf6ijzz9NkXV9asfZUs4nzloE08p5H/huZA3UWDuX
u/JrlY83/tH3z7agwGoRGnxWWwhZt9NbdzoRG6PvKdiLd2aocre1TQsEhsnsInYA
NVyhRTMGbqtw9MTyNww/YCpwfSkHRPtvOzXjX3baWzafTrLMEtkt/XJncN2YbqTe
BHRR1BCLy2Tw0kASotId14ugbJ9XuF5Ptyp0xAG2eJesW7/S7F83FDfCPPdn/eQT
SFyITDZSjuKF1cJDISJwmIkEPuhjBP18C9zRylj8Ld5Pm/lK0/f6VlpnrxZ2+yRJ
pockR8Fy6KPb+xaW4R2BQQg7pfgzEYViCS2ZLaVGCfT8SragD+1ij/JKZoln/fBE
Z4uXLh3/bKnIErCBcTk+vnAjHZsRy+TIaLW/P4AWdp+bmr/D61K1AEvynE1+KGbL
T0Hmy0uTuYmvqsPW34yjcvNcMxWXPnF427zq4l/WhOy9eSW1Mkh3jlWyZbzGyCKO
tBTJ+OX9dEB8LNk8BkplwHL18pcfoIGwNgJxX/qkpEsOLPsprP+y3pTCcLCQ3lXi
6cH4LVlhYhESpmWLbigZeRSRSJoGiRtM2uXoeWKpv1JDix1ln7B7Nr53kxWXIUbG
H/W2YTQmCk8G+dbXLP/vhE+ayG2l04eA524N4ZV3NtzBoJkDtSOcyVLxiFCnBOjC
YUvfm+xYq+uC9mUUXuAB3cMcjKd1v5X2r8zGjBiCjtDpu4nSt3HIgspGf72eYJot
G/zKhYOV2QQ9V3TjoFiKlbWFJQKXUeddeSLyCK/wGFfNus8I6xjdp1C26NAbu1lO
Iqm7YgSXtZO0vL6nPKwLO9GHPFsBWOnR3aRuqNNbZ8Eq4A72mW2WQPOm/lhG2Sxz
ssGYjM1h9UEfenG+JW0unBakVpkIn7THV0jDSYCTM6giMwHrH5wuyvpDzdDdY3FI
VMjhpKSIrM3dIwV3h07aiGQK2DhnRaxCF21sTCJMWCh8ZFZjmj6Jlcc4078eSAnF
OW3Mbln90Yk75G7vGC16Gf+WwpuOpjq0bYzmsuD34L43IuNuwkIHkbcWbzW7n4f3
V7WtZ6kW0vzLOUF72w0nbp98nIx1x/4CBV1BWXzo4Grtkxs8bfyKEs7R2wtcoevw
Azj/F/Nd2VLFnykue/YedQwVmuM5DGWRDknAs5sxZGphjnKyA1OP5DWoiDhkB+OY
R7W5IOysxLy1W6dUFsxPbQSWXACheL1Vrdg/cL6F+m+GZiBCTHDGoglXKz0rqHH8
qHF2th/zyJ8uHI3JXqtv5GsTlLQj5zAOLuf6qwp+pNbJioalsqn1AwjPUIUf2GH4
Q+/yuYXeihzCyYHW3iwmwcjjV0s7v9rK0L2qVY4/xnfUM+WXzymIn641tzKy6pVH
gcuSmBmqkY1R2cHgK8e3nmAy0xCELIJ45o3oNFlulZkngSerJiFHrCXIlwB+mzcd
ycv/cUSVKNckcPWkZBN6VHxmyzlJj0WRko0Df9TMmQ/6X1mTextk0v9+MrzQkWa7
wFsVAmtV5o08NaI2B3IvlHd5pAKQfg/EnPvkYsh38CG+Et7NDEFQr6p7pNoU+MQe
hC0LT+9BUbka29NZOak26LiDsHL7JADM28JKuFOsjZQ8e2/PuJ9dDdjkteQ0hGT5
AWliStsVgCd3uJPyZTymaXivXov9sZmxICqaA+J1uN3M+wfu0yVXB1bEvJxtgpZh
MK2NLFxKNkKvYgChtT+bCOfnPZIrn56Pz9i81jCeOstx2sHKHt5VdwIJ5tYJ2TTY
kYisguH9rkQiy4SmffMKQPobSnmoDQMzLy2hmGtYA6IA8/SC8c6+XjCaIsSEAfxz
SSh+AI5L3hxUH3WNYsznXE2Yt0xGaG8oEi9pjL+CB4Jrw1FCoyzwYwkxLWWzu4HJ
pnCdGLxFhgwByVdSdZJlKhlMlf3l1ywLdnML6CuOWeHUIYgeMxDg24W+YJ6HxyQD
4/UOVchVixxxYs7vhIX01WFADbbLBcX8rU1MpeOaeTe96n5XRjFDKpRpiudP+7rn
mdlGNSX4b8Zqi8EpyK+/CW+Z6sWl/oM9kblE7HY9ykl/Tml3W08u3fZ9xJXQ6+CS
iVv4jmIAW+38G0q+pyOf3268dFgoAIiY70GSfvNFLkugJOlFhEJrCJ8CNvYcTiYG
IB+yr+03XocVoXqKHUhK52lM+4PTu+C0t37xBcJWgQYNRC9qpDn3kn9+Knb/jt14
xngREcWTG0w/qgosN5jstkgfWYx5GXB1iGm3O5k2X21j/xQ2N5vX5r0UDPXXxENC
kGMyOLdUkpOaxqWlNGVZsA+6yzjrd56y5/rV/+Rz07c/KPHdbDIVyoYWneeALYu0
VihCqY7nn4LtfNUojMDDQBaazZE1OKjC3nznOUwOBL92EXDhkjgQ66xogTw1HKLW
YHZDkLlsGNnxzNn0BzG+Op/Roh3qazHcoyULOJDFbZR2F6sznBQ78ZnRdvUeBq8X
iBvekLNfIP20f7c+lzKBEEkn76iCVEhYEMthJdaEswMAbu1lUPEXeRZs5KS/Y8LK
yG/snK2o38lCPo9L/lYcOJ+rqENME729av/B8xTeNXdMHahAV7P9zHOCDpUOmpT7
UQuk5fD5vU/P7wC1M44J+aisPExxIA3YIYfL/t3TFGRSmmKoPIoV8TWpB8SJn6tQ
/VBMWq2gkBAJBwzJdMNZASS7RebZzXjaZWQ0wXKFpygEiCVCXUiBJIUWxQ6kgTIH
Q3zXZ//7my5+O7cn2U52GDN0lefC+UR1mwkKkaxIq9Df1ZXs6+tg9m5cSiaOEXuV
4z5cAD/XNu2FmsvQJw4ct8SY4mCPKGT8vAT82DeE5iIN7u34DagFlrgetHEE5uHT
VA8aCOmqIJv0wqJACtNiO4H2BpXITtDzdAzHcq02nKClBM8WmAK8qIdEHbILr8uq
Fgx7z4Bb5eQtfKV8i9BUuwxzdsn4y028C7beoOR2fHKMrgzQ31C1OvVQeFKn4ilm
3DcIIs1enpanH/Ne3GQ64/2SoQh6hGPa7jZCuk9eyR8lcprVxxrj6vJQPEZv8/LV
qAUMbssudGue8B5oSTLcUCColPwyaGGkcBAwYIr2lELs/fW/hvR6nPJCiXm2/qg1
sfIHPE0aAYkwO9c/tJkwct6e5EdUGsmjIlCYCxvSskPuxd5rtC3s4YOiFGEbn0pH
UOn/h9GFnCDpR9vn87Kwjbych7HWBhnEskn2wGm6ubbXKsBRWhYPSU2R4S2q6M8W
B3d/hDYi/66Ha6E+duF+OF/amSJp2WRdEU9HDuBRN6LP8WVfUtmHv+69fbPwdE8J
ummKfjeGPuN3CFQ0a5/BRtk4nAiadQv6yRB+CpyiSMwcSDL788ii1sUz8IoAa1gR
AxH7a3oM68OHOvDAVpF7WQhvynu11JFFX6lxAeasmI5NQVPqFAouYQWQk++uMUCe
qc19N/jBwKgNWXrfEHEMRhMKA9h1ySuknmT8CXzJXrY0AfjWe7J8woqd2+8lFM8t
hsr3HNKXHRmaH1hjnfsloWOkR3WaVYvUAuoeaiX1kfJD8om6Coqd5W8smgzvMqPr
4trxv/xRE803hFS5JRsh4tw+duKfc2y7bZW2QN7u8nOuEBE758tGBnT7LVlZD7y7
xce8m5Jz9yjSgowSFGo9yhKDDdMN1/siEUHRE2bVzWHoyYqYsYBoT+dON/ygTY0X
iEijYPb0cJfeyDfRmPz9buU5HjuF46qnyJHUQHCBjf47z9sg+H1zN/fIko9pcBWB
peNGF4Kdltg+zqexTjzu/hEU+y6VytsAMO5B/XCCrhOTJRJR1SgXkRCABrbJ6Ukf
6V1Ji8hA+oi3IfoXOiM1wgpF/OlETPrfmFl4tM01v5ZXzD5WB92yVfJ2T+WuueYI
h2P3qNRNNY8reKiW19ewv8vB6LVyM2mcqHstFlEgVQWYL6PQycuKfmu526PRYjrh
1zCwgWM8Micko7uww7mTDD/rdMVLIzmGOa69MIo4PaeufONUPr8okMsabg/EtP3F
DNSmJEDZqxOblVG5hvaL7jU7N2KGbaacLrIgcaUNzvqLwfq3daEh60IDIR1duh/z
Cz6+1iIi8lwkj5IfnZal+zEOEyuSXW90SmmhIHAGx9GZfrJo4Sa9cvYVOV2YizsU
AJBoaT953s3aQBHBGf76RDSZA0Xaew8hH+fSoTUCDrk6V9wxBRiMHOIQeLUFE1te
XpCYeYKLSVrYKXTJsj3gnptxZgm34R92AZXkavX7bCY8g2kI7PFSjqIaMeAxFoeU
1JXuO+y+2mqyzsMtwmkNNQCqsTa/qSpzxLZ3X7nMBmf3PMf1/plHW+jWh7Upf9pv
DeTJb38syosy48IEeGTHVztAzMhKp16vxSD2QvnMlfmX7Wl/8DtDV3Dc/iBKRUoj
/2UpWwZdPBc1ibJtjAQiJUDlPWiUnAoDbcMaELrb6stqbZBPEnlX/OGZ25lYG/Mq
L+bwEm0TvNp44cP3HWljzHET6iVgwqt75HoBilYyLtOnJYhw7yEXpzx3XaOv/OcZ
qxjbX4Hy+2IQgaKD8zI9KkdISC3rKokWx3yFiC66LBsMtpuz7O6edhnw14CZBmu5
uWH5vYO0dZzbGHv073haesSGTJiWqNfQlsUqqxg3euN6JmDaxQ79haU/rDzCfh1m
W78oADbexWwPdDy9mpgj9C8pFrmiy+XwVGoqNFoZpiIDl3OpkvBEpw43wL09FD1W
XjhqIhxaIjH55tCeheHtR1TETW8SlN+LIbDky9gP8aJJd2WnuNoq4g9J640gM2Qy
0FnQpsDXt2zCei2iAq3fbUUYesrzt4lmlrTJ2Q7hbqE/bzzH+5EyGJTHLbjGr+Dw
dqDko40q9B43t9uCSN0v61LmeIQKvAlIMDJwWF17KWhv2fxIFqOAP3cBMkoJoySg
fU2ocCPv1FyechzGDIQ1C0LfDhlS9JfC6U7ku/S34tIyJu9nSdB6lnm/ZgZzM0I1
JLe8RX2VDV9Ib7BfZLE+HADBSLz/JwIlPIpAtTevZdVxAdC5HZ4YR9fi3OcZ7uKx
ODBQerFGfVHvPB+5eQWXfx1rfq39AFTytzWcLjDFX+rpOQH1rmiWbnNUgAPCgwYn
mV8ezfO6VY0w2+8SVovSqKXGXLRiTga5icqSHzOv/K9VqrH//wdQYwpeHbdKGCpW
hi9KfMpGOlwQSRislp5oZgO7LSZojmOHmOC/LMpTvidLocVsN/9LFsqg9fmr87FG
Sn77ApJUvEyrMFcFSWoIhqQdSllhEHzNPYP29WU+Yn9tdf+XCOeLqSZZPh6lzqdJ
jfFECUCZI4+M8F6I8QOszcxrmjhl//GYNyNvqlSocpPwfn8atcOoyRfX1GjPULEq
4Dvs7/fi6X0RjVgLVIRdaiSqJQMHVxKsFe2shrpyGkN6IguoLSahfXZXuB971PAC
SI+qoGBzs0MqY8zYryJWN+VlsSeNiJMHAZsb4iAcnBZsZumYINNK9oFqhbb0Q44i
dljw3TatCJu7V2CWpjzJPWGgALYPucg0Crr7dMPW0LEUS1g3v971eSpKpKONbVth
sYCMxE56PbtaMcrt18VGqVn6NyhJp/s3ghALtHBxlycn6t56CZ1584F+hSNHl+Aa
yP+6V+r+G2FAg/WZ/26Zzga7DGV5EGq0wNuTEGjpoCule6MqtRIs5ODnPE4ExHGE
wja21qxI/2DmgsC6aMNfUJe4ooXg97BaLkw3rDdRwhSqeSaxipWnCcIe40YhEPLY
FuZXHD6RMGTdoReVIkVlKCxKmfeUoakvuRBLqZfl21g7+BuOTj3Hbg6WT3AF1z4m
bccf/MWmxBBlucpu0Z5WVMADnA8wR40O6n7AWS47X0XMhigA1Pq52KH8rgvv+Nq4
4MOpMALiDTTP/Gv+4dqXWtv/gvh15zlOe9XJsP2Y25YgQEa0SwfCppMa7YTmjr1Y
dzijkj2dz+MFw/oKPSs7Ss8KXQ5n79TgTHY1A6xej7ECsn4Y7NNQ7xdZZQB8/Lv3
4M8IjBBChgFIHMekYe4pSVfQDnQ1lpA73PPIJ0JxsHVNTwN+aBSkqZ+40SbPFc5u
NEDv5zcVzK05KhjUAaXG0GRwaG9/8TAXoJHOwSzp5f97yfTrmmV6IQV0041sI4uL
EnUsO+dzw007BHKLAUpoC7v5C36Mu/4e2gvpM/0LOftYlcWNMnVFavzMetTGKxiq
foHEL1Fx89/+lnoQV8L7r0BMY7bQFSNkfwHodpr6SLAfcBSGXWGxsC7Gea/xJjgl
PhBsjk2z6MDOkTHwnp2GISSOaJKJ7+Saet+Dd0UWG87ntfFRSt/d93NlwzTH26rg
K7YP5eSY0PL99oBWgXrBy+XhTE3pdWePvzDvZAlvPkpUX/CcRyFiu5znR/X7i3ol
NTMiKO3L5hBCIUtuv7AtvEUDZyT37CwaMtJRohgI4WBHVaMz/V33U82BuxdPizjw
bSoA0UPEgG/DPxGWGTuxXj2zh9SwE6+lNd2dbYcgjRWLMPNc1Z3r+EkN7QLr2UNL
lC0Va5KiBOgby/LOZMQSHSEcA+DvoYOQ0fG+F/l8Q1oXA/a6Ly5JGrPwwssVeCeW
yNPHNJexoiPQwIt/jslIHvA/ey76YjiFk356Bicn55EUJajXWzc8dLElpO/CfUPv
nd0dbv8OHOYb0oE93xO8BE9bX4CrnHO2seajCfLhWFYEr+zZe8LRcm5qwkvYcbUb
f806/0olYoo45CrROtpM/qTrV0tvgQRSBnk8Prq1B+p/1tkwXbBxAlQFIjAVmgFH
9Va1kVqa9DVJC9FQcW4+L9ntx+1C7IiJpV0AMwiXsw+cGjmQGz9gylUqlQ/7c5E2
zllmRwW0ENeT7meCk9ZsBy/4xzbGX4XXCENtexps89t5SFPUF8jbN0arNSKlCZrA
T7hcj6qJPRQy+Ijzmm4lPD93USx82AMDgA3ax8aPayZ2XSMudtdIob8X26evCtEz
GidLUsB6+GeuUZAcgskOJEHvwSrXEjeoJVu+gRioxrBcAmF7uicPAQKJYNExN2SB
DHoCoizQ7Iv+OnIa9NlXaXtK7kfM30YpenZm1WGigtBUsu3Tz+krXSqZ5uwn4ZRM
TIdHun0K0c0EF18VyIhTHL2q0aSDxOJEahTJ3Z28BxwpwdZrp5KXTniDafqp/6uF
fr2c+BAYNc1mW1NdBDdZRkGqVDQXT/A8owb8BKGOxyxuMUZ5xSqATUuK/ODi6Yaf
5jyGLkUnYVBTmLNntOu2h1VM02pSyywT1TBPIt45JL8ZZVpYf0Vq5/sUSZoCWClo
SOfUY9+HC7GWOZBuhUEizVnMWg0McUIPjC0tatj7NTMwtF7dOY9h0oap9Nd7UIYK
gdE6wvb1P++bJY6ssLPkItE0gkU5LpNVv4Lb/QLMvWJeBqplTa4ch4KRz0+NH5IB
QRX8jxQXgB3Frp9GWT756hdG2j9Pz+CNM6INzN953vI3PNmr4egziCoDblt35+XF
6a/V+3AxnRpz4bk9GyLbO1yz9oaj+9OW7G68B2DjV4RIbiKEZ2XKskTnZzp2ABiL
HlSnMzOmmVS5zVC08K0LUKs8TpQ1FIBjBiRMSkjeaOM5MZg39BzN8eYquZuBP23X
fudsyIe/m13gU8jeS+I1KuTk+5Y/q2MOda2DAIk1YuCTig6OjCeFIFmp8mGXySld
TFFbafgmJfocZ8ONZCRMk68ISTA3xu+J0EYv62Y4892dmWWsHmo91NvgEVP0rqP0
7HJbwZ6qeYY/P9IgkjtUH5ocYXU4uqpD8e+CGb4u5/o/ciPpsCnQIPFKdP2QnXKC
NvdsCl0sgem99cWEiWoj5CvKXALKyzfkw4Q01kpJX98AQrs56sXkePyfzbqfzaeK
GckQ9bgsId05xYJT3HxrZ5MGPYIh95x224AUvpkAPSRPG0pzQ1JO6kIJGvQ6E4Fh
OdKMCF81U7+CriKnMX39ITWL8DTEQYFLtG8HKxXTevYL9Fu/jnd/yPkX39QTaLSb
oKVoDdbaKT5rZjsKbu87ERP4ibKwa6Iw8Q20cnkxlLYsKglGRdeHHylPL5cyfMba
hMiWTseDHIfIuhG16Cipu/QSB8APRyjSGo5Jtg6z1ctoRBskTe2sPLmyLzBMTX4L
AwLYZWVnOJbn/kdUvABAbKHQStvlAMM+csGfvm8MUz337XNrCDxX9OVl2D51+FHQ
gF6H2pIZVliDAxSXhCfl7R024POSwDx4YT/f1HoQNH+JAW+a+oqWqrHajd37GRq5
dema8SZ6Mxid+KZZVfvaf5j9/N1TN7WUusm0ql+CkeF6UF9/r1aXFFTvIPtYAcNz
+Xv/Exo62rV3iBwvpKQVcc0hRg2Hqcv6tur/UzekEBXTj2Xm6CoIQZy/iUek0W3q
DjE+UCx34E8vUWO+47UFE7ryDMJLcr+DDXw8ishCkhoTOOE4HVlFqHep6+F+I5H4
PP8bUbRCV4XExB8U8o37HQFo8OeYXRERyKKarg1+BbYrnTjqzNMPjMy1NbX86yyr
pX8MhxFKSf0nTGHs3Lmje7ih32R2+y961330TNz2uSGng6tbbz1jjIGF3XAnQERt
Qr/H1ZInmf+Xz88HaiUj5AK8UTNmINDJ2C11NGHR2anCBoTM//Soquq3JktR7JEW
UU76Epfyryh3UXpZ0iiFLXKWytgG4EFF2nXhv8ZFR6Q8BcrHJ0vkyN6LgCMTcwg3
b2nVrX+tM7LU9mFdYExa/GGDPkQBF7LnV0eGzIvNEaEFc+5bPxu8bFx4PnmFKUca
4LEPARF6akCaR+CdI7h1MRvdWKJKM/2S2/LPgXlXdhpHM01jAj3Eh6vj5DnNHE2c
J2kMT7yH5rad5dhLbtXm+2PTB+W0L+gyQD6QZYnSRlm0gWv+jWogxnohyr2j2iHI
XrR/aonh1x3GO1cc1ENng1Jzj3kNKFrm/ARiqOdIIudMFjGgp82HFKvlGxc1pHCm
xiK2L930Y1PKWRgHtPjwcUh3yLcIEK+Rh7MFks7oTqGvB/p+asuaJkjge+c9lDHC
Gtahx0wlsFfVxB7+PySBCZZCVbxdxRWC7EQO1QLR52P/2Q9IxSUVW5bIlp228rpf
JzozFA4Sgnu7+IaM6/kgZ1+Z2bItSPO8agfsV2pKsayzFiWewT8PG3ASrhbK4kDN
m0p3ENTEW3GNdcktRgwmdp0Ko+gMNfT1yTt0uRr9lNsp8p9WMAtXQjK2pYfBCGkG
0+o872fXQb6t1D0NIEicah1wm5NhtJMVqY0HLROJrj0PvOHOhPLs3fKeGGSulpib
sKwgtFONVw09GGdJvTO/oH14j9a8V97dltFPTaqItHp19q93LuoLi9be4h3XtrkH
wHv3R+/JWlBBdGWYFGPNI7fW+e14twfGK6dhhTUFGWKwS986RU2Ps9Y1mVpe5koZ
qKZd3bP3Mq6ZeRiiQ4Jo4SalDdUCFUFodZRd+eUqx+sQl3gL+GQTFsIJf8SBpIK/
2Edk9/U4UAc5Ap7YkddxCYDBgnExncHXBHTEQgCXqquOqS70NPS0KOAfAe+2dB2O
ZqAnX88xsekDjDu1s5vMJq7qKcfMUo/NPsSbdHruoLp3tTooKMkZtYK9xaAwNb2Y
QfxYljjprzyuYvhvdhP3y9OF51FLVLkFCIgOzffmPZMq1y1QL46BMd0HOzaxnwaR
8UK3PkFP9NEi/v/cgUf5+eh5bAeptO6TAHCC37xYKDvronY4YnGpu5P6c3++ZZES
mBnLTONHHp/csNwA21aEOn87kOGnplTyXoxRT/VSVVBRBmdAaOMGwFt+DKrWfVEx
lhndRPesZC5KQ1fu5qFlbAElVIkx8ISWtQmhyyGWHIZMLo/FZUXwMg4Dg0VUQFXH
GePbwMiy7MjNFYJva285rvAymTQkoZLygPZ+0FZFqrjvXRVkPqdMNcYm6WUkD3lP
UxRuBManoBpdTiBpkM02166tgHYkZxtSgqp+oKWGqwfTDNvQmJzZqRS8+eCOk+VS
R9Vcl6odAebVly5qV0eZUefKtp4SCXybngRYzYrd//VtBdolC+tQqZ7WYD5d9/WU
7/qIAIdFgQfNtnGwcGE5qKMVhNE1Ow/6nvBwH2uN1SQi8jb1/stNnFjTDJbuwzyD
tYA+0QPkbAxsdzIVYDaEmCfnmkOV7wYtw2wmYLF00MH/uKmA4aKpMnzl8nOK5ad9
hwPi1vneySesJa5DDC8dMj4NMgR2zZF5HpM363ncqZmfzOSvPM0oTcD4QPvTpgz1
KNr/qjBxqRNLkro5lfBsRjpXhsDxhNdnQ/iw/HCHogHe9TJuVmlcKh9vuTx7LY/G
MZnRZXP4H3B/X5hzSG0utpuccYJ7j7Qe+e1YY7dqiSPJ/MiGacMbgJIs8OrhO1Zs
Uf3g1zrGYQtG4Rii2dAJuMNZWiVE01FjNrFnPqEpS+n3sRv7yXlOTCJMvErGofMn
De4mtNpcQwqC56KSSNGXNtQsx8vzzTQXvj1Wb/ACFAd6uKKg62z69u7rsSEw4mtM
h4wE3tBfebMYj25hFR05AzmZQksyNjdsGaexk9LTytMXA0lbC00WhRj35V1SUvj/
+70Ghtkgepo+GAd6XP2JyJf2ccDRt2sMy7M8ljdw1jLLOqtapfii2NVzYaR+W0Zd
JBefaZf/euN/zCg2Gs4yiCZXf55qvUWP/HfLAJqNyYCR2xr00tuKpKW/8CLfTdB4
a0Iuq1ZgELKn9ID+PwICAw9Vi9X1RcPL6YT9jkJAvE3L2piPnQZ8n5k5obCoA/Mq
GIy2+0FKpdsBYSLJVB4YnMY8V2KnlOh5mdBNYD1l/dahvLhHaLoy036CWFNKyaNL
FLo0y7W8ocUszdsANZz/YUIHv0FsiI3a1qo3OllLLNZHC60OOTejmJvr+j6CZKTV
z2NgMKMnQOm1+z66CGAETKm6rhMnxyBc99lA60mlYf0Pe9hhDqp794dwEmseCTgH
iEN+9fkXdMwT/4ZxtFH6q55mK72cBf+/xGt1e6t400mYVWBrYQoP5HVgGNUAS8Jm
j7em2JkFKgRGc2A7QkEuLxMv3PVbihRKZJtjfVyLzSVXflavEADIrE1b6/pCLuln
rsB9QKC/hnOqBvAzHeKLLkRQWQ2AXX1cAyiN8dBesH5MzdqQbPY1BJ1p8Uf1U3CB
wgzKdeZEUz5tYxGQXVkbS2Tdr4dVxhY+mu/eI1NZLXP5Uxr04WdrHlI/a2wZq/o3
VDIT0X0OqEhUJTdf2nc6M+7uuey0cQP2iWhp1eMFraUVFzKtJI9jDDI1JelqLc27
BEzJHNsqqm+JTxjibwFBY2JumRgX9BnBiBbNSs7ToDQwcidot5utlDGJpXz1Oqtj
RbK9jzpcTWF6DfVlE50XOklHxLr/AXEo5PvGejYYoYUalWy3x+zQWEtsjQVLGN2w
op9z6gQJbh3l0++iyS740jLhHzxpaUzX1qkvgdnZTl8kcKeJl49dhLZm9yU7aV0L
0dz3wFD7UkYNa2U202/xISNR6fqjT52tIYK7CdyegxY6MGIlYy1Y0lmXnLHJfHHy
DnJf63QV5oAUecmughBOs1J1psVk2VX/OuSj1uWVi+dCm4lTUcD/Ui8NktWQKGIn
6pkrtjwiWO6xIRajt0PpyP6LVyL60gLYuwMJ4RCD7gmpWcZz/CNh9iDDUlwdiWeM
60TZIygJDFukmPBMRHQgVorH0hpa2hV33TqauCRyzBx9aVEXedQHW9zqKmYTETQx
2EiLW43iVtSHzIUcAjhpWz5Wx+jirfJYaZij5Hue2TJLGGXXaRAG4yiD0JcmflPl
V6t+XNJjPfcGrE/Xh6YpmLSFL7xr0hwNG8VQvVJWbQ/Bj+21uTI5bldts26Pd3eJ
pm0l+Ao89md8J8NOeEOKMGDSlafebsDnPeXMGlfqMtLxV892fqB1IO5S6sAQZT6M
6/IxpqVqV1l1zreOGHsvbJwWgSllhCkAIBrS7NJz4SWdH18m5QGrSPHTkUxjQL8n
qdo1G+LnabhTBLc8hU03xwFlzSb3znfO9ug4a+hLkpcFTONYNazxRCO1Asjg5hNB
D8U5Re4E4EGVO8Qee++xjeVlqosga7P1G16BytRJnE2TTaEXRJJdSbssMGMdImkr
YayiNP2LZj5oamG0KpAIhguWROcw5jeAxqg8lC6MJSiBiVP2hTDcOTPYxzVJdN18
ktvsJl3in2zQEKn/djAMIk5qkVtbPSCnvoOtJDuwTi93LucM0tOYEOtuY/PqgRf/
HyMgRW7rS2e9oo4QXxMtlOk637Olf/OoSoO0AgbYayIKLPmKmbZhkQQUEjIhFhtZ
PQcKthGCrexlNikY6WiJpSJ8a2xocv9sRssnr8a6TkZ4W9QjxqvUp+hiZ31Oz8gC
t29aP9aRW1CGvf1ZbBPquSJnnAo87nrarDEmOEI5bBTY5+kk9J+8biituaxUunTU
qYjfYeKqyZeA0LAsNUsYQWjwNSnHHZG3kRjYq5YlXbROUNH7CqRj0ssDSYFvDFA8
mk79CZ25+zyH2BFsV024RKvUZ3i1NkkSpuIPmw+UK08FPw2znzRXaWtMlPWuiJNP
shpXnXNu9VheUvcp41P7TRovu6daCAnhFSehq9M2zOTorFtvcc2C4ymiMH5vsFyl
7oYPBlCmhdjo+hbCj0OmGc7Um3HlWRR6dI1x6i4oHppdI/oWz/B/ygzULi5IY/5M
R1FbgHNbau24uEbPSZu0NVpkMf7sLmMswns1sIqfazougPo6h2RO2T4KIrp0gjOc
DNMv+IdR3xSGL8ZfQ/G449J+RUJ4heL362M3WWtl1prKdWu00R2UI2c20qsU9R+a
GqdRB+ACh8dLCRyD24DD4rALuu0Bn7yaFlbW/l/twMKTOzwqDNgCOD6aYYSi0Ela
FazuuaV3nKRCUmCqlMhaeWpSRVydMqdQszeLjax5Vs5Cy5WhsANcrDkJiQZs+gGY
baflKEwBD/mxqAmkOvMDQlKkE3jdTm4Dv8iSAowBMxiIPARivGrfPl3rICYLo7Uf
eq6mpwMif8+xCudexJWAeYpTDPhgooQCAzfygRdZP23E9hurH0MzJhoNVm9UUyqI
uOImua42E6QhW1vtkUaLuPeMFxrB562sc24fKmz2kdBMoEIUDVSmaJVjjXrfI59a
vS6Knpyht9P906T96vOnWmUU5PkSUOMqy0mVYZ9EHZcDuKpBCnbZmvacymJTzRny
7mrkZrtI1C1jitY78BTFyMGBnRMwk0F5oPezyqPaHe07wxnTibh53aPDqIYn+jd7
u3Xtdo23XksfFKCbpCTJF0Rly1ILRbtl7S8OLaeJiRThfe84N9L+GEZKc2rIfr/2
7BZguuKvIfVapU/QP8WXDbZkYMXMdNGAaFjqTVUBgBXsxeo0rlVucKkRNlEVdMRX
oYCcrPlXasgKJWOEGEH2OenNdeOiCJS2Qx93qNBp81b6Vn1iWxZ7pmrNKeiv7JeL
ECDQrIK7yagQtxTUL7RNwyUHyhg6tfCAMtjxMnmTmg0y45I4v2s6JUU1lhlSupeu
P+e/hGsCPqTql+D0yoXIKBPabczm6fkHDZg1WCK6JBfcwCbQ4wtmiok9WbmJol0a
Ts0kUCbk9e5FJ66fY6ubwB7iB5KJfSMkXb1/sE8WV5h7Oj8CuMQaidcH1sqC5oC8
PLMJKjVH6+QWGrZuJlmRbaeC8Gq+wAlKDLFHbiSZylYUdhekdgbLeJ7jsKsyHsr7
KYoHax+mDGBCKxCAzTxvTUM2jN/Jie9jzhhKXxcU+kw4VO75DRsQLK4g8Y04u8De
6RyM4TpCM7vJgIUy7WVBtrXHh9Sg4vVoQdlAKddp6DHIwXKlHsU9DklzdHj9h9ov
dcmfLDN0+32UAH7w8SAzLOPb1nzKSI0M0jsdc/cfBVKJokSqrmh1cAdrOZoRonTO
oUF2SrkZ2HF3Pmr92uzUUg99AGMD+JyQKH/bj3NqiWuMlpX8SUKATiZ6uhFDNEJ/
5yavHle5Pj1SWyJXbctDigTGlCs1eoHV/XPBVuNCfHUbHn5nchhyqXj3JGt4jdMC
zFZdM3rA4vm5Q5cvuP5lWyp/FR5I1b95Vgd4/09pbFS3fVzg3rw2lX9RfveJ/OoI
3qH07SF0IjAfWJV1Q3MZeIAFG9Kyw9GY5su+kVYoUEwqVn+4iCPeEi/2jHKUIuwX
Yh22ef+vC07cc5yYbR1J8wLMY2BiqwWfrUOmQLHG6IQVU7QNdffM6FlUqq7uXx5q
e+4sm8mlznsSLIXvcHqxrgqk+HyohFFX/9h/fI4cvI7HHle+AtGX18tVvOo/Suix
zkyaUECWpLlFVnv6UV2C6DuQxgGsEY+/+8GowaYwbuWDJ1XGGD+C0lqsiMn66Cnk
6d9GWVi9XyFSVDvwGR2D4GV3meQsHWIwwwIN3r+2BCqFiQGnhCyQf2tI5pm1lifo
sh/hF9LVHwIQTVl+3TPROvJv6Vwh4+KnYTRhXZRU7e8nyVuEBY1hX8bBQ/iz1wfY
C8oa/uWIm9ZA5r4Wkh1rJFt0jRm6Zyt6SM0ooGYv4h8Gxlhle3GqNqo7h7DtQha7
qVSZhY7YzU5n7RpudwmdO/zJWQUG2J3iRRkHKg88+0lZ9py8lSW8h2Hsp2zfb+0H
Yajk2+5jBYO5hZspYRLZTChj52CG9RS5lbV383r8Ymv3kdHuFAx1SdGPCjcYoosf
1HWM6XWRSBHE2L01nla19XRfT8VT3M2Otkt/Rtq4whOK/cE+JCi/LHM6vHf7MLVb
bR0X0Gq5MXlypV5bW2Gm84E57IgWJA99eeJ6lNiF7o4xCQOLB0s0FHDZgg9m83D6
RiuN5mhMA2CsUuVB+rxAjH/7hJM7AWqwxV4Vqp9646XSNbKIT8QTS8N3vM0SJX4a
uH7mRx1/M2VBUBYUE5N9Y2h0ZfKvDkc4FEO97SraOcihWzxAFdJmi/P1U9O1Ez4p
eTbhiDQMnjVgZr2p724IDSz7P2nVHW7A4Xx1uZYnvYs8PGQU+clsxqnqaoZo3b3R
TIfjlszqFRmIZ+xWSWvXTTUwWS0zMZSQ6tB/Dr5NqP1Pad1jhMnMJ+znnDVdPENI
hPQcvwmDeLVuA0bhnRLnMiPcZV2MdqEOL0igl5TgS+A+/9pg2ZbNNb9LeQbwB2/3
/Nx7t99LJ8HsCt5B260GqNYjPVq1hLj6/oml6gee70yV0YNJANxoD8GiHqx+ZhIF
FGtOmzk/v9T7pGh2QqK6z6t7XISByOB1YjNKJlBr95y1t/oxHg2Cizo/Gl5DVHRE
oZLihsEKFIpCQDvVDlr80tZOG6+UEtorh55lU/ATPQmAJwLguY8JMgjVTlOMzqFN
RE4ThSJovq5imHHB9hhiwTkGDnjJMfHyMbd8nXSzdiu2gWVFxl7XN8guBy6KrOht
/EyqqqITc5Sr6QzTF/H6VIUQNwEzryyaC/q3fgwOI1jNmijCCpFLgrVe5d32HF6M
TlDhfIl8QXWxPeYQNq2bTvpKpCWSEZs77mF1xUkPlOUWPJwNGwUU7OvbrHBzpanw
If3iYW3VwRHFnz8A4i3Qs+dTKC4oaR/OuiVR8PnPo+MGmzsdlo7GposMMfnSA11F
MHMerAowXv7ylzb4/0YSEAk/3KbhkDm4V0VjbSXjn7dpVjEUSyyMhUlOXfwQfgbX
XC+tWn76AUyAx7JIMsZvZMRikEYNgEzVAw7ihXPi6GyA4l4bQaxPt4anhkVNvxot
KRf5JMOq+jG9B2T6R+2LpYuLkxmsh3DWPyzLAJ1Mjkx8lEB52fPqntbU4XBN0bwC
QmTyK9QJYq2w2CX4LCrka237oUPpMUpUUBIsV3V4RtvJnx4lw79jgwApB8sH0Ygq
2fYnOxlWjqA2VHHDCgqvSwHzzf2F6bUXIxnTH8e5jIiq5ADuNNoUhglDq0VvIucD
2yfY89ytrJieAPWIxMdNY9jraRh/KdZtoTsY8ms/JUxO/3LGDoxV/tRb/UTuB4d1
SPI4NmU62JH0qMSLxwtZFWcOeVICQ1Tad4wp4dMyOSSsKkfWjhcpSroJ5I91wULs
3cApbHOvB0bWvREOJBedorIfVsCjVYezRoMtnoCSGurE4FXiQnVTiImJQ3QW15Wo
HncHPHdHIvpjI4FIl25zempwIp02SuzzMUl+M33kpbMoor37GxYDSvZiTTtlJQyg
FHyv7zPd8s+xe8pA9Ik/rOWp/gun5iGKXz+P1iwvf5skc/smYo7ya9H2m+Y7EW8c
hwc6s0RVQdhm621L6LiOKFRjMWFZvyGKfDJBLzlToJAqogknpgb5RB7YUyi72RPc
T8ix/X514lkrIi1t+RI9hePRXCDTIg+ZSVWz03ADorj0pDAmv3CS8NycVAyIsdJQ
wk2IEwumnShS/jqkE1PCkqe4H9b51t7MB5VJp6I9lydeuTyUOw3FtjiSEJ1710Qn
Uvmn1iNpesR/1skF04RRwJ2cmy16VL6s/gS8rkEvCytAE0BCUtxyT2zhiUXwZPEn
Sun3o7oW4IWsemR8JXnLHHdzYd88KAlPGFoejcHfyCoBzX4WDALvHUOKp1DHgASi
CN0XO2q5NftwYll921+7d5mpH4wO3Po2jsGHi/nXxLNryuj65LqcucFzt07OfRoS
MtbXdppa2mrwCxk5cHpTlkTfiQOfhQkMEabenpfA+HsW1NU74n1pnvluDROh+3A7
YhmNHzYPTaElfZGS9uoDF8MuvKA1NpeiRyPHAjOUg41TcLNK8F0QQfmdLH6oEBrh
x8GaumkyhoaOftxilnw+MmgQ3ZcL8kzNKFeIW1rbNMWVpRn8lTD+YWRc+2vXL53V
8IDtrWCU+0/evdQP0r+/BEwAWDXK87LNxA3hya58yt2+BBQPdCpIc/1nJZx1CBBI
hjqMfaTXvVTiVQn5+SYZKcLgZBHHW2HTpBMKMw4R9c6slwdNGjvEeKxY3XFJL3s+
I5W9JzAl5CxZR8N9uZmGs2AF6SJ3AEjwhm7BAxvcF34otM90dBBIlYsvMLZ8YHSR
9Om6710RUEY5v62mZJ2Ip9Q9JDb/vGqM5UUbPF8cyPtY+bjbT89koM5Qsp0u/9Sb
Twp53+6lwQgalxJ3SFEBoJQdjCyN431HDsTcfIdAdncvsUeaGtU0hOminxC/ayQG
0kpyPZtlBHXFtkQZkEiEyRl5GWpuEtyqGiOAkZA1bf0Z0hLQxsYyvfHRXJ+gARBb
olCkGnmjsIfZ80duwEx+Yw1HaIwOZXgvrNeNesQHBHr9MmYtW1G+cQJUgy9tT2tS
skSCYFUJvO5ErSjpRslb8tlh1upk0ZUUA6NOTGvpXf2f/4RbOQ7wsBkFBfXCjMXu
OWE/HBoXrAIzcT3sljyIxNol2/hiVpDobwHePWyM2fpow8anNo8gu81tMOMW3NRK
KSsr4gVvia27ersRXEDmB7+SvZEqN1h0MaoXRJgHdRKilzQYdw5/5oU4yhG9zfSd
ntapIB+d9k+3joA3S3jxagNrWtTZvkp/4nbrtaC+RaA3NOGbTCq9L5XZQ++aspVW
mtpgYnvXE/Ga7zqMOEXxsJ/5R7atQDC3eseYqRR7NgDOmbx8gsPNKnJcgylPFOEc
sskZsV+fPGDB41dMOHEU1OiIpwuwHnh0jVkDoGo24ssEk4EHZz/gkzHoLESZx5JZ
9+R9GJSnWjSVzqI8r+CZ/KFS3F6AgqDDdSQM5fKzxndKeZA+Txgctcbdmw8klbNO
upUroUyvAfGH33x5vtPVyc+MlKT6159MF+eLE1bLNy+4u72zf/H1GOej8SaojEfJ
imqAwFOg1Qo12yYDSvW6re+MbaZD3wB7IsE6vodBdTjhHbXoikaHGqVLT5ehSEWl
pH4DY99uSCCkVel4h1XO72d5d0nOelP9gtzWpZfql77NmdOrkBtuj4CS4hQOh1KH
yUNdAY1/8qphyKgLFU0bIbb1mgVpIsk2Mzp2VWKl4l9fLOA8YsRoaUNZazjSgFn2
0TRgZHA65ooiFkRHU5xxYRFWLysAb0mxtLsscK3VbkZ1z14beGBL1hBvju74U7gC
iQx+IpE9HS3EWTiCAgEGATPyAX0neJdOT00tl+Lq+ey99kONYuoAwtd4DSgu68Cz
KabzL24c/X366A57wQuETPBrFM4nVTy0d6GAZHo04aAbHk6e+tiKocsb0F2IYWWa
5Ct3HgVAl8lAbvA09UGQqZTNidtSgl0RwkYvEvu8dmIXEt9vQMuvi7p/d3Xcl/dU
p6XU3iK1e5N6GcngqrWKV9uZWIZofh9TgGo+2Yy5pWvSJAhQqY95ufCQ/jornLlN
RwdAsJ9CgG/l/O35yrQgaLFp1andzJ2nBZs91zXY+CzTPf5P2ow0+6S0uIU8hVPO
VNkIFRAVTvAyoyGECxcCwLq7p3Ic2B2V6cIGuNXt7Y3PvPIKPQ46MNdCFGos9czw
FQ7K3YuKKekzpVrutUeS1+0a9bWKCgZQE+Sq5tY74CgbQ54naNwLzxNPq2e09aV9
9r3UAm3jtgzz+X6+i6CcD5WFeWbCN3HPOKDbVjZS8/T7hLa7nL9yG1TUTOLD8C5k
twoDnGmpX4cJouqiFldE/R6w2ZW8mxLVqC6rqow+GFMwdq3JFvEIIH9wlCLd+kD1
4LWDNS6R+A3+YhwEF9Mzb9uwU8VOEECM8AkqOM0K/Lq9JH8Di286uBZSzBCvDALR
ZjwEKg9LKIhepS3jtFtUvizHGAoylb54HfMmw55dBdDc7ZojbPJIaIT2OAOL/IWi
Qt1JCh7g1tgDgSv/BBqxSaZEXqzIgRfKkLBI9xIv0ozYbasxiFjR7d7tI5VD5nSX
ZCQ7wlmwgfg7x/3u7U7r977b7I6JpkfJdujca/KYpWpzhWREsKMh18Nu9Knm/9pw
0arPO5InjeOWYXIfp0n12r3QdbmWRV0DrJkdoVZhOvUtIIymRLsH39d7m56Akdxm
Jgk8GkvVeMBo4OS1tZMvFBapWBtv/Z5/EvHG5XsnJ6IIjIoPWgbs7ncUFAmHVvRA
7ZRk5NkWs9GMS38G6bylBYOgNyd8+8mQQiyb/rxw+ZXlB3TnapfYALjXtnNN8aVg
jXYSTG/lOpSu6MEgGT0MqiK+YByuM+MbkvxLzILwmEIGQzWDFZ/hR+ORZuJJyTPq
Ugmi0wn3wRYEP6Dn64kGtoqd8Sg7FJre4W6R0Ez0sRe9IlYhIEF1AzBGBTxshgHH
BkDdj+2Sh6BKtMIofAQL6JS0a04rB4GSpiXQXRuxIZsmnPr+1hQEedqpRtMYrWDT
2s+5tNkOzawIepkAay4Bs5g+kZKmRoBnBlIanj+Ioz4mNrFAzDG/PvGYQwK/cXHJ
wocu9MPtBdyNGpqrR4Fjg1zDHE2dexckZAtpQof10kvLpjmk8BxmjD2TGzvOS+dJ
QlxdOJmdp+1YzjBm7UKz5NpzmU5DFf8z4MDGEqkhF4I=
`protect END_PROTECTED
