`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
korMCLpShZtRKFfs9og77Z0LrysfydTtzMJ19JjoxOo2lhbbtUrPuuFzf232mA5O
Udc+pyKEmF9nmyRim33YTv1L1SHFmQA60svRbsOtLe8ser6XwS0YPD0JXCeQDO5a
/fNtpqvvDzt0dLmnwGrw4x+SJEBKs4VMxsWDubmrHj6amFG5UCyefdtNjcipsN6x
ODquYe+VHezorhhsGe9adl0ahNSyXgxhej6eIWqbO29f6KgrZbd6TzSc3lW5aUWh
8vxNZZ5OMC2letOHMEp0+cGIjOgRkLR43PhNFtyXJJ8+fiPoAC0uWSycuQhJWeM/
V2JzzVKJJAtsEaiXzzXdMSzW8PL/GbqdyYe2+RTFGFzgpmN7PF3C5n05q6MlQPKO
u8KDvT7IrRbrqogzNxKfsJTNuprXDXESbafnWbiDUGPGSF8hYTFXtOrM/11brd6N
Jcd5w8WI5f2YFbAHyCKIpoVFczU0Kp9/Br8QxvitSAJ7GkxwkgAeANZlMZImDrXs
joqochR6u4QPQS8H12l9HMxu29nirdMtDWPUNCqx45wv2mFcsJzCOt3qsjOenyr1
MtF5/pNDcqVg1mUoYirNNs/cJs+kNXKc7U3kw5F3QvWAzZXnhbN0N8b5+TuNLnoC
5tcxeSdDPaAkOx1RDStWtqOOt+RkpXw0BWClCJr7M+83gvjTgpDSwta57QIUFlll
HEbtCsYzJHTdQMmDmdkrkKSfqc+nVqiR2FU55Z6MiFEL6diosU0lE4O3tJf1Ni3+
M5x4mNmxpxEW0cSIRlfg4VLyxKmErpmZAhiYjMuh65pd4Kyqqm8ydzBJdlTyA5YL
/LByY5zm7MFPS8pnmuozUfq5tYT4g/FVPelq+SldvhZXdX9A1xj/Ndgj7PFiCxrZ
iRoN1FEDE1xRjtcJJFlN4dY1Jnxpc2hsTfIxRKrXGTEwFiI1jFw5lFB2oe6H7Ghv
pBPKBjjl5GfvsMdlqIql/ny5PUxTelo2A87c/u4pWGg21/tLisYtvMm/gh9xgAUY
5MTK6arvOxJIyTc/OuEWH5c0Ul1pYHxyFjatDOUUvdNLr9w45NlOtxpZODUF7s6i
JgRsV0E/xjY+6lewbEYgeuZxPIxL1VSUlQCW47NG8nhO3DI/ON5dtaZyUVlzBzTX
9U0F1SGNyQ9QxPJWk6g+XaWCyjq5aclk6UbnUtjE1mmUkeZ/NphNs7u7fUyfeTei
gdYHFige0kUZTsyRjCLEZ2vM1Aq/UaOrTazhhsG797dZXfoz1JwN7V1gjzM7wQas
6k5Y/DICaz10ipYN1jKTDmnWzBOjEa58x8x7Z0fLHm384npjv3yPYMI9UeIjfv6x
lq/2junMKsUif2cikbYBDQ02D/UsREBa9S/7qm9UQ4P4i9errfhXtw3oENdO5xzA
JtSGg4mddPO7IIAFs88AxM5GNgo1g+pssfl+rEmIZ9Il513X2fLPlyuX5BfosnvC
E00qiKKgd4cYW2mLQE3kkrpTsk39vil+BwfotdGQiKFTsLHBlWyisH7QxqWDVQfq
Ael3djg5OIUDmMmrInuSkyn81KOzJN3Z14Z3zv+Kcg6zfr0vHaNUcsvhygSl8An1
QrOj8iOzciR6EJzs5fgj43RBX9MpQEQdd2zoaOyUMwof854NYZEM/2qTpDQ0MxLb
rA8Wjq6J9MiOSJMPfR+tHDksjkUX6wUvNlWgUlSx6jsqaQTFg8iPzIrXjb9bMB1+
cr02GdRFtANE2hGgMfFZrrVxqSYBhu+2C8US4WW3uUiwMMdXjlwFUHjQbLlhdReF
/FK9WD6yaYy3HBpQleB8HNs/xwl+Z8BFnsGZMrurvYuxHGo83kj+j6Exqt+1D3iA
vrmsRYewm2Gcsp+Drqub/dCo8H2os5uTaZKo01ICmsVzK07NAo1O6uy57ZCu64GH
6ADthLd5s5L1QBPXYymd05p909eb7N8o7OadrQovb/pn3NVxROwrvLg97JSifKCB
7+q5lysepfN+AqmS+T9RU33ubm/dqyUq9OMfk/cgotSsoTZ88d9ijTt+IAIXNxeK
XmgjZrWifdqfe9HRAAr2OK0cr6jx8D7zu6Guc8xBWqZlFMt1ZIV6uN3es+1sASB8
dw4M7APAk+37qDlwlTHWhSLy1OzoUQy+EjpMec74wEGZ7X6A55FhSM+Ga6sFJeBd
`protect END_PROTECTED
