`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FEkYg2eDf2aYjQPa6KvzoG80oVFJSoa6mhg+4ZkUmObZJDF3uJs2fyGaNNoDkeeD
QawfIAWQAIMf7sSNTg+j/RSuqMa1Hx02acNk1sky5/smT+mt0xDRda0gTHceS3V0
VUoRALSl9ZDizPtFEyvqn4/V+5Ttl8hCMD1qlUY/JsCEAWcSfHpTUknDMzwI1aqB
lNgJZ9473s21ahHEhAaqVt3VIcuOo1u0q8+LypQvjUBdxSb9P/ANGL0OXa/bKsX+
6p6pM8Pl7RjLV6ogroE9/1dYi5BBd/7xeWZOhvLrk/HrN9Rc08oOOgpg3QwfbpW1
a6wJEHrQkbbesHtS0z2xqw6/pE855Vt+3Xl0Q8IKGQtYqMXobSZns1VWGZqQujCc
2fhj78ZzURBazwhGV/PuGKYHizVtWuj4l7N89++QXtsXo3raZV4F6qfi532SZnHs
798/Owtj2fm4Lo/4CSMFzUVYw9XMXVl4tt8ClPMk3UMfTvgHh7TciXoBjpOL91BB
YPYqdktgQuD2hTeRejAM8A2OxwK9GjU7uzxjS65aDABIgUn7DXZwJk6yC3YbxmE/
JjTAebIGXxiSsE8u0VGBrPVOwwdu1SQrpHPSE2Tq7S6hFTl6gSNdxhraynQGEqYU
RG7NRf7TNeel0urDVVzr+EjiP0p+BMYVwAS0UxYsVkCGbR491MN2lA7XYs4mkhDR
mSnOtRzjYKhteODTZTV5flIhT42HoTk2Fi2phrRPeuAl/MoUv2MzVbePxq5bWenw
0OfR5FsPum9MyCXZ8fgsyvVWCIJ7gaJSQ2MQSmSHw9pQPDKyllO6hr26UyqgKjOX
ri1X+bHxGeutgDWIVs0uCRz6wKCetzxAax15p+ajB7FAhx/RR7VgJzqJ5C72U2ly
H+8bZaoytAUCMM1szwYkeXZeEoZfIS0JZiItKLYm5L8K5GEUUfyR3f44MaU3S7Qq
Yy6obJF3v9Bz7+Y3owAnQJ1QmF6Np1hBo/GEOo9O/UWdVHuPXuRy3kNDuOATblOF
xum98FAfcQnmGd9mytRD/ZzGwwIojtUN85eEDjSTfz4kMfg5wEzhNoeR5ISg94XC
ascJkFBtQ8mqXq4fJ0+3l2nZHYmFEsbfFRBaXr8CAQcylRQCuvuPv7K/MXXSr+Kl
LLHmgfALd3snvwlR/c4ToOXEtTNl5Y7JsHx7u/xxlTImNTpyjgGno5/8V9/fWPxT
Y7RL7YSu7aI8Q+N7XEg/1ZTvMoIXGMNDHU7seiSxB/ngLuesK9zRgGrXYdBNY1+b
kpWMYTa3EVbXfEb+niGPAuT978DqZxh17KoezOyxa3Y2/TTD6ur0lAHFCnVca9ie
vfLcjAwypFaDnPJFPF4Rs8zV8rnUi0XZYZiHFwMbujqTmrXmBKTsOWwWPRmX7wmb
D1ul7f+xFiKTKsaI7V0n9d9i1kjnT/MjopVDr7JYZT5LI+lfa54bgNzq98rKrZU3
pGyBdOcIThWtpAsmE3MFXfoQfGW1o4wsy90qUM5aj/GnImG2n5g/tLoCJ1hdBIZn
eCygovmKIdZNR535fxBz06xQugFqUGumibUILdCFRtnbAedeMhuiBD0uuGzh4veb
gjYlTmtXbPVbJFyUOUZIZlp0QQEl0oss87rVRJtLB4vzWjpdLI0GEaVsVrB/lLyT
uRE4S5AWOQwFkLR1Y7RDTwVxW7oFMSlSX7tp+Ufww7YOg15bOxQz7QYyTenFFt8F
eB0alIiMgU7Y0LSKTxMLLrSqT2AhE7i/oUnMzppS7IH7ZaNCGtj8EwNStk9E2Oza
qI96W7L1/wgrxlzUoxR/yj6SLomVC95MVWx7Of2mw3RbyyoW/D2+FRMrQ8uA/9s9
PzLmCR3dS/W9T/f8BLnt/xkJ1yT5W/DSqzbtOgdJw2zNqBUx7gd3rYvsafLNqR/x
EwzC/GTYE/2aRLZ3zCxZyHkMpXgzKgJwYLZF1uiPOXI5fjuhMh2w3QF78YIAIFdF
VO3WH1qXMM1emx7XCYgREleWVExswwjvNZzb3fgpwttTVVDNuo2xV8+gWT/B3tGF
FV0XD6xBncVrB9YaCIsYmZQ0bqtjjhKIi2phQOls0yH/dYlrZ39FX6diPwPfMQ+2
cU6AtrvcZTRrxpTJaNQa8uYvuqILpS+NmQMFwiJ09SKxcydXWzTAYlnvjPxOxi0G
4R7sBATNKDOapz8kG7o4AIh0r5qRfh9XpdZ+hYSgV4zW/D4rdg6LkkUkBf/0rHJF
iRcMYZoX+9+pvc2gKbU8BxpTMuWPfAXh1poQq2BN8vtnQQoRk4gZXqqVDLhYJpoN
50bC99JRJyGF4Wi2CBxvjY/x1stUWoOKl9LONqprBjx3jTta1qFFXyo/PzOG8QW0
dO9BnP62Fxoj0saeKuGzEt/l8L/oiH4eU6GtMUQh4JmLxNGdACQklt2YXS9qcxWm
mfQdX27R22efER1Zfy/f2yvliRNP7YKEHcfS5Pwc5nevo2JRngdmQJOzO2abMdqO
RCEhXAIqJw5McuI7nhS/Z6d0fYM+zsmngTCpR4u7cKjC/e2M/i0SbP9XijEfCOi5
7mdpbqUfGtBB2qv0uGxYtm/xfhH8nI4VYujpK/ogMpFc5t/QTNZeFgTsZI56pb0P
IWFf/Rj2EirJ2+FtYA39CWQ48Q/hzrdRu7gjxIJI+3BukyyphjjJtIkpmIODWBo0
Z++7P9tSY9wsJ/ui5njACPVU/U3eiT0MYYEAHvfp+CKyDRA6/906D7fRSpupZMh6
mb7xvwfJM7bufGHhIE7VNjNNqWoCD8IHr2Mtrl2hUxvukiC0o8BfAmf7dVcEpmaP
ngfHpLplWVKLje2eOl8hYPeBF0j6NS5KctC7SBMx21zVqaujD+JZ4ebsqZKPX7oD
naxIaitbyglNC7QiFakJGA7fFBWPguom9eNvc1wvgdB/kiezb15z3VRYhB6QsMNO
uKhggYnpD6E+tS1STDIC61HA/gi1lUT8Xpc0Ao0tG5CGzxv+gmKFEiOwjw6A+lP8
d53t3Xk5f9Blxa5fmlAo3Jt6oY34kdifa/a6RizshUBfJXRJ/OYzecGe9NaOUN6r
JxVUE9vHl2e+3AoqOHzv7VxEDZvzhKUsSes/wS7O9F4V3L1S0DcFwa0fIVeaKF3N
T25zIPJq5ts2roZF7zGTS9fI2I5FYzVnJpkqeYNHc3KAtwPJn3cpLOR47C68l9w9
SMg/YdDlvp9Z0NG4IIlp+Fl8HBIkexGkhwKfQa2LPEGEylI1AYvWJtfGnEilZnZU
CD5YN344aHKgEoL1aQPj5gJIipXqPYPZftg1+r7NdXEP29kQur1iKuPi657d6D28
hr5UVkaoXfQLSc31e5nOiXyP+MemNdxrPE4FT4ZG4Ix6FBF4MtY7Fz2qhxbXwbgj
mJhr4EcShst+FPWn2QZEjRTWubrRBAcOj7uvtcpYho5tatiwggBsgTLir4jsVz9L
TufQ+/o7dWZGdr6mAB5rN7N+0vQlt/+01qOLatzFOwGFsRP6yvJ9sGWKevR9oZrK
tZrPgZQVihT0HCTHOjskwT3nUEL7MQX5F+nTI3awcSV+8MGLjGjU7vEP7yZd90iW
YT5cTM5q5PlwY56hQ5/DW8OyQZp9716B1OYaV4Z5nrCRD5b5lthjeF4VQ/Tf+ixj
A2K9heAiBRoNQ+4v4/NlN9aAZUieGfyGvotGLYpshKEgMOblCLIgka8ny3L6m/Eo
Tj5wKKcJXB97h04OIKK8hQzvjPqNh78mscjvzDmAqXiKYN6Rz0w1dbH+Q46+zJ2P
eQtCIPnXkn1eqQyAnHcESlG3MbdvYtFHCT+NJY9pTFmhVJFAmVxsJuUacB90tM3c
for2bAwqNiMKa7zgxl7g/pkcEYrvNoXlGSzLQKatvaJDwoUGau7mBQeNFnBGHaqs
3D034ZGJ6uAukyn5j9tOQXBSoiDaXAcqHJwXcni0LITkubz3dBsBgfNHdOT1oxnS
CGhuqwiETxLIuZAGanDQvX/ICOB9RdYMjmpEsvzI5nakudzl6ZdasqzookrjsdlE
d6CXTTRGGOg40O9K+Ji+WizmHeJ4Oh1tqShjYZxYs4HS3RS/1ZI1DfbRYZp0Yj4b
IsvZUiHp1kP+I1QwYU7knSFe4Nq59HinD5Re4g8YoWgMzPzyjoh4PiA/bGgXnjEr
pqHVwRpx/SYf2L9V7ANEvVNq0f3BvifoGYEuxbqkPDzW4Sf81oLmgPHGKWMjhC4N
YyV4K0TBPirsP+GBiF+k3lomvgWVxzpw1mIzLNs9DcNQJhor30QoYjXfo/yND3lV
fds4b9/5QjoEwnCDWb61b+9HNtlI4ti+3+PSO5ZyMSQJnrmhv4jOYHeIWqdRGJGC
OAw1B91Gu93zwW2KCxZQkxaErrh/Zi9zobomn3uOY9D78NKLdvaS1HxcjxOkuNop
KM5w++HI8LLm1XxNueDe3LhrCaGRSFXacTqDyYhJiyMsmDLroPUUId8MRumFk+JH
8cUyFQk1/PqeovroP1WJjnQgY5HnVvig9ZKxWEeie5ebXjnr2BU/TR2nQpYWmaY9
MaC2JFP098J5nXRhmImtcoIZcOG5wsiOEGnDBbluYlWBjY7Rl9IJNQY8KQQg/9nM
m/H5MLbJblcD64WyxNV8OMLV38vgVeBa0X2uhS3w9pJdd1MhGZ4iyOKwJuLtQeoZ
JZ6zmNJmzQbOWcbeT5GBT+ie3rlnmkM+b9YnR5CYmDcetXEy7IqeK7iq+Bk+F9XB
en4uyIs5VLV2es9hMZfEyEGPpUnAS7eTKpm0Id0gwUHnMRKig/PzCaBMnz6SOgKy
zVxI6Qp+4D/c8BF0vWOUPPemLTShav1NnDkTVYONL+pDUEsMI4WRRIpIzsY4w4W3
vqRY+of2dkOfObQbpsdwrXWH9Df76AEsFohtgbvx7CToWafZ00w7ylspvJELsl8z
fxdlMccAw8FB6RNlw9/hxvBaOtdpmGVY/M9QFTDEN4KKZYI66/yxFDyShqmde5b+
Mz7GlfJsC/EIWm9xtdoHPpyqojvx1NGVTObAE5iZqee+WJNx6D82P0HnzsNDf54m
SlFjT1LcNdEzxcmC2qzcSD/i2GhmtyzhpKufjEDvKlmFyfihEZqM0XX85Qp79yPz
gKaCAqxJi/f/QY6oTjZALjPijHCfhJYqhK7EXO2AOAHIFlqagz05wszwVkmVHCGg
PdizeEVDZgjahmbExdr0tYViqHDjGUiAuOChHawWeoIr4W20/V7NT3Fxizo5U0zy
Haq2Dmb6Be7FR8KVk21KQreDmIw/6RJWw0yX2TD7moN097uGcrwZRbxLaD9jR47L
mwJQig3AxWoum5B1Hemqz08KL7HgylLe8zOy9ACW52Gqw6pa/kQFTEvdHabh1TWy
E3lRVXhBAzVRJ9CTGK+fstxEfhR5mLYE5kQRLyudCOaRev/Qk6ETsR95G75puvBj
orpFy7n70u2y6/E68Fv8KUg3ssBvdu3Sza6jCyRrUm4/8ATLRv3hRSMel77hqXvk
afwgYD5HFaCknDpjPFgFsWBAcGg97MhZeEeK/+ojnwXue0eZZXx4IUhDPKqeH1KN
nJm3zUiNn0KbpFk3Mg+slawbbR9a0nkAfzSp/CioRYpp1uhD7ouvJ6RiHERizm6Y
a+f+ELAQrG7YafYApOy28A/KorO9j4u4wa9dDBAnedyKx6sbkIiRtwYOYHH46Qkb
q1UuGMZIyHLyAdDqA6IAA5QImnETMR/KpmsGoX5xzga3B73fG2gE52vfRIyFB5tR
CE/QVplPAhg/LAw3VYM1Lsn1QfHJHYiOt5kh6YcB6EIry8USd9sV2FuIMl6avT5G
NQlD4PEqBPEFCijg8QVXzVrqaY84aqH06WLCprGQPJTY1P2WGmauu8kvZrLIIcbI
BL++ISxiOy7k941kkCZjvEVK5h8aSh3AfXI6chNKTGMtefMufr6DKGF3Q8dP2Ga9
mBZWZdjPnnchEmXcPOp0mKxR3Y/huFYjBa/5V5uSIFA+iXmOIkYzn36r9kQqZ/GI
Ge7aND1rp6HWmP4nDB7j3WJS9y9AcZdgFXXLXUfrWT80wApWVjyyMyn+VWZaLOcD
APhKPaWJAh1U4sFhVbvhhmWeABOdC7GXvHOQiVCBY3uoIsixjxk3WQlQ/OFXtiMg
zuUqZRUGpNapYw7CqgeuLaruV5YDLSn1z3ybXVG8kF2ZBG03JiRqUS69T7FxXSKE
ZVIkoVnNIkqnOQGvvW/GbU1/2GF5fAoeg/Ii3wsNiQ4wBv5y5hkQpXMp/FGcgbG8
WuztG8B4BhnE4HqHeQdtkQPyNYjgqL1rGAw7MYbaJtHFmn0wcR6ug8GMwvBInijE
VItwEjcQkxH2cITaOMFs9VvvLBCG/srCnYdMfx1jL/aAF+ZSs1gKM0NFzNJ+SUKS
qIJ+lpDHiWPxWmo30Kb9GzgS2qJ1UvZGAzFjcw/ZGMeZdSLjGhpDIBYijvLDRym1
zlo3zu77RDVNonCbTs/RECFTwbUCZa5zPe9+uvyLo1PRdAW+xKoVol7zak5aMSLh
vw5P9zE9mh0fq6gtRwripT33n7g0wf2P7p0WzksPSbeH5N4st8yA/ALQUw8t+Q7t
WFvz6PM+PltepJrRUAa2uX0DdFmGS1PKISnsuUu+TPlpZHhYTSw8U0Zr7IY9MwBu
9QaKlQoe1H6/vFWLRRHMxOqBGvnfYVdPsraMXu/3IFiTwP5unQrwd6Lk4OcuqG4I
uNC0zGVvFFFm+cDQIEcMBkmzZHXMRzVJuoBP90KTz5/JCoNa4NOTuSCKdx5YkzO7
D4Xwq1UkP1u72CPt6iyiirXccNTIJsi9b4eiOyfKkepxDc2YXAGHUY92QTxvUP1L
hawUP9L4gN2Kzq7VbyvwJLbEQC7KVZpFthUAPu2JguIMDLmSWkYs5/CjxsQHkSGn
+14/cExsM3Ji1L0Ph2TviV25dsxL12/wmiI6wY5ubaglifns6pVjXhLir+Bgv2kz
ZTcGZc/TMtog1/LxbYxZdQZb6C1wBlF4cw7VlpRvfAY5EYiWuK0ipMjMUv8hfPCz
VuLrm+vUnjVZql7wKHxpTSv+2GYpA00FCqlua8+H7fCXoXjnM1J9NmfzNJIZXrej
x8yW+50z5MY38tWQykRDaIrDVoNeT0fak/MLmU7d0qTFDi2C3PBqggYuf+iGgg0q
zVCr16tM6gCYVmbEa6ppZsV1YGHuBLJIat5BEzciDz4wBROekmXKchQqcCLDzHDZ
VSXFTqi2DVx7Ga8yPAv253vfzmvv5zYpq2uEKzD4ddicYQsWsMy2B3yJIvJva4xX
LhU7uRK0/qqUZnPlZcgvq8FhpV5iut5OUu/9jTgjsto8J9inmyyoccieLZU+7xzL
Fnj7SITsRs5z6bBUJusyucuz0vspO0EXausydA/t6CSzbHS2YSqsUD2sflKUyKr4
8nw19J4Q6ypMsXqFEnPFO8eIm9ibC5GyfEG/DCry6dA/EDayVpg7fjgWrOGQl7ZQ
lPBTID4Wtx24GyrgtT4TiTkg8ad/59gFOFhn5YaNHiR1p7vs+N+eFWQH5/i/fSeQ
FkJGfYn9myGhAYKYmQufYR7ODsOi0fcgEdfHe4UUiwQKJ4jKAtGuc+Huk8OU7J1l
QrxxnuUmJm+Z1dy9IMg6HcR2ZfABuT0o4lknI/0EWO/erY3zSiDvxtrXQv0RwClf
Cljx3u7uR/HJ2vlsCnzt0hvYzzmYhYe0eYiNP41eXHB+qXxUKqFToFmUiPOzZUgN
uR1F8HuiMTLQUxXa5U5nxA==
`protect END_PROTECTED
