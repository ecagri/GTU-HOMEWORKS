library verilog;
use verilog.vl_types.all;
entity cypherDetector_tb is
end cypherDetector_tb;
