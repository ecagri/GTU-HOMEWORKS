`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k6gZKFzl8q1Uy223SyN9rdzZxflWKbyd5hyEDHOyP7klg/1IzF5haMqqxhG981bh
47AJWlC+Kynqjyx99GwlbGhBt3WGDkTtbd3Ul3uSIBdDsuouWw2o99H+3z3d//yc
gCjBtbybu316EK/8K2YgNjGYlfdNS81js9Mv7BopG/FFr1Y7vem2BxX1hFKRp/I9
Ve9xb7DIQcvpNPHYcQVj/HTlDdBUgU5n9xJvATLXS0esLRARLgegRDTP/cv5ziKN
jqKH5Jabn1FN0/2WfWD5A4tgm5pIQJ/OMZAax6KDHzQz3wXrE+58gTJ6hjH8sUVN
5kmo+zRj4daZ8zfT9PlKCk5ISS7TSl49TAu1ipwaoI+f4kGlcqdRWQlbUN4RPuNQ
kWf11+ACd7gPbdULS/i2Fyhcsvfn7ZnCbOYv3JlDl2ZYsbnfn/4qPKM+EP38fIth
1+orfXYExajlnr2FmlgcSi1YSzC4RSuHuXo4zB0Fn4monUvCBG7sZEYwcFT7tEBn
`protect END_PROTECTED
