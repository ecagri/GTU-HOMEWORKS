`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9KgXb32sQN4nvDWFn6m3FTYo5ElOOTlUIIe+E9R8Xz+viCsS0Tmi5bpI6zR5U14s
PHIkNrKHGx7qeztAOAZFqCepbaTvopJDKrSt4SXgBiMJMtLJUZfoZD8WkI4/XQmz
20odEbewcF2noB+5CLosdsFoHEkfCUcZx3TiJeNT0q8U3YNAMB/eFE10IM7+Tw6T
zOdqKxXgOtithb9zw8KWpsnwowM5D8Ps2N7/v/DlfIJ9FKG37kayrcdExsEd4ehr
MjVuxXGjaA/Xaqry9AecowCbdTTo+bTEQV/l/tj5b2wq55mjvL2qMeVlfFBhSCsY
8+CqFxkLUu57aRjC5t3f1v/3AYNwgbCkVKM8+TAep2UC+oeWuYSGFa8CKpKyy/iT
AsYd+GGumMZv3J3FR001onAUuCQCpsE40/5exoQyR0Z8j5y7DfWL5i6Rnb2++R33
Y9A7BmR+hpyn8yXQ/8yESHAC6f9+JBQ16KXtqaWNIScIrlt7JK89bhsfqdauirkR
m9cl/7mbU6VY81uCoKGrpZJWFmU7TNXhQWf051liyT5ncnOi0Z1AOyuhaNKzdn+x
DQyYY4eMyOEOmC8TRQag8Tl1W8FhYH5LowLiQ4uN51cnwlbD6I0NbuQM21limvld
CEvyK5fed48V3oCsIgFK+SVt3BaAY52ok+w1hBy2EYC0+LZaMHgbH/zFM/0qkwbU
ZB54niNLHItDOxQ3KJv7PWK803Q7/mwkoTMtYHn7GH8+hHW8MyZRUmRJ4hY7Igs5
kY2IDGmbPN1b017jtUHYoVfYvmlIAXfrH/bZkpxNnZ8FkJPGQlaEV5cMs5w1cMDo
lvwgSc1E+4xY8QNuDD/BVw==
`protect END_PROTECTED
