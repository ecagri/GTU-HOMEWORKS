`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5MIv3EapMC5lv5tQx9VkRmvZ+O40d7zJE/NmSqbWMbXEp6lkVKapuoiE5TN4lv8p
zvW56W8HMtgVIEetzpBRoiZ2vXsZ6Sqm/ys64MavajeWiLVDVFBDGvO4m8v/ZiRL
slH7DmfisZxrZ2sknRxOzGm+TvQ1yxh7au8ZL2JgmbTttcv6nwo3kQ1Z+B8v6pVY
in2vUwIygY03Ekm9JEsqBNoNk60yH1lmr53TpQzF/+Dk4AyWlTT/YUaPBcPxF6aj
0RkANE3xgG73UAbLYAc/6rCAZ8C0VCveqf3T9GWDlF3X2CFxO22CdKGcEkxz8md/
eeOQOsOOIrs8VX6YYvlryi9Z/BT0U4LWqh8VyywCwhtZj8z18BrA+lkHcXuOyKgt
RpGjYHcS14WcxGXK24PtXSoLC47dCo6+wPTM1foGVOA3KGHliHiSwl19Jjs8gUyH
LXNF1KLPU1f/fDSg23MaQruyh/Xh9NSr1X9wczGOXQ0Hr7+Z9Zw+u0ohjjHWPq2o
y5LlvtO7pqx6UYQBxhMhGOewmCZZ3jml8W+dKdKZMG5rNgo4BJkZ+0M2DkpZL+ZX
8DQhANXQHhTSRip5gvHB/w==
`protect END_PROTECTED
