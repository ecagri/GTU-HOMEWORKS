`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GIpQHQT/Etwn8bmwIp6OziE1v+bZAXk/p1EUCMYpjE4IY81iVDSnIBTpeTx3Si6h
m6K6joyR5A+LNqmjWiovPtbWqZRXgSiA8Q8mYAWQuWys98vQW4hbTKjM+cyx2pCz
SRymuWpMogGAmkTuIBcphr0cTiLrfy1bTPdJBEq+AM0EQXmAOu2MyUCENQnBXLki
VKbaDL6Hbp2Uhl1cDIlLk5conuPc3iGoV1XKAc5AunqufvbmcD2eCiOnEBbSsfJ2
fxN+bWP2Yab8Z/9sAF5SSpmjAeOeXG46JglsrJ58WbYZklzoKRj/r7Fi1hdkfDAR
BBvKrZFXUJlAUv3FUC4N5R6Zqg/NgCu6y0MaeiX2WZO+CSCQN2amgdL4o/1aNxeu
`protect END_PROTECTED
