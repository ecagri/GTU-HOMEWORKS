`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k3E5iRVdRdBWYBCkSgeT0RWeOP2gi10ClNcGhtZmzBZ9Rmqpz+o+c8v28OMWwbcJ
eagcKcYx/I7fH8jLsErW/adlES1SDcNGU4XwBQh5WHrJn/egXu0tfKiIu0pGrSSc
ji3lpKV6pnMeEZ+Iy2nI/x4nEORP6RKiINfL0/DW3o13c5ZLloxhzQ8L7AVKZM7a
N0G5wHEJjsf+JhqzIxCXqlvHoPXES2X+iFl6o/HM0PN9FzJ0D95+3aN7p7IIQ8PH
azcwukc9bGKadRX6fYb+lHRq/eR4lQNSNhE5qhyuJIkv1PqxD2IU3lcAZq4o01m2
9EteaH0WvGaXj1aGwKoK1JuW/osOWDWFSUh74lnRenFFcObAolW3DnMqqXhRyxsE
Mcb+yZm1MRt1QzTbQk3bSBj4MxwP7/kDkExMLBzNs9/YPHEzV8oKi97WnDOMQT4s
A50UPdY+D08iBEJJNq2DXGHqxscj+8sZOaXuLAB2TjTCY/ya6alyiLaRDJV5eVJN
JCrmqjGDK+Gy7I/38U0guquxaMSURyyf7NPhJIBOg4CInCRCrcROuYl+bzS0kDvW
8wdlc0Bbhuu1rL5lexTt/tQWZyvvX0+bUDHtQICRGwY5TBiP3g0lAUIiCxeIPkQ6
CzayAH2DSTr+QqqW6eW+7iCjRK5tWmlkREmUeK283sVQ4U7JJ7WfA4wZqYK9FLA6
sMHaEERfTNHumk93kWFkdqqoQfWVC6QYUkq360v6biEUhe2iG3O1SXl1pB6WU+8M
3BKY5XqOpUIR1u9SNlhaD+/nr3Ln11z1Nvd7birh8VJWFLGNzkGJOeK72Tmn56v4
h56iyiYSMPD1/S7PMLSv8mvDw3EoZyXNzoV6PYJFS6hByeeH64EDMpwpts6Mr/Rd
5ZaXlQS2UBRjIYR4maakYvZS2ptmf5QK9DD4Ux83Ef2z3lxME6EDjR9fGAmZpOqc
CxnQBPnxYZhwzTh4OEzlNeqpPrCFxnkrUUcU8YPNBbeBLrNW5Qlmx13TfGHmq+dr
xCK4btk0nOxSd26XhDV+yfupcXqyb4Ho7JsCHTFY18tuNFV3Sgs9DFuMyPR6cyyF
swPJ+L1N6Aj0zQasaAQp0PLyHOWswhBhsovBxkW1ZzEM/amL8nA/PkhPWh+lveFj
gu9K2Ejd/k+6jtBGWvOagiEzOVNuR1dhcqKr3NqoD2/E+ARHxwrQbFHgfr3h4uze
wll4lSugGZDgAq0DUDCPQd4ftF5NeUzxV6ARmFD7LrDf8+y2TpPYIKeLcgwTcS1v
R3FRKW8/F5lj3axyo2ALXw==
`protect END_PROTECTED
