`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5NJ4PHI2eT90d38/GJSPA5fdp4RXITT7ovfk7ceAX+UI8ZeR+3f4veZY9bf6NWXF
Vv4JEpR+GY1u5VzBeocWIMFBuD+yelTykA7lc2Y4mZFQKurzIST1n3aBtUCYrsnf
S63BzE9XXiQzecr50XZY6oyTyV1tDqMZ3vFy9bZuaPJZrXCoIATI7jYZEBszcQUe
QzXEbrb/iTb90B7eGtMf0cL48hzKlza7p4aCqHzW9Jwt3+fmnxnlRJxy2kOpMscu
64Q0s5S/5RADT2jZIUCxBO9dGp54I3LPDEesl801OXZkyESbGKaYjdTdj3iwNhLA
3dMmbepppaGowxyyeiywPeRJd/xIXgXNAS0yeE/V/AHFQ6yVCZrQYtWpF19sgpTP
k4nNryZ61KTkx7o//kmZv09KNEcfTRcGrUrMecRL5yjntCJ5gBCil//YYqPXhvB1
FYc92rf4u5iFcLCot8B6bJxVWDlWaKFtxeYkRPq2rmR+jTB5oDGZglUVfnfBoQrX
ouC/HHhmUasH2pSAcdXJ0g0yic/uRZQStIneXHL2Qvopc0pHjakga6vEcY3yr6Pd
9elhnMD7F5dJ0aF0yZ4NLv/Xy3DMk64uQWzgjJUCFRs6Gy7qAxVcci0tZgzFhcuV
x2ob4KTc+v9PeF/WJNjbf8XPfcx70DTQA4m4wjNAMFWf6PxeLED186+wBDigpNw8
bsOC66FbKSVSaKNsFOD+ehMq3qTqSFbYyZDNcxYtO7p5BzEioHj42IAeRJ6dHgOn
e/JQqliJQlAHgnvvI2hYrOCEnWgYQID+S9XkHDw+K7Zqm5QRZWwzqERXyrQtT0b3
oPZnYRouVVS1+HibYKwDpjuhNCXKGjeQIrXZBG9WqOOekImfqSGgwPnWNBmxLMlP
hx4c5FpFnMI4XsRmwcAmrxeTNYPOowosQDkgpRR24fM/uoaxmuQV5h35nwIGjyMs
elQWX/+1LiKTEhvYoU9eyGYgsHqPkYNTmdkNcqvC5YA/JhKsw7t4LqvC9vQAgprf
PlhOzG75VDEij5rBN+FSDotz1IEAUq+cwj7DhcpAgpQ23JsRGoFd5VPEg4fNQdYw
4t1rRDaApXFZpjMSNl1i/xcKlkKjRygW1rHqkRxGYA4o4N8bGyppAz1Apvbt/95j
Vlp/m90M1eWG8tqIMZFkI8jJjtfMLXOCcEt7vOL+C+h9F3F3vDtrS6yAsW3Ad2cQ
UpH/Bmf50g7NFQV+6IX6xHv2obZ8eJrOy7fgLtfyWVMYxZxwmp/RsTcddVvAH5JH
E/X1Og7U0Vjk9/EecaSOrIFOsX9UejzaRQH+kT57WsA87Dwbc0e3A1nGT73m2rtp
364wF0qoG+EaF5PM4M0fK1mRmWukQOdrwI2rYssC3RalxA5aSLnXE2ka/WurV3iP
8/PnvjOIV9BV0FPyHrftFlgRRVjdf/WBPU8R24WUmBn2op7CiYQuUxHCcVj+PeSt
iktuoFqo1zepCTYPtmHOpwGDU6tTwTYVDvA/GushgLY+y5iHQazR+I6EtAc8pIon
bwXfbR9XABtxuLRbztd+p+VoMwFUojuTeh9Ru4esl632BnCNl4i6c5OrozvD9UUr
K+KPADy961huEE9n1+0yxryNP90rf0b+17dTdr/NWONrpU1msfewdkC41+YHarRr
IQYWCdWpVEqGA+HX5ZyCmWcpJ6rmM7NXQY7tbp/FIBYGf2yzA1xj6u/NlojFJmq6
m1LR5WH8J1E9okJnta/oltqMdBbPuiz/nD5rIz3jtnQMCCUNTrqMCXoj0f9cRflq
/N76uUfX00OMeSSQAcHjAwrD+g5G5jbFy078zkbGu243dIz+U4RZX1uqn5G9P5NO
70vvL/9kaveX1JUJcg15FGFT7hybSxoFfJjfkdm/rZ1hRsekYAbaj+gTou6q6J56
VftTjBJ9GFG4npUCvaD1dhOMEqLxQyKQ0yITxuN3b/XNKB5ZSEvwJ0eUPSuUCzQy
FvtEYpSlJ4lqff6M7sVXzyJvZvYJAZtcQDwlezuVtcY+GaPAFjL6C8ih7mxzhQLh
gaotZuoAj8qTe/OmhGILrPqSt7+Cz67/DHlum3G84cH1Z+rjwGqKnXzFZkryqPuK
Zfb1nSnLNeq1GDd/2GmFhzIQ/gCXGXZUe+XAkQ60B/RimQvU61MDw/ibcMO8iSrO
slUQEhqXRwT1OKArcZVvdjAXJH83Kjoj01nCM+nJcqabZTMmSHpGd/phaeR73P0L
nQA0FsHOeAxHMwVqfXwXEx3eGxkaajsoCv3ZJDgY4IJM6kEFxjWhE44110wWRkRR
ng1OqG2MyTJBswIQ+xKimpzAaTpFoaIpvuLb1UtMBvF6K2KLE0La8+nnuRWrZrU5
`protect END_PROTECTED
