`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hsj1i6JbPHya3whGiREcmYJcYXOkD27TSqQI/0tU4Uhu9JFOTnhei7KLVrhz6Bl1
t7EPcK4LL6wkcvzc0V6V2fkznaxHpASD//Z/BOH7bftcM7zm+uCCg+ZQ5FE5e9qt
OL9AJzHWfH7eDCfSwFPASOq7a4rWQtJNAISt6kOtRPIk5hI7keKbUKqULFRyqt/n
GADepUYRo16dR46b7A//X+HrbbtFL4uXJ8mHUrY7xthztz52DcZnxnRDePx8RCg0
W1T9Dr1jiLaIR0Lsi63fKyZLddTrJrx5ulPgsjyd75dRMeDfEJJlSRc+Juf77nrh
wScFXlOCipqL2UoVJjbJ7pEg8XXt0OFU1jLWPmoyZlThxEKNRCknqcYaVDGcWMHg
6ZQCQrHFHq9kiJCX66vfELTePhhVZ7RlkBs9tJ5eN5RxD/YLxu0Qz76H8kh+jawM
3CPclydR36cQwtc+TdHqRYoZMYshStf9q3jENkenZvbsmGRvdyQeR1mlKvs37+SD
hOJy2YqaCt/GZGTd+PlgYgf9DnS/9qV7Ba/6yMITn7qh+V2REG6dllRiQQl0ofXN
Owid0jKgRZmXdK+lk8NLyzUJx+FxZZD5D+wRXagTCBkjY1mj98U/Q1lGj/R2ehj1
qXntrG9TqTPaQkaWi0X1UPmGHND4Wmz85mzMtDhL5zEzovXZUt10I3H/m3FRh6ux
CHcA/HlbQfQc9JYSIFG5PXWCR00VWtVQyHI1SPi6i2qCJAPEO+giKxBSVxaBtuEB
xd8WLjVrLxdY/zRDF+UaE4fbJEWi6W505bd+cprpkDoNkqZepvgK28D3aCJU8p+W
Oynk3T2ryLG/Ts+SnicCyTHnLlPAOcYlM2N+n81g+Ak=
`protect END_PROTECTED
