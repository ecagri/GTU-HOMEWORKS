`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HQ9wOhZAvDN0hpTnHZvErjEMb0EAEN6U4m0TWlfSHdZdyoq4EKKUUa7ZUMtThfB7
KcNOfgh6gc0BwUY+NuelCUO2h1mtJsUhzqTU/xanqFmzCML1/dpa1sVLWlxGFBIC
rEnP7qizhEMgIP568tLXeH7kar59JwpOa+8fFxyC7a/Qt4kLtFCdC0WmTU2cmkkh
iJCOEz+Oo5Bq/kCnFEif139Awmh/OymDgpAm7ZdGEP2sHWQ8Q7MQX3TDj+V7z0bp
pFsEDKLuzpYkK+LZ+zdUs5vtwGIqovI5Mq2wLB6cMXd7kF+CJzOjivmVz1hQoPu1
Xpjvjx2LV1iQnmodve0YY1BlhAihAQ7lcEyar4l3agO0VpYVSVMy8STYN9zaZhk9
1TY8grSkyXX1BDJfgpH4IQDZgqscxQNDjPMh3SmB/94NNp4/bQiBQbARgox7lMTJ
pGGZIsPtrc/TukpAhVZQ6zsEKGwa+QwxSqg7oL8+d+KRJ7Ej6tK9IFtepKGKHQ0o
QrPBs9wehVt7CcfxAQ9slqKLybPFgjLQ5XjPzt60hOMWIUiyG/VfM0w2MUMjg3Bm
384upnNh0Tc4uxee/UJOVn4O/BnjVSwIFiSkoVNqN3D8YNSVYMIJ2szH5Uj4XQzh
lRK8gYbp/NNNGI6bQTjIZXUZXqumZfo5co/PfViLb5DnGrEfkXolL0G2O4I65QYF
xH5ziztHb5gg7cn5MeMN65UyiDtBa3pYUItMW0YG0YpCiMzV1FXLyFCr+PAxZSPA
rP22rbW+/t7TPav1cKZK/FBPXS057v67QB15JDj1quUJsU7AT7zKnEk3giT1d2F/
wCyyF9+aUq9MhTra8mvgjyddItXiXsfupF6gCSl7FIBglzxtCeO5tLPAYP9b7hqJ
zTWV/4XRebYjmPyFpwxyBIqmT/FpGZ2OHlq6qldN53Gd3SMjFkJGt+4V4HgCbmdD
QnAFpPsFDv+MaWul1BI8kCpsq2FDYfYthax+Hea8ZcFz9hP+in7shYY4yEZHLiVy
LKMwO8EsCNRku9dA7SiPL6XCpik1d4G5v5I3Z9h6ggIaxpN2ZO4ORi1GD8EEWbjY
qD+4sWQIa2dY4+GrYcKne1027Vo5HtXA2Lzeh5JehzuK6K22ll2a/OsShootUgzx
PPTsZgs8J3shD98RDz4zC6OlYbg98jIBEEq5UQtbGcGvNQC7qhVBwN7L04irFRZ6
lSWGet3TQl0+uWDS6gFcKPDPX4msqr8fuTRDkpojbXLVmXGaO99IUOnZ1aZLpRBy
kQA8ZW9n2uivVho8DJma4zIlD2zo4EEkp1uvPpwD7Fy7wJ/j69Rzd5oIV3cdjsAF
yNmZfm890Rik2eKQCszZVl4Rkhi0fFQtGGiHZ+qp5Kf0U0hvXUfgUgLiz8so/pYg
DSZTp7MGrEDRPq3WAKT0XDPD79BxOsA4K1mlj+3LCLx8q0xNEze1dLJPXo5XsGMw
0ZuvQBu7/vRC+0OBuvmeWw==
`protect END_PROTECTED
