`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
240xPRa/IlJGA/iS2uyGVlvTZCMIrI2j8+vVzqC2qn45C6aFL2JqsCoX78XdNzJU
o6VhDK/wON43OaAqkVAt7u6HxCCd+ds5eUMpByGYvvRn1mOmIh6WutSWgej7Svd3
b1f948SW75/upegTtA2OU0R8Q3MJKrDptDw9CYTxXVBfUug1J/aNSwP+RGNx9rxt
6XNTjNsIGc7SqTvpedSuA9mgGM2Pny5Qo57A7Lo5ChogcEB0+flv/V73KmOWt7SY
z2+Wh0QCixg89icZ/ikLPrwzqaCqeDtMUT4B8tgmbiGUiQB1JuE4TQ+T6yB7pXNz
5nOdJFyQicEAQwVWchJt4Y39bJok+c+mrbXW9TnapMukO8FL//4kQNuC6dsy7lry
O+fbMfttA0bkvYkmR8L6G+xXGJHAlgxg4p/retjdZ9q0iDgYPCuPTs2BnrABd446
m0nIryiXliIVwKC60I0zkt7/itOiqSP6HG20rYGP7174ahlqttxZb4ZiQOp/5wnm
wMwPiKTkbvBhGNfzEfjbP6uCCirccr3Zc0ANGelOTG5XDfWaBq0LvFtDTxIwP3Eh
uL+zbZttBEs4HxtqZMRzJ73ppRMilJN9jS0hGk+gAYk+Ceu2v+uKmuMCe+OPgSBO
UT+l6l9grUFMFp5bH2dnCjGS4cyLvyuUSdEjAxhlgWDsLYRDiudf893cX/SC99zC
tuW0Bu6F71c+07OEcAh2Vyen1cUfm+W6rq2pm5H4O0A=
`protect END_PROTECTED
