`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LBG1udEUR5lP4I6ZLRuqjRNZS+Cr69wP3EtB7odIqoiXBwnwa2qYfTSgV9ZHjyvd
y09Wnfkg1Dw9nZgvTgbF2uhaIFMRacdxcG/IwpqFFOCt5ZenGjBg6grWrjvt57d3
3MzxbZz9phYfYA7RJxrCoPEiGk4HNG9TABRoDV/rGUyxfJBCikxDszsa9dQXghOy
Afv8jcuutnPgqB+RjCq0pB1vJakZ5nbpNNlYVZtI1wNk6NA8bAZt4Wmc4bjazj1A
qTdYrOw031/xFCab1Jo/FejNjsQOfBofJRR38770rB8YBtiGnbEsMI3RX0HiLROY
zXnlftEtl91TR8MoirOgvQEHJ8FPy1fXHixGoVW8QlXv2PuKN7DonY5jmKvePDyr
E5yz3JjW0YfdKO3h/D5jcmdUgTY3bF4tUHE6jw+RGPxfblnvPGKg/fLV1TMPgpBa
SX3QKg9KoLjED6ZFRO/j8WKxf9kfMp0nwU+rqcWr4VRbcUepRYfgPaQjjhKoHIFk
T00BT9YHTYOvW6mxLhO02398ertTnlnPasX1WNlptcSCH1SoLvHe6SREqzsg5mSU
eyp++vQ17DbJInaGqJxDreqIr45ySGMG9fg1hKKP44B8ZU0RGPwvtTco3o0HCux6
pLa1UZXTRpGrWnxnI2RjwJqjJluAhcVcP2NZq3OWANitJeUrwrP4+q657qdbXf+n
yJkiNAKi8u3XRJf9b5vuPA6qosCOyHOA5PFF/Ri0nX3j+J9ewGH+kRNbzghJuaaL
H/+PX2mayG4jddq1sqGI0bqVh5OMLE1tegcsPdRyZZLh+AymQeYRDezgI6YogkCZ
9lmY54joCIYqPzNB3tCXAGR3g0KY/izUHah6/cZWrSspmDy3SjzYM8ismmimom8O
`protect END_PROTECTED
