`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
38R3aVucfEIZMky7rS2Vq022sXxxyCXmq6/d3Qgd1GW7G/xBdtb8KMNaQ1YvxaqA
6A06yqL4W89LGOPXH7cfw2MEr6VxeMG5cjwsRdbqUV00Gg8UqB9hGJK83c8IIV26
KLImEtZ7EHThFmXmmPJyL+Q8IYwqzJHCfNIdIO3l3a2xBacaulQGOXnrDnqvELH5
X/50rzahHkUfO7psi44wuR/zi2UEphqzOfXkwqhm18ceZE6yhLth+YRXdK/qNg0A
XmmjfO2YBtDpggH0kyxNr0NzeG8Gfity4kPxo5UIydnFMotUKj5SfGxu/xu6UsZl
eqMXFG3bo/RjZ9UnALcaIc5ix+T2/4Z+FR/npSqn1Crj6caLbzoXaJDaVNgv1IXZ
kK7X/kwXfmKUqK1MR/ia8zyBqhvSxaNSUw29rhVkooTPhEMAu6k9AlZ10B4egw+8
aZjiQSFPPB+f0ORoYjDIIqMmpo9zO6KXAexLWTeJG7v83a0/jyY7wQLbNkEKSb/I
yztUcSUbG3K7XE9W3u9RgRKFhw1fGZWtNVwJOCZWycw6i4qnOWMp7Gp4GjqIkN7i
6fgP+fD6HBUgTk2S7ayoNSs8L6rsUkvkT1Vxu2VJXB6oSM+0bgE/SFHBVEgEaq3+
Vxt7WmNYBOVbcZVTgB6sRRYZoX/+qsUJs+ehAHcB0Di+ZGKA2ZaqwOVZxThIV44m
IPcGge5fbw3+pGxjmIpFcPhYHOi07gclnvpc5akrVHXkolh8Czjke7TyNte9YvWv
CbxKWql4bHWGht/dx0DLwh8rjr/Er2Y739H81N6difHI+HMwxETHfvKydtjh+RfE
otw+5V5CcLr681pahR+rpHiDGIVaAJU6dUc3EdkarVPaT8qr0zSiprewBnBoKvjR
Gs/4Mn41EO+M27jUJMgacBwNJdl8WLRGMog/0Y9qHC1XidB2eIa2yw8j3RLvX/ib
oHl5eJF+uBeLrEJWffuPWP8iQzDbtPLS0ZcdiYtvIr14VXvAZ/pVnaGV/RGvemvB
rsF7I9MheX46ZhYYeRnkfvZqWXaGoX1ZESTaUHZghbb/0Yd3vt1cay4X1HniJFkl
W2/w6nXdrk3CB1vmo4G+JLYTn98/jwW0mIYUm6v1998OxqcJs2tbmlo/TSUo+zhQ
yEjSIwZzDwH33Mwgzxm3XZyWjyG2OUtLUT3tup9v2yW7yStwohJqwpu7HwdSHv9y
LxML6419rH2iMHQ76dhUSGAxCNnPGVvyvK1+G9XpnT+QO2KSkEbZiJicjSp+CM4m
l4o+cqxM2sdM3gH64qrw/4fo7qdP9cth9dK2FOqUOW8TBskBu4tYJ9fwtaFExfR7
3/vhCyqD9fMH+hojGGaAX9BUueH8+tWNHSH3gwupu0693379HXRzTPTltTDkAdXc
wTVH8gMUEm5PzXRiPZHuqowKItaoGIELSri8a5ALir3zj2VoBfpiaNpxxRdAFV53
Szxhd1qbP5FgVPgJ/vyxKWnsLtGMSkTa7IDEGAml7ISWaajdw0CELVsjMuN8WYZK
iBcvAL7hDcGlNj3a+ZmiCsA5J2Y3UxCh/f/ip1scRdxf7iy0XSoYycVWml37XWbf
Nfz16PlTCpxAgH4mI+v5q+xFfCSouQFyICLRK5jXphfiMKL9C5ixc1riKeY0eCgF
AzHxBY9S/hJrpPWWcToQ6Hyx9Stog0PaUDrtIIFpC8oXJ+1YPzWtHJFMn9ocbFAt
aBXVrO/ce48RY8wDQ+X+zIlQHy+DLotUSePSJnn8wgdabOk0gLR/42KKG+A5CV9k
XMklmqQPxQfD3T5X+T997ru0wTeTgZL8+iuC47VvkNGjqbEj+fzLMbO9JK9UTJ+L
EWGfE+Xn74NLLuiLFI9e1ZyUFCnAOndL1yBHUnnStdUwFa6e0thSNXqeWalBShTZ
TyfCxPTqhBdvEsdcCO59NKjjhBmpfc2rXerQsN++KWMCiy4sdDc7UNMKttK54fVZ
0AKQ1yiiLhdwnOAwQoYqX3GyPeS1vRRELas+y7GnlKjQ3Q1HjkROA+m0v/CFyYbj
1MK+9xODQO5tpzOSfmWIPaOmjyGrEQKtTrakFDkFQlwg4Crwy9GjAZy7QoqgNKvo
kXPhNA34We8+0/tFJnafzL0H7VXNeW4vP0sWq9AsYSHz9M5INYESTgLHWwNLXcyy
faCL5eLDIRPkx6iVYgKXQtH3GcNnEWz5BwByoF3AH8ZhbKHKF6qbV9597r1qtH4U
68hXlHOdGESRJLXpIydrsBOS6CpMebpfkPPtCCQZE8h4SzOTjJuQEZB9/CzPj6NF
ee+SgqH5V/xBt0NpbsFkft1OEt1fKpa49r3eF0qh7lRXug6V6lo65lazka95H5M7
GQwTKnuf6rk7R+NepxkSnimQsDlLVB0o9CTLwi5KHypHikq51UxHM21Z14LVwSgF
BSRY5uNrZMwUzXDy5PZwy5rQNDepQ1Go2YjVAgIwkr3f8LjzeqehE/8KTTgzVVpS
d3xCnK6CUualbkUvawiaZ6ELjQDZ6H2mBB77yK0MTUAHi0TCVTnVha5qTpVySgqu
aNz3F5m8jMdna6Swre2yF2kbo46iWQK0euVAKS4XYoyd+7Z188npwXLRc8OfzvcN
vNKzGqIzdRGxzMxO72yz290JfYaU+jl/dbAu9ue89YGbCvqhkCE4VwFCreiLyprH
LWxiwb8hUKZRRU8NZuTejXRn5GHAECIh4wds1iiZyAqsHs55/cSVlV6PpY454USq
3yOOO+2HTDrAu6UahjQqeEC1fa/4Y5xiz9GE+BYo8RItEb58o/2QEV/k8iUBKVHm
GiKar9tCYUe809y/bk1WP7VkMJi9XMEkyBxzMnDiYVqOtH/LeYom3f/f0T0r2a91
FznzStyDCBDpvluUkh60q/tCZusl1ff802918sKhtZTqzELW+jLnIJQDNqlPPEsw
JUlRz9/K6OYthZt4DcGgzZNXMkl3WdtmHq1xXLH8+Os8WfL2iPePx77S194pkQeG
GzV4OE2cYyM8BN3Tyd4+yBlsVTMDNWrsvZ6bgwcWtN+OJeycsocR5vZXYK5WSzA8
vLIfCmee8Nwv7yomNME27/RDdTmd0uEQX40vXknFtn5v1vBItUlesPeVVbkPvyE/
LL7vLK7ET4J2b+di5EKgzAfbpWB176ND5QSM5eVSK7oOuQnJUzArpoI8761P7TIX
ilRIWBAQN/D+RUC46QOW/LUreLzbtaqIhq7owkW4bFy0urN7/Iv1R7UT8bemDgqI
Yy0s8W2Ap3609Mri/xDxb1pL7LYD0p0I72x+yNOD76MxrI8n579hdf3F7HQXaMur
TKSR/mSOfFHa3OluZHH8yg==
`protect END_PROTECTED
