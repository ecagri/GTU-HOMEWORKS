`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3/R35+p9ny6w7+DlK7QSQ9gHiOo+FMIJ58nXiMvDx6r+sC9PyzHJvZfjRLb2YsEp
P3h4TRt5DtwZgdMw/TPmR1rmbLx6HhfD3teh6PLQ+9DDoQzJ/rzJ5Fwev/F1vrmK
I+bn2uHstQtfOJvqsJm85R/cYHmU/uSPq6FRuJGZ4ZRo6mP4/zvoRsUyvx/wHF9M
vqhwt0m/v2iHCeciCJ513+TI5LfXntFycYQmgYYp4Yq6tVia8dnbvtMR6RjiNVLY
/BvzyNaVp5VjWfQY5V4n/plRQIpvDRM24LEK/GESLWoKh/bB8Pl7zpm0qWB4X7Kr
VTxp5jCo6bRGVHPTWeBVKAFbUm48wPiVi2Weq3zvSoAbkK7lVf74wvyvB/537PeF
UUcf+BOqMWC0X5as7QEyl/hPkjbI+xrwoSk7ZoCIwC6OHExjEXGkYbzNg4wbxnrW
IeJKbzjDpP4lRpFt0csixD9T56oU8IRYnbwD+ANhNI+Xdi9OdfmbPiDUmEZ411DR
eQrIsnXO4jLo1mKTqxI1bDGoJaE5Q/seWGdyHc6Ns4jvxiV8NE7lobcr7afZQvhU
fYTabV7ieJNpKkNwUenNHCaXdmwYoR9IlX8n/Ky8ptje5c/jNuUNGBFaRdICsv5F
2EwDrN3bpZ54oD3vvlc3pb8AzHxMXudFAHeOT/MIdWUYKmbpFpb967SkcPBRXQ1T
E0eW8+otmtX11WCQnTV3NxzaM8ImY7fVsF2RHpOe/7acvk+n2rxD9qYga4a8Yz+T
rlYBqLQgpp88oyMr/k7H0LtNneOWfkfChCE3VZBlU3SQgtN9OnYssTLfbrc5NZQo
pr3TLlYMNJi4vueYgYd7cU213iL+fg1zYFHukfcVrdEnjTYP0opa/5OGMH+TQYab
2twabsvTirFWNUn6Xq8Af3YW26DsBuzkX9mLi7ixGNhS10XRyj7HFv0x7ELb9Xb0
db6avwb/OTZ0xBsv6ymXULHpIyUO9qkqVFqfRhPcfYzF0BLz8g1/u3M7j7z5BAys
jKPRBsPHEUkV8LKe/3xPhgiTGPU5+mYu62otiUdS3cmL3PPPcJs6CCeVYYp18FbC
AsnOE91pWLqwuMI+3spK8JpCSQZp8u/Q2D+o0nZr9niGiXH/iQ29fg1UGSQa8TbY
gRfWKQGXktud8TCG8MM2P3YrQVWUJrRBMKQXDMhhx0dGmmRq21smmdJbmC/YlFYC
QQAsEeb3xZ9ea6AovtSM0OT5PfiVBkyVNU2QeQyUD0OpAOZWyX4KL6rS/4nF2HD0
cyngydTlpzUUvaFoLuo9hkpUSxsgvF8Ys8cYh/BjR2HhN251sgcX6/oicQFrxN0C
R7AFzZxdSOJipcbss02hYW/G+FK/pNtYZK72G4CqQq4hwf0iEsQ70HkMKMcaCion
/CkiAGckPoRlMEwqrqdu0BSdz0wKnG15C2p3NP7Uy+NALxGBqv+ak4WuioAnFh/z
`protect END_PROTECTED
