`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fX8pnwv1Towx3pZMbUyLwwVwGPhqpsd3xTcoOCe2BruRlRmaeoeuZikH9sIGhfVh
aQOomqyABtOAzj1JFAQ+CzW5N1t4bLPOIQCR0iVd8l7QxDIH3VxyjxO7J7LhgIes
vwnnZzSPdJFEPcQxL8qfPF8DzQ1G9X8tIRCzhIOvriXzwVFBQM2nD5uWgOJwwt1Z
Oh+SeZv3yFgA4uKYwPsnFUQwG+1adSy0tsRPjUraWNU1pOfWpbMLymnueVdFCxpM
LXEqeXjw7c24Gz0ylsCFKghyqT8d+Sk0asPpB6N4scCzm1orCouwBl2URg92Oa3p
YibyF5K4LJ0sWzEEHtYDPfVoej5aX/ok9pIDxhTm3LNPpWw8Ps8+suh6STn/6Rbu
aW8ibXeV9K5nGEF5BKhikwSEpYT2AD/pjmoFVnU053pTB22FpYz9vXKg86ZsHn4A
LmizKNtWlDhwuQhMg/RUjAw8Xs9RsYsqpuLtCYZ6635OYelmr94CPuurxdxWvrki
42mRTriBpEwjMzUM5XgDvz+sVQG7fg/w5hZS8+WovoOIQX6+gnNrgxjA2hNVgyxP
YYs2OX9t4YqVgbNOfT5epLfN1xtpNfkTFROt7B/cqu/jB2aLfK1u8VxKpX3g7bZL
LkILvle6MSLpUYO7kKd8h11lAQZ+9kysejc+nQje4K1Od3TgRht8hC8+UPc3oZ2h
jbmrU13PvwJNJykk8LEMbdYraOElk08bqETxM4Li+/cRpmHOZHGVVq7A4+VkBtY3
mN55pifJIBSfeLZ1getQcMk2waYPhAKp5fD6Q48QtebnkiFc2tsIN2orRQxEE74e
6QohEx0nXfUlvPEv+u+gWGuOvOgqZzwpO3huzdpIPwzXWnKejjPoYrv0yp4xgRqo
OeXpVrFQRqBl1va2g8FL0/+sSlV55XA73+k88Z6jOVFkHGt/9CP9yRdK1X6FEVD/
C/syvMxgjRtntFJEQZOMQUEbFydQRF8XD3/fohYWLXs0EHyleGbXg+c76CdIo8Fs
50KxCwPr+GqNFVKOzARRDHzOo6I2DW5TNfhAa/pdv/ATGWOsSYEfo5nFItNRFkip
Lb4OTCu/hiIoQsQWw1PHovhNOlW8wpA/tWOr4TgDCrKFPMTDU22FcucWUglrjBeZ
FbwHWkKeo/3F/XZ6TlucLLr1mTxR3ljVQ1IBDZFJi34pFYEfiarq6FM3z86z4Tvv
nm8vCIbnO8SqZd8NhVvKYz2PdcV2gdXK+s4fQ76B0b6DmyUQnEHWWEve73S+6L81
QE7afFvH/ebCbqNhF7Z3/XG42u8kyg7KL4deRNxl2d2QMVKUf6ozl9JM+0FB/Wqu
3V1Nt6ZiB6na04wlrppnmI8yRwWL0ICsCEcjFGMTkzM9Kj7pEG+qfK5Yb430khho
oWsBiUFqYACMhSuRSom769DeRroPfp92un6+QUEFPqPz106MHt145wtz79beISiA
nkIjIZuFRx6d24N4Dcp50GAFs19MjlA/NxRuDyOGWJkJf9uf0+NQvnnIdgCyrdxI
Y+/9NpWmT+RTtO2Y3Z7i1w8OzGPsgYleT9xC0uP6HZuzPVJQaz0wNxPO2zFIC2Ok
8vy++OAOkT0R0iKueSoXdsbJD3Df4F5p5+lwOZL59jtC4rxVaHgDRzX079kdLcWu
tsqv8CR6x3FjBr3MIYeKNJAT5MMzeU+C1WRHnasjA8+a8GIaAF88ha6yfCS2Q2Hq
61HgiwPNvXX2bvEbfBq8sXW8dr3zWDC1inuNxnlNmr4V9AhQXDqcZPJF7jJgQdh4
NtdPyrk93dOQe++tfWKRBXhVZVKBeXo4jp4zXlG2AoH+0PUUWeQqj7u7iZwYjnw7
V0vKZsZU7efp0tx+BcRtIdFf9ag61pbm8sOM1IysuiDPNpK5AN5FeHUVp7uOdxAl
HdjKARc2VEY7pOFDrfuZLMKZhigre+igCuujWciZaAmP+G7rqWPYc1Z0HO9GG+3q
8/G+Ns7SBStq3B7ZLjM2CTxYA5WujhYe6wk4tRuxveLB32TAqH3pZEW1S3BUB1NE
LSILe+EL0BfTEzKwFiXa7oph4QYcCJGDzz9r2mPvwNgjV+P8TVJaG4YE7WvcAY+5
114FOou6QUlMdjR73WJ84w97x2e8pIaIwRoXgnqOM1AJWO1K/lsCIT03MXPI1mJm
NXW4E6/f/DGOrwZ521CKsitwKfiir/N8fHwf19I5Q2Fbx3kG/YZDpv3GAtqa22Rp
O0Z7AYRHY0daAetnYH1uMA+1+hZ7RxyPC/Da9WWVtq3z9xJ6WGw45oE34jQBMjYV
BxE6Ws0GrMf38NBSii/75VCFMvSJ2ismAYisXVOO+PM4souAHWNSeomPNLf7+asX
hvyVu5akP8/YRUoWIlm9g6DSa1gFzoAHnts95tPnFSncRyyC567+Blo8EfhFnkGi
omUCY9+CBmV7cdF3rMi65zXWdrTQBriC/Jbp/LnUjeeDtMQlYD8hFvm8w23UszSv
Kd2oUZ7Ym1B6TbS/seGUvfELtnuqBiMahANogNMhaZJg/S1FSpSuN8MCQLs3AJn4
SyYURTcME8i6uVBTwjAB5dxUYeg64ih7o8wD6dG8/ELdKLq91Cz2sW09IG8XiPoH
y+0jW6ooxODg08hv+kx3hM3n/r6CJmteDBMaqSnUC3Lx0VdYhRFYL9dBEKLOycmp
Gbjs8vGxnuEHs+IvpmasW0HK4moCIz4D9XtAG4U5LwapxJSJDwsfojjFGI+V+ffw
2CTx56Cab2hE0zckYFN7d0xX2NaKg7tDZkb6ypdUcvg4Skz4uzsAV+PedWLDePi4
qYpRDuKMTFF/6KPo4FtZ6xbKM/Im38tdbEP2EwjNIPglT10AK/I+FvFe71Zipsk+
S0WbsffNFop1wCUXg19UsN60SDYQwIaYnGhl3XNwZnayW3miJUnbvnW2HI2arPj5
i/xhCSsCNi2rCnzQ73QT5wEdf+Yuf8vIaPSMmqvyPjc0BDW6olFHpjPOZbeohUPj
tDyBvGys0K97i+BZoDvp4eGbJy+6ie6IIviiF4kL2rfbaKTvrgsinIMn/uvWxpnP
8neHxo5+qs9gmY94vqcXtHGw1osM3fHwJI174NOxtW5tJ7KBVoe1ubQf/nxABl9Z
3Uk0/zU1SOgWh1oz2I3uTPiFwWpiHUT0OTkbcYa4GczYB66cFPkzhSUH79XVGCjM
nhqDpTstmIJXTvUgLfFMfeYqq6fEA1gCEHJX2WblIbzjgXWvwGObWCIYzOx8QwaQ
brRGWKGx4YGrrvA14vY0k/WV4/oyUg23EDsUv5Ir1zA4TIUjae+7bm6homml3vxy
OxQ2LEZH6Ric4SqrHIIomZregXI/snT2apK5KLEPeXmdoG/FcReRDUztqd3zULkD
J7CL0YxDY9l4A7P4huLUbA6SBmnaHggHYP1Dwqg3uq6JJsWaokol45z7TmGnvwrz
/mC+8yiM1q5O35Oc5XV2beqfyPu8rPsK0n5Ai4nuCVFasQSZL7q+DtUR0SoQl6iZ
owWfFmzixAxWZBkCTu3cYnGd3VnTOP4kA9/fp6UbUdDsdXaCeJOAa254LchnyRZ/
N3zvVQtuTiI4d2PHSdf6Awr+1Vba41USWKQC7rAhijnqprieZ6tXGK1C9584I3rR
zQAgEbc7F8MVP7WDEZXPC+FvegNsIPSC/y2s/mIjDRkkAtI/7WN63mLLnEaRh+M7
uRq1q/ipEBvsHCn7Cty1cMDsOYqOMBiBcTi6MfK1InsIyWvimTy4H4AJUsOGgdIn
vfK8s1oiYIDQKUpXGcF8HZBItaMhCUfOPLRxkeJkoCXoApKDvK7Aa7fuF8QHjqSB
4LQxqIuG5pmTEP50OeEBvPcIhadGOiT0pPqn8UTgSenXadzRw4wC3CUpB1kppr2z
69mhcBajip4J4FOscDmA/bFTlxT4MZfTSvohiAG3oNEPqzAARgot2jQf1MGN3aH8
L86qhGPkn0j5cEHBA20VxJ5sqfrZu2j2DxxpqhDCdzIy+87pvFi/Q9eMw7KLtZuQ
I3WYBSL24BUmIdE/yJ6cDMfCMfxz64AF7IT7vwhDg6Z47KC4j9SFW55Ce8erBu3K
`protect END_PROTECTED
