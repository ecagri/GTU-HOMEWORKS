`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EymD9vlM/8iBAbFHlvlRgJLAGwxl+s3ZQ3jyv3hnbkFc5/67g6hRcwUxktCd6pvS
JkV9LMv5J5KSuihBjugKLsGDiZZmAaCxDLZwJhXWz1LsWUTZmWlgHIZlD2tmaMvS
mnhxZrtlATRKfVgvS/SLZEv8q+djS+GDVpHyrM6Pe24VilYgG18TWJbKe8ZUKYmt
zyTdPz3dJGv5EptjhUlSWV3KoclZJijHOTLXBvWPby/VNAb8ee9BMugb1v4bHFEX
mRH6eHNY6keMzNabRWCkeMbRwaN1YKZVShvieqiPZ4cXCa6qWjwGx3i6r8diRlXG
NcjSDIJALg9wBEriR7c9k46x4DBoLDIL6hws+FT34LvkEe2CU7YLuojmhop6pJGU
egjjifF9EthZ6A7DmOOhJM7qh6McgijfR4e9PMIVz8NpA3+C9Y1ciLxOPnexYbIp
qui3bDFV82nvGVwJsRUGQsnkvNsrzPA85wYExo+BW98ujXRiTyt/4fRxAt0R+pLu
laKvc7Fvwx0TkGS6WznB7Rem/Qhz3Yc8h8ylC0M5yJCQlNIq6jGyIMmusHWXvVLK
k0KorRWWOXKGJ/DZz1al8PH3pbvVDzbux2iVdpVLShaAH1XhPlXS/xrBCxXtncrZ
6drI5/PU31KY+oI1ZXY/zgJBJVWQDJrZRkciDHctmQJbJrpRbZD/agzPd/+zDI4r
SrLYA0hT9cVldJN42EzADMNFDGXjtgGjQrxMHJ7r6va8I53TlNKQC1V39eei3wyI
pioO6xEY2S0Q8Ca721nsLPAQkbs/2f1muLBvOAg/cZyW+7JmnfkqV0JvEU0TJgHA
GnWYs3WT7jrb7jakj4V/7EUGJ54dGsK9NX678EsF96MTBjFLuk9/qTsQOhg94rsf
YnSGdq6s1x68hDgBWO4nsoA8G8OevsXWDzG7mRNGJBoNxzKKSh7WtjwP+o/Laz+a
X3rrWQ4Bc699Dy7OSql4/CmZ7wHmXiUVvUCEPjB0RiggFjyegmomFSMLp/nqn/vC
CBpdyrF+0TO8UC6jtJhpu4jig62zqcDNPQIzL/PLuWn9Xu4YbU37Qoc9sBtQ4ZmK
sbA0qE4kWs1+5s0VxT1StTww6vfacYWLTgP8yVIfYMZgycwg/dyxgarKsUN3vaoM
NXFSXffbphJwFhbyJl7LMhJXV5OBlAq8nBdzPhaJIYAaxGChmvk5B7hYJi89fg2Z
rwSH+S6ioa0sYSRKEzJbkGHq5rrp8VUPMJu+ggN1SU0hUnop9aB4YBQenaDD0556
+HPKYWNeE6WcJ2cvQQ6hnCJY0d6nTm49yHl4A4vqoCoHqm3+sje13bMPwGm2T0JT
gouJtCg3jBBLI2PsMTe3ryahG4z1wbd8IvfaBHYK+qIhideC+ddPoytyB511pWj0
MmnhBzD2NnCXsRXrfzLuR0scIBw+WF0E4wM2aTt/3AKZNs+U2DwBNYCaOc/+sXbn
tX6YxJf0Gnq3Pp0GzHrW1Xraz2v10dev9tJluDKRIkNPurqUk7V6sIqOwa4M0673
JcByircIkOQPuGW/9g+UtRDJ4lT6A0t2rpZdbxIxko5d+XDDbpEd79Y/0ie/iZZB
WU95J5lLdOx6GGsyzoWNSyht+D9HRT6/eVQqXcym6fwnMjNX7pJCU5VVJjGT18XX
yRhdqIbMFnynKai9s9hI0LZvO9QBmtmU7faCjKTHsnFciNIS/aZionljpsK0ydy4
gOV8fKr23a56ARMbpX/zcwpICOCnIxTcu3WixMMNy+Vqjj07W+MFDh0fvZseesl1
eFtaGIUY7fqzqykOlrDlerQDv90zlItHQMDaJ765gMpd7/LgRpHtmXoOF/bmn8QB
gHfrxXYNt7NJfTF87afHrdAGr81evVpXzvu1sS4KJhmIRIBsCZIGCrBmIeCOrDTJ
KIe0ddMJfAOoqMQedNWRzwhXG3LZhJX4r2/EZUiCo2P/pEZ9TEdAHDFi7yqrCT5k
VEDanfi9h7Fb74DWcorikTVg5tRA3atLD/YxBNwHphJ24f1hxKHfsU1AQKOJMH99
TeOImXopxgDeOj+ZDNATJ0OPlHoRdF5GhjJ9HQF6SNTd4plqs64ieeS8vmD6PI1B
xcFkS5hxhXq69Y+dqlRBUelBYuLPlbqF7NQVa+GzzrKLcqw8kOxiVh/XCSm5sGsj
N/jp+zsoO30hJiYnfkid47Bs9fQhYR3FUSRUfQf6/9tndBy+ZxnuPm2F09VXHGTU
ExvGJYGTIDC0Y13FqeZBHNBX8KqgwvVOnOA1MAl1SGoXdTJJcwt3WKQnA81iNVoq
VCeVK4Eq3aBou3KW4FbynSRDf9ebSeAehJEeWJP/szgnyKNUGeKIi3mRGkrFO3u4
RQ9+jCJMxtKVldiNlyd9P6VoqgluIZeOCenbmyafrPG0JYTcEBbJWqsM+68AZ5jK
F823Z+gEiRCW77IuuosQxKZYER6P90Eo4RUDTXGM6PK1yupsVDoeZh4Cc8hkW7s1
MbnlNHDHGeNkEG1+6MVFtaFepyDrJczaSxtPxsQpaGMvwumUKhtDXkVSt2E758Uh
GEQOsOeFCxtgWuzZpKHNhA6I0qWvgoLIbIxOBcx6OWhb0i0yfXoACQjmyKMmhYPK
QtJZ5pN9ieKGz13ftiproy2RX2MVKcfLwOvEPGIrmfASKu8dOgr6wm6ZVzm4i1yS
+SlRhjxJ9coRQ4/E2DCf3n3/oaTFNeN7XbK8MUAeVseBhkp5dtglu54hWPl4FZ6D
+BxRYBrpiKl9qfR86DuFEyMzph0Y+032Wd79ZUFpMjJU40L4Cwat8C5+EsDUrxXs
3e9DxToYjfnxUzEFhPxhCqiwfCfJMPDRz9R+9YmIg9qyinxjzTfrrowTOry6Uwca
WbRl36ZNSIrEN7CP1wah3gFc/NtPDPzuTD5s4VO0vd/8vZd0Va5zJTdT8GSx0qdd
nJSmrTQ5ruL3VfmLbY0gtj8Py4iWMQDptES+/pLmFsVQcO+hftpnjE0tMwJYL7hb
KTE2yWygEocTUWBdiiCljQO0BnD1rCQ49IigEN4WHiwIfBLlD8r6IY+LY/XsV+1x
h6xX9oAXs7g/bFoBcDSEK9d3dVii8cymUragG7t1fu62DYiVvArU2mLLZ81hTJyy
FxHph/7iNL+uoCQ6hUPqxya6B3eckAwZ2evwnJV4DuYCZfMZXo4uP7O9+9i7BYuY
Jhv8BE54WWXAlzfVYKlHUPOAAkK8pzpY3Gm/G421eDpNIIcBznLReqrMG88WvYk2
PYlLZIDK6fHBVIG9BrmHYTCDlPy4P4y1w0bcsnRgWk6z7Z14kRqMrmyNIxOekJSo
yoMPOfvhfAqbrC1ES1/D6IQ3CnWyRHKmbGU1m95tOQ6y1X5CuwzLNYFf1FvHRAbT
/q4YSKXhd1boiIYFutd4Yg3ns/y1D7CQ7aIbAz+ckmoIm0syPciVnDwft/2Nd1Ky
Tu0nxAmQhJrHAJ9K1i8Vj9HAIHOo2b/DChZ8Je7VohiO67LdhjYZJ2N6ZJsrePo4
FiZNskv2O7N4H6FXXUmLY9KwO7nEy1qL5tqmzyjSii8T4EogyZaEksYO5cU+Gkhn
PxLfRur5fABLCMoav9Cx9CRHwvgOzv/13d+bWGPM8WslIsbFPZvgag/0Ycc2zPH+
dO88icd0NpY+jQkdoS5s9jzu4kNUzeOMTxoo78DwR+JWr0h/6vZqxsBTEBv7FQnw
ug8yNT+XqedzuHr46kUv1FHLYhCGA56q6hBZgNoinv9r+9jBgtAvcfJ1uXWJA+o2
XNPthQr+U8rWB3YVvmBTw3mG6N7tKzghtLNPiGFGcjxrwGMIpqNHN/wWX0d1tIj4
MxX89X3lpCcoEd/9LS67R0DBMt0jX4zLr1xqN74O2xcdvxGyUi6da7hU1IoFKJAG
uuPLpKX1B8J5WEpENPGzcgzilsh0p4vfn2ycOduroYrpzT1NvE3kEnXZX6xLfO9q
9QLUCkKbIwiD1/2qLlp3B5U9M4xFnewW4zWMehqRAa6vYNpPovyR0SUpMvNpHt/Y
BcksQYF0VotL3bArz9Sl50KfXdUbOvi5CNy2HuqJl4I++5DjMUZctM5NLhtflzlz
/HnGwVRWbFiu6E7rGV9Sx2dU4hSxWEHMcOU36Z60vJ528egf3jSDIV3vs30SNDYu
`protect END_PROTECTED
