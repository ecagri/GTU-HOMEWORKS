`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LrzvQKwASe/ba4CcIsaAiikmQUexSMsueUMliWRo6YWJ3BBx2LOwMIYFz52MPF6e
56KRLMX7/n2AmcRNa2gqDD/w4XDG9s9xm6O2P/JzGix+4Vjr8gruFH+3iNq8WQkS
t8cdCVzXXGScgC98g7mr9kYDJ/xkzxNkLs6dENBzGHnHs0JRT8Mkvuy7OF+KyyFn
Q1QWxzxSyMisCk2Fb6wcN4yzprvNrKRqsEhr/sGDo2Xu44WUoiQgGBea44+jxbwv
QqKHGhrDq/KT/NOaHQtXO4CM9Bzt6Ku6ZFKfgLvp8+Xzx9eEWZj1L5CSNtr14FZr
FayIBg3sbDtldvhe+dZy5azjO/CN/aOgc9QWcTaqjLBPmIzahDOhYBjsr6pLLBLI
EIV/vcvbke5gNDJLsVdAo4pHfF203cAD/f7heC9YESb9c/9OYZTr9RXP2Ym8K7Ql
aMGjHuR5Ep4nHP7jhS8EzHrirnOh+c8TgiBdZtLp4h7VBhmltf1tMwuSqmgXAhJV
Xl0fEUprfnC1LqYF3z5VNbzLO/WVG1luweh2sRA4RAGGpRxU3l8oscb5QA/K6tkP
6JafBgJI3fSfeAJp1C5Y5HFfSxHSmQvDyuDqDCsmsO8GNyMu1r8m0V72PLYTIrZO
lLkHaabId4g1UHcPHkWyEONL9/H5cLqFXK+dHRnO2sbXa6uV5WBYszNuTq5Sbj9N
SX9xUCpPERVppvB9b8z31P2HtDZRb86F6c+u8yRvKGF1WRF2YcZ61eDfF7ZlJhuI
UhtSInzJe7j/pvRy3GxuVpC/mU3AY0tmUynXeh75syfyVyE1IndjiCPVhiDk55Iw
MFWNH6H3dXmZIJDiUg15aKkDdY9DQs7M4es8fZCTfeinKArExb/dsNhnL0HVvDxs
/uwcE9YnQHMnS4TBxBYuA/dJtPN+Ck/4fp0tlNydKQl85Xhnl8OqnTNSx4Pffv2J
wDr2/cCr4vJsOcwMzmmnf4lMvCNct7i+pdZljB/BT7G1YNE0UtO231/+XrrFt/dU
vBks2jCsNDcebyU0/Roj9ZlCdplwkrXxykooiL1qXGOKu20NktAEl8V/rDeGZHmZ
pmeqUcCoJbIbcD4LhIXqIvlPYyNRPC5Q2lSPPx4H1D79+nvAtJ/p1aR6wgyExuCH
M0KO8V7Ps3tFoHkb43epswPWhKnL7tq9geaU6sFAi68/+x91nf//m5REkcA82Ix9
tK0ELY2OVaKqLN92GcF6iW2eE0VmHaUYfU1Ksj8n1+rBKvdNnWz/ctH65cyBvyZ8
WjTeDTY3bnEiZJzxMu34r15lkdjy23zt5myFlF2fWyPlxFnQ5zvOr1U3pa9053Og
WpqghsM+inF0ol0VyxRlKuAyoJ4dlnYnPobYdBMghvfXnQxdO8vWzjjpVz5P+z0k
LKb/rfthnvZR3IdCwxCxpA==
`protect END_PROTECTED
