`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f2TyZtUdvJ5aCIQU8VSxd7D0UdQcJN3O7b39eodckLKKmQ42aDAq3+/L/HAi2ww9
jiAY7iiSHRLwtAsQuGjufeAeesyCA2oACoQSmwVZFWFi79S9gTqGkWMO1moWIqvW
MUIP+mqHKRMHc2ZuF/cUBdSrzytV6/puFsG8jefICKnRhpPdZSm8rWtFuAl4yA+u
eI/ATMvMl0gvrDCTdxEJZ/+CkKInOIaDMmexPU41MUJogVPelyCTbdVTNEx9gi0X
ALPGAlN1Fs7mGSry5lHL+v7aMDsKblUV4EWlqGU4VopgZh8MVx0mqCE4YKS0mZNv
Wr/kYgI0jdmRS556aBlB39HNnvlxL/TPW3zt1ljnqKvkOjq4wdImXabUFY4aSnvs
wjpLh6raN/jE3pg+TQ53T5/Tk8bcHWCxU3fchcQyA6dYOY2sG2iDeowoueT4VEPa
3vTGEdcq/+QHaBHnRMXR+rtITAhdFJ9mFzNCAe+zsrQ89YPyxeTkDjYBtm9sq3qK
zN9toUirNE3CeFGBtqMWzV61xsS0yyrZx5wEEgMhvx9F2h9JCyjWty8XNT2ZBIc3
JuJi1wRVitsA1TaLR18xTmb4bvOk1GlINeHjEgD62SX2ff/s0Q62eNP913+RvgPd
gahqgs+ghgZS3DSot0//gkmsgQf+PvDJB0StEhEn/FC22AHC3utA2h+nDncR4dlg
6Vua+yLpAV9Wbrs8YwfDLGInmP2Oa9g1GFIA1Tg5Zvozz7fgpSiKsftQTCAvTVGi
r8cm12Df+CYo4QOhFBG/z4vhzn5VWPlTUGnMLBV+74WVIAaHTN7FPnWnE/ehfkSs
GlAk92RKrgrt5fNNEjEGxP85bDNNtMoQcoBEZIIejMArUFjSLyC/oicpwgjdRKS2
3L0oExjUCZ2cpJGv1XOrnwaTf6Dfi7mULh/pbVqM+pklmCmfQ2fzhO0vLreeGpTk
cDffW1Fg/+G7PaN0soo7d71NclHG8BHBW09Fhufk47NvvZQls4FgPG5D7c9gGCVl
zW/Q3EQgigRTAAE0D2Lq1suGelH6Qc0dJ7p8ROxSrE6UEpSeLR9HxXgXkCWVbxYx
BmomYGHOlYbH1otuTTN8HhCPhINn5eGrVJtk3h5twnxGAUGJtUUPZ9nP2Iw2U/Xp
6h2K6rLE8jCohcwmOmKWZI6yz2WODfMQy/a8Av2jvH7PbIrAdOY5EsumAUzS7s1k
o6clqs1RgMoq2/hXU5ZODe0fj0t8PuE6aEp2bGWq5r/5Tfp6nF++0bocm6oBhcFm
JY+/KUZ9qCSPrSgLPFVJfxOHr7VuL6Cg3US6Jkzr1TWoY2uoljGjK9qdyLhssHOd
AAK7GcPEAkc56NgSbd6kiWwQgPT8dio07hUgt+NIG1f8/KrgqO1unc87I6t+f9zT
c3UavLHm75gMtn/v5ZMGErb/I7pUKBAQI9u27SQatfRASK7xwcgfyIX6i2OHSdDn
Cp0EVqcw8QHKVaRoV3+QLDZXG6JlngCxCjevkCh8U/9NtZrhB428I0oCDL9sbdSh
co0nXYcFjYnpNYwufwWNwdvTcZ3OpgZXRjrikc6hye6kIIOYE8kaIkAtPqS+o0CD
R4CVSPmJiaHElLm7NWh5aaGJhioaMmCzofj3yY8NiUujf4hNxSRLC40ZVKR56PLb
igeXqtLzbps9Y9CHdQfmQj1mcFrRtjTH/9QlaeUo5PpBXdTf08ufWcNOaJvPBV8H
5pCIuuEwZ8/LixiUqHX61hyrB3eUsmMLMNiOatRt5zZNtB05/455tdrypXJa2Y4e
9Ra8yes0nSZpnXzVDFWvxbVgKpHiZ+staH864+S0ohguw5oPrI2gcM32+fht48bb
4ajLeC1H0hg3mPEt/waMkyH9aag5Srnh3yWNNxLehGubMELSdCW3urzCcJXD1oo2
saC5ghucYbjxA/vtcbpbZSYVvB6oeQx/Ka0u2JB5Q2ALHMaThiqskVSoBCGshMMf
kk5AzPNgMdSUlt9/BS2zXcgDnlM/2vwfyNpxby32AyjDmWf+ZXqLKxGeDK9S8Lou
7MiUqaYDK2yCtfX6W4Pp6XMGB6TXfexSA1ClzpVNpwJn+x44gL4G1KgZHNmOwVOB
zRTbKM6E4S61Fnjs1FYzq9kT2ml3WW7qiI1qI1adh9X/mZeMgbVhMQfd4WXhQPlQ
oU+0O/PdG74KHvrtaFQ/YtpKPhti6jC8LD3/OUmdR2s5vXDoILGIlwJqnwtyMJzj
OIbhZ0wWKAg8NeKiS+1mG4bghtIodQg++iFK1wuUfKp7O68JR1V+GExcnpU5Skj+
I+Fp4+YX5+PXo+v1C2uXaNUo5emB+uG4FzJVD9X4nTTsngehAfuacfvNrpGoV7x8
c8KfdehGtva9nPYj1dBMwV37I0jXucOUX6yBgqNQoo+O04YbND5ClhT4Y7WDudSl
zVr0npRJFbstdKUbPhNytARTFZiHuXz1qc3ptcHtmZry23jYN367KOw8mYK6VEpG
MrCFHg3NMstf2ZAFPcCrvPxlN0ldUgWO6qaf8bXNMUw7X5/8c9Y8zcFP8OsKjcFu
w4adlovnWw6KsrI4/CA+nOI+1TfoA8xp3agAXhGajOmzS4KB8tEPiTopep+k81Ua
KPWicsICjq2xGKS9euEQPg==
`protect END_PROTECTED
