`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8QTq2tK57V7vQbytJkIKY3tuUsNaseKFIjhkFofklXeqUSeciMwXVU6vFVaPWfPg
NHyXkYMufPDgMaH6ocZr4ZgHCiClL9MB5sWBKTTP4JZQojnPOhcw+L37ZVo1FXWb
lla8sHEqn6TgjN0z7ESpJI/WJ+RUoty/WgtwpiT9U6FZr1V8I+c+hsAXKBWK7iZ6
eZ+O9fzbQq0WuySeScymEduDvxVNRXueqeTC/hsgM0EGQHIMH9hgzoUcxm6C8rm9
dLhGgwR7fDLBTCTw7YwWDNJ/3Hn3tPb1p64sREbtyU4pkBq94lsOapYfSkFZk1ic
gZt6z6I8tKWB40mvG6YXtHjUWXvVfw0uOEMd0g4aWV70yA7lycQcFSqjHWlFGwG/
1Gtl3Q7GhA4uC0F3R0/nim6ATP2mmM0z8cQdAqD8T8Lq3oJp/b9tG4vccMuhabcm
LndKywwNqtwEpnlkKYi4gUxePb7FPFMaL4UMjjiG4HEAHy5uNM/hikwuuBMTnj01
Pg8pkWZfHoipipFkA39M3hjwfH5j6Pog7lO6DllYcDg=
`protect END_PROTECTED
