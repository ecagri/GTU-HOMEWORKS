`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v+upjFvg16ulO24L6cuVpXJ7QDUbPpKsUQEft0f1Ifn+ZyTLX9L2bxa0dHJjdV+B
erVycVJW4JaXBmvyQvQvk6nMae33FFuSlq9cYF0xkr+2ZZfVeFc/niEWjZ90AUeK
uDpBhI8cTU1Xj4DMDnvv9tcfyjCrjmJO/Rlqb5Ra9acCSXJ0mE1dJPzHaVh9gsrK
NTz/aGs87BW1MOosVE5MdHjXv4zphUmGN1WYiG7ZoL1GigIwSzB0DdwAgf8kQtYx
CEeDGsQZkdbwFOTvo51kkGrfsBwHeVNJnNi9wj4TLKwXai0O0gwp35sAEZ2nS2io
UuxeHhzjPob0+aRghJ1r8YUkL1rExrorPxWtZ4ZUBxx/ThIfUIznnmC57MP8UiIV
i73hthfKpOcgBALfSBlRW6osnNtvsM2DmSOAKDIEJ0Gr/qML3LS/29H45D9zK8gf
bVHF02gj0UMkzkzfjRoLdmM6JexS3vdHCaHU543HmZgLFZ52LZgNpfJ4QuW7MX6T
GM2yxzuLr+NxM/yKdV+XKjDT85HejvqRONQwnZ6oEC745Nm4oUKch3EBTm0o03LM
RHMf9+C3KuOWZC9iq0kwm50W3HO1nZ/A1fR0El1vIcv1dWBHNTLA9Mvr71XBbR1N
+CV/1B0uDFJOEwiCTfEPNVg1tqM4AkXlM5fwTk+fgfF/jcke05F9YkwbMfC8+BcA
qzkIjxaKJgsU7KJ68w+oXBOYb/VbYdIT5McRvVAkNlEovXZoITshnuMFpgiyqAft
jyVAAGiaLk6jvhsLKHqre6eiXNH1OcWBjug5Ah2ShGF6+w/f3uHstrB+y+iU2AhM
KqOsPpow9QP2FFzMzsgkjlHogXgDs+DtGYT2Q2GNa3kt1efy+vcuoE7MJVJWfjIJ
8kVIvpD3bJzY2a46twVCuv70Zx/EcSTv2m44RbgkFSZLMnBIx5zqn77TT1oUKNYA
Arikh92DSQ/gIRzzAT5vCE+coz2T5766GiOrvOVgA582sdeekcaJyjfnzi8bgtg5
+Yi+wLIehqn3V2SVz8p+IC19+mvm9d85yCh1X2y0KXtPdRwPxuT5XEEtpJnWGkZ2
gAzS02zLWrw5OsGTVMIH/lLHiBm1Ak5FhLj9nroOnncjSPP6FP2YgZIF4Jeu3obh
g2mZHYd4o2yXAtUkF7D86K0J4H4E5r1h4tql0EgXeMYYwiHcr0W3HU3G/rmw3jw0
xqmiYj5/1MSb7GQePXaoR7Wu1ybKSdoZjGqMGap3cx9wJboEI+AiUlndwnjLztMv
S+lBa/tP4c4GE/CFcV4gOjn+D3v1bXco74YHvK9ilTGXzB+ZA2L5inVsrJYQoKP8
J2d9odCWp5UWNhisR7nUuL6zraiTD0s6htRkn1hmb2hxUCxsfMpVamETIYPkqOa7
TyPCUgGvX9TFuQ/p2JAtkeuKig+erGpdw1zHcnGaYEZPEHIu7YKLKEFMaYKLluaJ
KDfAl3xyc546cYCu6LRQZbIMAmpWDfDYoy8rxbG0RQfDyTxJoN3ieWgIMbqpnapm
oZnwJwn0d6crBddsMDywzrl7RknujQhka0mExHnjFoAb50AegpQoFbLRJur19Nul
wF3iYKRZi1sjGSXuEbHBg0hFifnmaBVdt5P1069FE+o//RomckOinfYIeoyQmWUZ
tvW1CNVoRdD1KE0Gh9rB4jhUfucUsyt0xph5XRcGzwpAxbxUZoXQ5lK7ZthEUfJk
`protect END_PROTECTED
