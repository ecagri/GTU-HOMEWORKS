`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pfRH5HKs4gURGX0C3ITUlF6ZFoTKRWnXY3zvJuFrcmdQu4/pKggtfaEPyVxCr/7N
anbaPAlIaQ8js40MAvHzuUFqm1YHEaXhW6T+MF4u5MhkKtJeE5QHHz1fZS0GwH3y
aTQj+J27RJpabLZfpL53XH57FF+PilGNYYAuUw6wKfP976r3U5qSEMtDMbi6zcuu
tQ0AOGL16Tk9aTYh9NHovmMduJWNwVvV9LjG7pkexR6A/P4SY3CAX65DXrkTpaxs
ewg+lZX9mCGGkGxwSkpY4uvCtDkDZZKatFE14AdqOJu0LgvIiWG5EpUaeQjEbIKy
KP6KuvEWV96S1+MCnrt4k/2OquI2kg3r1tDhWdS8oryey+dT1OTBOUG7/TTFhfmb
jG6EEffDj9jhDlzavgyuouEftwPwLarzSD2u+Q8we3Jpy7zwZEYv02DLcC+N2I/f
cDSBRUC3fG8ltLc9OCVSzvZM6i63dnFPn9sNZNOp9BPhIkpANiT89171B5VR2z4f
XoT8DHsMj6/vbP7poD6uaCjkL/8GqVBaQEHrR973J5msNC1mLMe+XMhCuzacCjDA
hubp1/DVayze5eg+yQ/37x/uGMzMztS1bAUIxBqqJDh3ftREbcgASESUExK6ka+9
epY8NOd8JZEekoLLX9l5aht1SEIwA2t3K5kt3V1lKJJjlwAZjYKOm02vuQmp/Xqe
NGrAzf01+WUFPSddUyzuiocFfF+dF2UAVdR40Bd/buWHMqxKHTTB45esXMREgQby
TmnihOMYKa+XVP9s/MKuvYsF49+6wOQtv9CQWd5dCEMlshi74Pu53prSMr7JQZK2
Fc8GpkwSd0NGzhUpSXi0sMxY1hxIELyuIdMVc8SApRvJLdrK2BTp7j1XKfLlocnW
Buk6fg7PuZQLkb6HJW3+qLgoXfXJqKC4lAm0/YTqs1Iok/lgd2CmuMth44d+FGk9
EXetMlTHs0EAUisNoGw2A+a8Iqogy5WOPbFkLCDXwwAcHyokcTSl7e8iot1pgr2k
e7ZDZQx+5vOB+bLL7qNDcEQ90GySNdQG2n5ATc7rMqoVbwWuQbHov8opU5MK5Tcj
esYBCe1nGMfv2LfH9XuYjQQk/sXh8YU8SnuTyW05HWgC6MmOiZil9m50tKdAZFV+
obGJJD1gpnxSreWIFZ3XY4NabiJKdZ+/kG2kOKZabwRkQRtuYY2Q1L4lJqJngGCT
loMec0ee5Kz74N7x/SYxF6yLR8kA98iwQP8zNya49jJ4hFm+lM8Dra6N0WE8OURE
IT0PukeaKOUSfoYIncHRWIn/EWx0Sp02YhYTqjUQFmrsUbSEuSIVPATkm6mHDZfb
fBy3rQsjScH6S4+eurgSaiXUxqRX1JmS+JcSQ/nGihx5gJfJgAlSjDfUIOwVNK5h
RE+09cqqjzpUlbvOzoJ/4pSudhjwH8amMWvHsNP7/J31D0/eHehHD2h5G2kFwi4K
D+WMvzPd7xiaBNobCtrJ36uyiN9OyvG8FnTYyICLeolV5QFmr2W253bNj8ekGcnz
72jMhcv/V/s5Wa39P6cySvkClksln9/MQj1aPTroG2+8S9bs9t1WgjPXSAheojUd
0vHwXpimuehajrqZJVL847Lzaj29EMY9sgghPugC+QuSt+hdcKETAs14vYudRFkf
w/dHQ2fCzS7hkBlp2e4eVU4dpVZDb1WfEPGfOfHG3enT5PMIA8fW9VdVsc3K4KUi
m7ISOEx9vZ8RMdF1+U+mrgcCPGF8yDmI7qG1uejY3comxhMju4yfAO+aFoQ/28WO
2mAqoM1jKG32S2jtTDJgpBnKkYGqR4zf4EBw+q/1LanjWF2CzSYizfQza3tKr/qL
1GIS2Da+t2tHe5K2VNCZoUOW8Hg11/AsTI0niD7DwhfLseURcNYgmYKa92Fpfl4V
ElMg+0ET4a2KGfHyXNpk1MiveSXS6DbkEXrySAxIJcxagYo1YgsLRVnbbMIkH06n
JFn4nTynrZkSo4MYB/2Z0sFfWEvm6E9nPEsDJTXoBA1JsnVDsBW679AaEUo01bW9
AiWLRscCq9n+yOf5R2ep6CEpp7y+v7jn5EVN+oJBfdIstGTuqdyVAzyGRY7vlTHl
HT92wCUL0/opFjTbdlGj4r5NwRPWLacIEhtoQ/ABN1S80oJyaDw+5G3trw3AY52M
MBKTtzX49jDlk3lfLNN2lAf9dQ1u81M54JAySD3GpYbKor6q+zBF8p0lWsbguE1q
nQ9qtJZdifG1Anzxm68klc2oYBRdlu1WjBSDdub705wJT+pj4SVKsu/sLMlga6Ro
XowC1d3cPkCeXKhTzSBs3TqCxJWY5McfJ7ejz2ModmX6723S+ZmRhV9Crc+Vkb55
2qFwyCdcy2Ef0fVgeg2QRkQlgxvUp9IjXS76VtLO+y8cYSN0VQSzHa+gAhzTdGBm
kj3LiEqolETXHDe+GF97AxhD0pMW/F7raVlfXLmUKzXS8Q+2Uq5GQNi1Xj6gcz/s
nv3pqzSk6nmbkGI7dtT8NCv/GfxSYzL7yZSCBs+91/QPEzPhjYyoCZpVXtImyFAt
2kORdoLx4AW/9uYODL3kqw+wCywSaCHa9fAe3rsChsNc/Wfw0D6KqqXLvTZzMIy4
0xbhLikfgVbpNi8efaMN2beTd5TG3R/RosLmLmuFMCiZiJ560o0ZuGF19tEdpbZb
m3+T3tjUT07SriX834qdbf74yZAfHky8ogDr0/hJYbTRfgLHJHBaog1e064RPNnL
ucbe5tEBB1nXdju1CEthiETVv79u8W/ysZYqjQOR1JN2Ijt3h3hBcEVSGK6BtxL5
P+SfSFB3B6VYtShzgmCxJMVtq79JEWPTwFApWL2mvoRVo0VpdIo0KyAb7LT7e3Ue
zcV3/guAYXlI7hmJCZ2eIeAAHapLBqTBFikY+YldIXKwr7P87OsuQ5D1Paft4C/R
M6r+L3rVzAmCwz+T8KpzswcPY9yFb35NEGZe3o+dl1zohstL1MlN8HGyQll0mDYW
gK9FMKtW0ht0G1QXtA8Y9XQbLduZOMgnqIjTGk1mXA/apbSi5nqlHbLAfrfsNT31
m8+S9vQgt0LJORlkbI/WA3WY3yIh3JlJjPUlYc9he2sXn7ay7d8XT6sd6K/FAy1O
IY+gm5Y/dpnbd7UgFIS3nuDw3PgtIIP95MVxhisdDHA9ltRtUyRBsuYZ7VqQET1q
Mtocpa7mqxhvFkiy4Uv/kJ2M3RD4a75xz0bfdmHjGRuX07CmYcQYP5dWg8p/fKCO
JZGipM5VMd0+CplEG7cOzW+gAq63FKzzyEz2PPis+bQGKPWRxpKp7+6/J7R5jEA4
rYEfngufmwODtsoneRwcDRcOkJeocJAF1ohz6XNo/cBLkT0z1VPKtEkG4IWu38Il
cLtqvEXrjOAyxkPYij5/Ij8yh52y5WO7HnbFqjkgrL7oYHilh6aof3vLQknlQmDz
ZjBmnttPCaDvN7NolB9SYz0ecWIJRj8hbN14krfENknz+Jp08tGN1VPFlyKg3Iei
uXJUIWEXPhT049S8Q1WrdqJ6D5IG2cydw1bx7cU7UbMRmJDaeQPN6+gmsTbaOUv3
f0xtQePFJ2C4KQiKjX9PnT/QhVjVoJVl8Lzc4rZWFC6D/bfgCgW9Km/+wpXqjOsY
kK0b6XHtrbEDJ/oH7rdslQ0brmaqJMdpt3SB0J2PKum8eYd6+s98/q2sPWign2tP
dFgzCKMo5MJLJBGcGyMdu9hI3bz2GpiLaWEXHouewWkqJFRfyEb+wot5NoefMAL3
BhpQLVSRw78v6wJjp55S+QJxVk0tGXEJ7MAHNxmLsp53O0LiJAYKhT0Zo60IAMsc
pi43bi0WLtwrhFCRp6HFtJZuvZEc6CazXpLLtfB4fRWG0nEJCsHoL8E/QlLbNd7Q
dd6xNZUP6u8mJXBzciSj3+oek1EW2rSvM9FqTVe9B6VO5f4iu02BZwYLV09Y08L5
EB7Dnm3QXalGQbv18EewNqlGyoKL2rKkjJwvprpGR8FZFcw6m4exsxCCVPbeFSzc
S0nJCXGLIc72VK6zY7Br3EwfKEgl8GO9IKSV4DuGQsmjOKbDL4gZx6LRwyO4xr8U
o82jZzdh8rkbwNBTr5XU6ffGDEK8dJlbi7SCg8GwU34wNgi+NX70XOH84Co6mYZN
SGeeTWg9e4j4hCzxSWNLwo9M+yRlSo9mXbqROGnXigJVwQX0UYwzUj/fDghRskkf
f6ymDn9zITjh1Zv/Apw+xTCm118GVELslKJpUSOB7xCuYnnpF8ruDokDdXl7cxIs
baP2DLhUjjMrSll+GFAgOqtK34sTGZYmh880/BhPMQE8zhEXf9EPvP2yCf2q4Dbv
olbBDpQL1XH0JW8IslNIFiNDMQawIfDtiBeG0D3yPFmp3C7dtf7Anxl/AUHKGRdc
hEE5QTwXzjM5/QIpUrd8NrzSCB3cJ+V3WWUAh/nEPyEY7gj1gm5Qzkgju+0QVXc6
+zPUvta0KXUP3jpeuDjN2GyWc0K3xj85fb29p4XSHXiMinHKtcXVnxEB5Ovmbk9I
8x1pziYfnJqidZQcHzi+98Buhg7tQs5rVVq35PEJkPFZZtlU3mObNKOQ3wNyOeUz
MlwveSZmATVXtv7OqTWrHBAZJ/CJsRseCEeL9DeVa9MDyoQhjdN8Nsy97/C/ozl2
i2Gi9oqXupQrLcrW0q6zbDzgDK4LrJuJI0c9PXp8+16W4rEXkdZuktVG8DaGZp+K
bIv/gSasNYwMKYA4VgmX75Uh9vkiYGapJeeJccbupJIgIdghTSSqtW5MpZVceq04
wxAvenPE8bExzxZMy9M4YBAPuW7jNf1iKDUYTALHL2auqPYdtYNIUUA4BNnnPRd8
n8YNlbBs304oK6TM+n/9Glrp6MR8XrvZO/R4+uRXFj6Yg6S4hkXskBhC68QfiDa9
u81axIz5dPhko9f/J8bkqXgixoZdmyI8xLLGxTcyVf11RaonUFl3kL8wkAzJWUed
yov8nNi395swWuoZdV/OtusrPbTI1ha68JaUgAgdbribZ4zvHVekO8hM2bqvNEje
zSpFynRl1FzIUUHwVPcIiUg4M3xxT5Dh30mGH+vof05qVUX4v7HISTNeBZsMHeiR
Z2EIpyFZ4qOpjWpJaz49I0Ibp9nbfqtmh8kiHpzGntM8kac3noO3SHWNAbo0Vo+f
3wLH1Zd+Z8O0AdfHT93wFOwcZvdAluW7OJJ683SNwUDRWJQI5pvN4O4jAcnYRg+T
IOn+uPRrHfp859UfaUK7EDdgmhbmSl0tmXinenGeQf8wHsgREKDPl98yUHIRpBMf
zui2ebFTR6FZJwv6YZls/z14+FnxzZ+s42MBa3GEklH6tHyeDbwJDmar4qqHlhGB
uCmHOaSUCXILAE8s9/awa7eoXSnUepkbeLiBjip+EcyqlLDoT4PAtihPbU7Yly3X
enFuJVqC+cHr6AVAUQs0N76VCmEg9bq+hf/JSARvhyuCaUs2s4Oq6Fh1fMlLsylj
MBTgXIvIGjD1v6E6SeEMMRnNQeIpv9mpFFUbnE+rMrDnED8a0UfmEPXsPxvAgbMG
UKsh8TFEvi83+4955BrUf3sFTzgQOC7X3130I0M6COiZLmDzyhDsXDz9bip9Pdca
nQYHv5HIjjgsxQ1t2aKwnoAD7UE6RRnx3+gcKqPrlqlzR4fwpOrsDSGxyrd3Detb
nqMH4jl1kNhD/lrdWGFnqyiHZ+CnKAN45PkMwoUVRyRFSTVTm+oWbabkMoyXPvK+
F+h/PnzLrJn4Z/bzw4sr01DbNcsJ86VVpHe/T01U78INU1nWB2cju+/t70whcxjb
3/n4RzZOzUn/y8aK68TZcJCgJVG9ovfLZEiujBqjJau42yFZz/W8pdA6BUXZ8EPn
Oo4Ru3vfHg/IWT3JZbee8GlDuuHX9bwXEfHCno47qklhvy8V97ntkFyaDxFGCII3
dCLQj0i2bOyTF1ODZKKF+rydCCOh8TKmGGnhSNQUS1lapq4gJVhe4Ex6qxbQgfrd
+7X304ACcW2i9DQit/qym6h+3oKYQbBA6dHxERszoApAfDgdYPI7f5AsvNoU0W2B
Y04McijapbARNH209VwVND1sIoXq8F14ucRR3VGqfVMX7+3EF8bDw6nqQmXQJGPr
E7+zs12i1UcfWAixoGH+K+lRxhLecdBboNmafN0DN1lGWDRGVmz5cA7hVa2cQV7O
uYbWDxM1UwaET+WGnml83F8USH2ScO9ds2yZqZ3TLXJMID3RypFP0iEZ/toekQGr
yLO4RX10Xhjp7+i50r8AKf521KHMEo4mXWd23CoIgxuLxB+GsWdmKFfBqkpqgv8S
yUoMUhZdvIXp7GzvDIFsmVeq6m6wtpFmY+kUeQX1nwQPQaJrsdER5oQ2xbFjmHK2
+zzXjbl9vUPLuu1X802Nyc2FagbrKq+fpTnS0bp2FW3xO/fXUofvbmgnmmZCwrK7
HL7s5wJiq6smnnfp9Km4jV1ei6hIxqNFBXdNr6oV5s2NdMJmug2hDwIJQrLIfK+h
mgFyHhVTZiDPNpVO54nXLBj2Re5T8Ng8FNpgHzC+NYxwWE/k00Bm0fA0xOgxEe8E
j/8P3oW14mKzzIZCvilu15pHMN/adA98CGfuxmurH7YITn+zPV8IErQkdDzdWB2T
Gy4oggewbMx7lxS0iw2fwBMklhuqTHFgj36vXp6pxjj3y3kaG2crCYK7Bt48KosT
1glMdKrziyxPjzgWlHpIFK8lpnJF/qqJTY0qvf5zLH7NjBzz+XqoIxx8hNcIPh1l
ZysDKUb+W/mJlfVo6p0T5nB+5EFrgqrieOkcVksO4j/m42YHu5nEHwycs2ut7bgm
yEZ9d7vVqpJe7JRFs4QYsuQIXAleuigeQ6GeDjc0MhSebPYOpx+lJWOQcNLWOZdA
Fe94lGHl0jom6derK6oGVge8I2Zm3MByz5MIY/IXOXE3eJnblnvUfZxOFWha65Q/
hRWnU9PpzG5rBzv4kdfJAZJ7fUksLT6BMWRBbbXfaMSP6fr6kmMEMgRIsN2d4i28
p9TGmq59MP33/kDl57s19ateBAb3d1AZs/kQirelXkLvaN7WhSD1JP1VjhM7m8lB
91a+v3T/fTFOa7rwu9+g/tQi1+VxWtw+ubaCWXFCuzE+MtL24TLmP12aOTs4TRUO
hIKSSR2eOrqVQyT3e4k4/2eqCFVHib0d4TUTjkGxxZOIEx6kSkeAuR8uRLoGj15+
XBUJ7RNXusGhvZyCvCQ9SxRO7Usjvq08twAZ1XL8m+Rh+ra9y8hD1n8OFiR4L9Mq
kq8LWj9m4E7OA94OKdiIprSxWW8wNQKU6E8DUteid2b89U82ufb1KLz1Y/GoHlE9
Ix7pM/rBuv3wKV04dtVgT0jsDsWDNkir6XMhqVZ4YUOZltu5mphooVBeVsnmnfZq
02yjIX6ig3+/0/RERD+S3nBMIqvZVR5MJFcsLdL4SiBlrB6V6P69ATUBhJR1OgCS
GnORRPz6ZqEneOyZg1uOIp3HaOcTsu4fHe08Pr8y76sxQruiC9iV7zLdshIilRhW
hofYh755YC33Z7I7XxEX2MeKp3LcOA/tiPHrUIw86rgkNS+UpagS0X+9k8ynnwVo
xg98poupAHJNfcuYyV7u6piyDqr7dXlAv5fJPYactZt9MrncFxmiqgzSdiTU0e51
v4ByfVk7Yb+pV6uxdHT9ryEEUuZJyUJxm0fuvebEXEsUgolF6tj5bvdCEWQni2xJ
yDOfGUcN+RhuqUrueIdvzLhoOyC8WL0sMLicogKQjNIdAQd6Im0v5g5x+xpi3kPd
jGXt/rZ69+kfDa95EWy4V+KTnsDaLdn0XdHDJEG+caCMi5gyrtjDZeaV7/QgF5Eo
4RB0mqdzjd++Z1s2WXcCRM2LTD2uBqi6hqj/aCXV4vyATAx1VJsu/9Q6ckzNS68a
9W1kdEngt97oQHa2mfxwBcMjzcED6Bvo9T1LICYqUiycQwBaHDWb5L3o8QxKOhAE
vcctHVs6NpO1mvt3zQIox3m3lpDunbn9+pQzycDD0hgV1JaGlPR7PAjfF2Y62ZWR
luUB6D008f3Xh/JRtyODKculwFezyHv+PNEK2akK3DgUt5j5KYt7MuXbTXoJUH+l
Ar64vCrwKWFxAQArGYDulYUC5IBp2sD6ydkYcYqsSCwcLFVHg2ko3tWz6cN1FI2e
Jlr4tiKraf9xA7Ft7N/aTuVgAN6eCfUoXCRUHNPPzZV+lNhOf9vjtVxargM9HeOR
cFrLWKHXYzIZW3VjuPeaoyt1rrubHiFOwT9yy3QjkLmYJOQ34avz5/0gtsaXcc/b
X2PNeoWA6BeCUXYGYW9+icEUY3va2vwVEYWu+uIE1lZKH9Ao+W0RXhsBOrZSchGV
0BseRcJ4ugfNInYPAf1mOjFgO7sNFJ/kOhj3Wy45dnZlpsIWBUwiT68CJ8MIdgf3
KMCjtaZiDDecqQsT5wFJQL65Uf8Uw7tney4o37RTe4CsOyO0jzeespUrKamY3MA8
DiMBDzMa1ZI9Eljtk6k3H1xnIfWl3zMzfyQG2DuIYDCoCN03E4NjXFan6Dkcq3ED
wAf9IpSRHoCilTJ331BYaCTiq++IKtiwsNPC++iLJEh7qcmZNAXL6u+nuD3tyhEM
4ymrUTFJ0de9gCdVh1puNGV5yV+zeVlkvNcxKxYyhXRAHD6i+m3Po/m3axZw/teB
tZcPGGGCrn0qF4Vn72wRQDIhsw4WIAPecfx3fwGzGiHL83evDHlaxYCqwaYBJJbY
r4ZzusAfabNOyWmJeu/vtYWm6abam9YKddsDHQObQ6DYzR/Y5sYXJpbRfIxAliRg
EnJjYhfJzeTVebi1ZCkdKM2gpYG1dwIJ/8Lk282v3QZ5JlxdNGIb+Hljb88dyNZZ
coo0v6z6SclVxPNyCEkj0hMDA+qb6pIbL68NO/tLd3KkjW0Q6mXT+RjqRjBUn+xu
kthK2Z/yNj2/SjblYL5gdpnMBwMpL5ATAcE4BcCwAEwtE1RRvDBOeZXJ+VAMo05r
LV7fvZtZxms+nBiBlezJiZUb9xB7X5ZPqT5L6E4eTcNwIDA58QYwlBcXfdtjOCtk
SDCKh1uowXr1WUW80knDwklQGpblpTnfAzAxXNysWg7dzG3QPzlzYyF6GJwEtCd3
kMXYIo8y+niomoLv/hnK7fgniimGPgjRgvQQN5RQc/lriYYkaZly2g0LreFkdqpB
/MZmiqDmdOAobOZrHVOfqvfUhZoQSlzRNfkd/pAsbcOelTw5cQVEsVd105C2bO5L
sl4qKhybcSZB5YJjUO8yve3tLLibUE/+19NTyL0qFz9v66v3lbnY3nAIpLdDPJKO
AHErHXb7pqpw3h+z0/KdXvqkhVH1O4SwqJVPD0kUI06RJYBss2Z6tK1gFBJcTibm
cQTLCjYwuZGlRIPnKd9kSCTPqpTsMxURxPTHhXfEh3gHqckf4ZCJ/zFDBQoHoeZD
l6Ax4DUwt3vSgqiWwkvysmjnmOymxAY3560ItL8C9LOTFyc0mj0wibIq5JAU5ZQx
b+5tHjC1c5f+3VooFYu8cimnaJzv4wmXivfa432GBWeRC4wcYeABEIbfBD6Ex2Sr
sdnAcOnzJSC28RMgZLwA+K4Qgzpmi+OncCf51F+KG0FDpc96Upvzzcv4og3QeH76
rBm8Adev6FVNaVfDARzwaqQ9JMXYySim1WY2XQI+zCXiboqmqgU/4jmD0Kfbmepl
9HhwzXxb/Ixqh5Hm473AhjGN14p6rUJ/epRwJwhY3KzwRQ+zvyLTml1m84AFCw6x
DP3FSaG8xsxEvQkRCn+wip/TXAZnau5elIEWbpzmNybcgvdrksti5au0i9AaKiz8
lIdwmLX7SWCSkE5uG8BBUgdjNi2HrXIH0CvnvbgEg5Hdymfs+AeYJrZtV/XiNFSt
jRVL2fljgPhLR2lbxmSeNbKE6TAJH+19U+yGLxdTIgKkwCgHwL0gKHpUQaNL++Yq
pHlWe+I0XTAvVugXKil90t2NnY40ayKYQOW8mmMRKpWvAf7cXJWD5dgdWQ8C+9bx
r4N5UllBQfX4aXjYE3a78V+ncC+EAD/cuhbbTklWyzXS8CgpHDCrqiuLZsdx33UV
JUDvM1Xcr9VMmHabqpzy8E8xLBrYu/jQBq0HNCfIu5nMFNxFW6Tn6+WTg6NBuInM
rwyroH+bFyDp0lopbKNkFWUbTnDj8nOKgLw5DRj/D8gSFFx3lLgjo9aFxaKcAXXl
gCzUJ415n9U+GX7d89lBvenxz4qW2wvit8e40y6PJ+mlPNBlIDStjNXx3L0JSfAs
awumENTbJuD30iaN1KTrLz/uVJKFJVbQwdhRikIGbx54QV2E9KDrb2q66KptDYPf
as9LNQhbsLWfTTGfjjZNVXO1CgcHlY91wnn0ZLTZUxOPQz1T0UMWl+VTOwX7g2vy
IjPUotGco254Gf5KG1rRbLKbZp6v8XC0PsRMu//PAEHjbkAUPNtJRsUolQCNE2k4
8sQCXjXH7VELFk+6aGtFRM/KsuFI4hiDsyWn9ovV9ZCSePyN1JulLIqyXQGYl0s2
Fm+7noKoZ1nQnLO5gN5yEDwR3tDh1r/vFGN8lta3PiEsJX0BTsfYkJWgehL9wENa
1SRZonmE/PX3M4Dah56CX2MPInTSIAuV+0Meok0qcJskZxKfcMnwEqwVB/QLTfDy
JBCXpy4U78Ij8FuWEqUen8t7WzPvni9QrFtVbirOzNkoRqkPicCO6vZRaamXWYTI
JTid3EEh9CaMOpQPnSN7LNJOk9x6kARwPvKyqR1susC2GvyINZVy9PyvHALHitQn
B7FKO1YCVrjfuUtkcEVxYjDzMvzpvBEaoAekKSwcR5N/saEZ6UAyzEXdDo5bWHjT
vObwYetv/c8InBt2qSE/EEJAJIlKSmnd+9VbYwWQMNe46gt6F2EpmtE6GtMtUWag
yTpfZn7biq4JmIzHTPRoveyeqRPive6ef2qNAGaXly8Xaz4HzNAqMXLojXH1a2DE
VbnRV/YhTkoCv6FnSo135+3JxVjGJjzEuELLz1Odf9w1slm8vyd7WpW0lH95wNiJ
Tku5n1hDLSLB/2SZz5IybC6/BHtENOzlRCArxb3BD8I9ghYV43Vn8SFhX1c7yS2U
vwIEScKv2i0wXpaKCrjAtwE6MtLr/y4O5otGUyTooX26uEg4xwmrWgXOCzhu064R
M0s2xGqX5BYFPkUIDkpqLhO3TZ5SY5Jkq0jWHjgBYQLZCbPiIesyWi5J39Y2SIIJ
gQ+cN9u32PtpmkrVThlS7NXijzYrO8HPceFPDTOcWr/YJvkXczZnxVc9y+KXJLHt
d4JKdKkV0nYXXq/+Hec98+FJqWuiP0Gl1N3cnlujdOLGbjoCo2E1dpZ8WMbYFtZl
LnykTNfRs0FjwgQ4Lc0sAjv4d1OrhFcV1xgg4uOHfgiKIj43wWe8zPyYOrk4mtIR
jbS8T5UOb15Epr0H5aF0OCMy/8uqBaI7zQ5Qms+88j4VkJHINKhz948r9YGDHRF/
s/elyDhu9fRNeC/UVoQm5l2lhAk2hxQfhV+14eyCgRQWvm2oQMW6MlnEolSm2fkL
NBn3ikxB1D6gjLyvJHsLTIP6rTlhA5DFlK9y81kIYoNWG+4xVZaSREnWFVPktjqi
2easUjCPokPsit7WFigKr/TQxWaEIfZ2pgMtA616c6hOB3YJ9lxt2jK8ykld06M/
0JHn/XA0G4aZf/gYFpPHH2oYeVRlw4g7SOnvmi00K+jcK4F8oy9NRlsHpmi4GZ1z
C68X8hu9tWKXmPXS+G562ydd2wDEaWMQ9VYSvAyQUsff8qCqgUJbJecGmeDkOIZG
4m3qWoaEEhu+bLKaHn8bhBKGO+f9HHhG3/7+IqkZoVWNDmqQrbL6rln7bVQu7srr
1OzUcqKLXJPruEpLiJ4HXODWnrbrcWATCK2hd4NNtZ4EZOnXvKoJ2IIijgtFyQvF
2yGSNfiLDA0DzHW1mZVa2SN8PIK7MxItoBe0P+Kp0xu/iPhPGJ4W4pD1xihQThxo
kFwTUJelWQxd9RoklVL96+OL2w4dNWcss8Y4fsc6KOOerYhEufqwSjAU/yqM+ndQ
jybc3uY1d+/jRCo2H5GAOHvt3p78m+awSB+Dm1GXlnFppu+uCrLmtLjevjrb4P2h
8HhKpP4zVpv0SHrCT/PBqDMAQHAC/yGNIhDd37qnjmLrN+eoV2g8ebCgKDcJhMcz
tDFbCZJ708bZPC15icXbGa7l40tN+YQ7FbuQ9TSrQMs42yk6/BEKU8l5t4imw1CQ
5jSAA83Fkx0S+LBbVGsTc8WN0rAHn4LC1i8L8CKJZYXJEsSjDuUSgfus6LC2W6qI
Mj5yXsRE2VEgTvio/9Wjakb834inwWjgaKQcBb8TqEL0nsGY09CBDQw0y78kcK/D
/rz2OfoVVR6AiBcKSX+0MI3oKgSi5mKUa8WGkdH8ZfrxEhPcPY/Z93jVR8Jy7Haj
apAjcpwveNclhm6R3lUC58c9zXoy+WURe1Gr9CxPh6u3XCgciVtE/siDGzqvV79c
Ds/8Wii4iqZvkHaXFVofR2prbeNCL51OPnUJhW5nd8PxWCJEx1VMB06Zt3+Yov3D
Ypz8DTiqE0qNjePQWp0gl1mf1Y4zwyL7+T/NMc3/7hTG3R+UsPQscwI8SgPeEAFU
n0YnSsjuV1gvz+ftDSF0Vp3Xme09kdqbUHwt1k/rvkv0Hq+h8psCvzy7xGBJaTO1
BMDmYLA6/QjEfmPhH1Nd1YNlJZcO8cHQsyIDnCHpzpEmY0aBX94G7jLlj0Z2JbYE
21kUwRUcMaIeq+9lNYFM84G/hJ3ciejwqCVVOwHt/oF3/QtHa8BnJRuBlSjPc45y
8YLWBEJniT00IyAcKn3OMdVHXqojpqokJt6P6qfxv2Yc7ui9ckgEpaJaRSE9RbvS
MnDyjgz++6a5Ihe3HdGznG3tNTSL+Tlq/A9uKgDwGSBbVRDm9ZKBGSEVf5bMzW0k
W8V5AUJLftE+ktsWWNw/cSviDInmbnw0rUQIJyBX0BUSThfLJggKfSJn3Ew0wycc
ZFS0dsnFTWHtMdXNBYQCFJMbLtSVG7TuVIU51W7OYj96EOUMc2wSaCJ+t/a84RS9
mDE8qyCN+ZkwyUVTCo3C0abubSLszh+GwSLBjuuwAy5JhkUceyy8zhHLNNY8X640
8+wTTyfgYwtSjVwkpall/oaBcICbOZf4ReFvFTDkwWuLB4+6wDvGGo7ioc+SuSPd
VDOu/sYen0c92Khw9vwgOqH0LPfMB2aPDw3EfYHyNU1IlR92KcJkisNeSNs6anuQ
bOYuEztPL/bgw69PP+U3wcOTapJbnz/Semgev9elsluMnjBM03s6AUWehQC+RSoW
LOxo3oH8jNu4xbD4vMYz+en+nN+r+3E883Mf0+Z044QMNxDMdc/+s35g/02mkV2+
cElxOFzN0AINO+B1XTKyXjUnK4VIks3xkNe9uPlU7iFtuWt03hlQROiEiB9ffGOP
sTpko/A5veV1D4slX1yxhFM5XVAEaugaipEH0cj2ARE1gZI3PK3ccfURmthT5rt9
5EoxK35R1GyOk0ouEY285yz52XlnTa48BhdCtF+ClnAXp4UMvrd7gsl2jQ1ySNne
9irk01JlYPUwUQVE0Wz56GqLGYbmVHfTfrqflgBIP+LcnBKHxEPaQzKx2s29TPxE
jHPdYYrcl7DY83XsQbCoBXngoh1KLaT3MOAqAvnrcrDVrTnpsIitkVTN9i5oqmY+
fbFb3lhxl3Nc6jAFJ+f6a1BKk5mUOBegUv9edP/PGO7c/QRSwTchCtmKwXPtBXtx
2UEb7y8kcJqPJdlE2cutf/qH6JOg30kFP/OxEVtt2F+TC7tCRs81OEoMcE3A1MRh
rmJZKKlwc0cGFrXUCBdQ9SZIaIhGcZ86ux0rHz4roIzNnCmDZuoea/hWGe1LUaUk
T0vqphH8XjoQbGyBGJid4FYyqKh/eETVRFo+LOnft0heygK3Gg7HItkRZXM/Avdc
Q8HghfUFBNXRjQDz8naoMIwGTMWEg4nus+j/pO56fMrK7+qe3xiJZKJ3+80688AU
WUhtExQY8/7mNrDH+qygXWbMvy4bN+/4SjgqdZXw3y7xA9G5fsW9kSdoboqlmrsd
cswg4dva3LwPVuhM8Vz0h0XJkyLwYePy86EoVOW+lpjQ5jnGvGCcqvo5sWiFS/a/
q0pfxaRV8qW3ZJCON0c2kYilKAjOKUo8PJKt5Gj3N8xLAyS5tOL7rlZBEPqYTaU4
Mb0FvGSb1gEyaR6mFqqvD+q1COhS0xquWpNMv+htd4rN+Nnge21/biqzPCkCamad
MAqdreHvjtVTmEEAiEmg0n7cke4jiYBWcjyrpglhiv0XPVW3tpifEtU2t7ZT1SkG
CU8Luf1LfufWcdrePOpoJdtPg+CiJg7FE50uAMA7AsKmYCCS/fF3lqkxp0F4g8HT
YIJqfWNYRILKlsD+Jh6unEWwYv80zfWEBzyuXKy1y0Pybf2Oat2jYd075sqxCOUT
ICAWRmT1pU+GHyjHesBvvJ3RC+ZV9w8hZUhw02tgNfvBT4eJo2zkjYC5LSjyO8ju
muntK1/vEca02wF9bUv4Cz4m688w68lyjxgOhL+fY1RqwjTrjwPZRGPEjC7WaaNl
qo4yGVdG6jjeVnCA9xa3vALGwKUKUvpgUxPlOv9c+i2x2VmSgxAoP7fS3CpxAyq2
FOjY24Tj4iP/+wccZTNq6cLziwSNXbqIFA+eYi4O/9QWFEQFSEWo9wZQC+NB8AI5
Sag9uhqVneg7K+FiExNfhJKNF9ekPLC4n5VIJ+rHnDhDgDD9HhYZa9DBAtGQaBi/
9IAFErixO6BLOQz8TDMvPWB/HNUq5gkFtu/HdJs2mS4IOCL4TMM42EkxwF6VD3P9
SKiOzaHeM0F/ZUJqTFSJ1yT6LD1MorCMXUP9PKLyJFuJ9c1ao7LfjejtGZy7ZVRs
5OUFR2WJYSfrfNdE043ZWYrGzK6kmf9bh/mVtt/myTtJiEsWZQI9+ZzySt/fwAfI
1NJTN851+GxznR5wEJj3DxxqZWN0H4v81aEZzRlvcPD91GkTI+bNrvATudUJ5Gem
Sh9P3OgdSbaqrZ1ZtguKiS3Ez+77pXxCqMMgTN8osVyRcBSQSafnwq9bkrie1b5g
gkl4bhgdcVOL6EcgwsgddJNth7l+YmsJaIKU83TfRVutpeHM6IJymzdGpYU9MwA0
m2yWPcOMkdaI7omjAHe/xG+VR+mzmv43auYf8zrGBj5LykUIMlV5GGOFYhqL59kv
dR8N1KbQ+QWz2KrC9pj5YgALzsdUD+kXrQDvIfqCsD/KV5zL93h6+NnKtQ8chEy8
4L11PTp7gbPIX5PqfI+EN+kFHKfBP84uP/hw0sIXuLlP+x1ut9nCkczjOoYMZopA
XkfbE1qtaB1UAupM2d9Fq/4gXFHa3OTgrza4lGpYLaALpuEdKkVuQNfGtM96bAMZ
SKjZzNkysHDeRjTG6XzMOAWgH4GyAtgSjymJD4r1hOJ9m62DWHvNhBhhWSf8D01m
qVCy3GSWdM2vIBw0jM0CHqB0UU0hYeGNFZzmBKKHn3GO9xP6PjsXK/6G8SeCGaFi
BEbhhkMKhRE0trJCBsjtyHj0MhVVcYlJxoggNrZDBi8bhGZ2OJbvLbECcaEVGo0X
WhgYMz91g5sXaCnO3EDZnYsNMKPImA8VVP8+Uutibr3Wzny/a9rUU6tBxbdjK3dS
ByhkeJ68mGqb6swGVgqKpwCFbtGSiXrI5CqpSWBy8kTLzgCnrjxqiw1GpkmXyxDz
/dJkJduRUUE40chCEj5weedl1ldfstKD0ScML3Wh04POfUa39USzRZM3KTwDxVy5
e1K9+ZpB+KH09u5LrFpwDd5l7/dcEux3hkqaBvH06tZHxhF4i8QG/28zi/jE0bQu
xDNGvRGUhceLjYE4VCjQ+z0bDAnTofsRIBlmbkp8xnfOHWsrDlFUHfQ8ouCteVAE
pbLcAwT41M6wpEaDOXz2iURgUB+dOM+81uH4/XtoAZFv1yGz0hodacTwpt4idJra
t6hktdXsgOoLanVr6tOgFR0u0DlGsgQvPAto6YTFuJf+mC+FAlqoROWejCpw24Fd
DzQ9EGkIFG5fCsYy43w2Lazso0Xb6k8nPwyfPFigxtjzzo+kklQg/3z3qs6wHpUX
6OQnbzk7BMRP8Ec7IP2h+LYIHPB+plTvmUDn+ERzz+qQqLUkzSv//KknxD5sL2u2
Ttjadl7y2hifRv7z8YyjRbMMCkbRKa2FrVNdr6p7rdZLBCickR5afVhvkVjZk5Hj
Aa3U/3CdBH2H2yqzZBJNJotM8DUxMOAGoHz1YNxlp1mcVRD8kCpZ1kuXxrDhh6oY
8ZladGuk9z87Dv0vU98d5iMRoTIbbqsfeakJ7req5TKm0d4fHYrh7UXxyNQezjak
8YTu+pA5ERAhD6Me5VKpdJoiobx4E6FaYQsScgqqPiN+QoQarXnwE5hW7k7Ft5mc
TOygkXdNSNGDcYIIDGJaNVBXdY8OwGxNVbyHC8larMI5zhFTVgtymauyF4LSPinv
rYNu0AVhGkZEd+R5amoPKQCAfnZFum2Z8iE+PuAepxIXkgcAZVBCRCXcERbEPnUq
qdIWhe9WEjF+B4uBDY7Pc9T2RdcCMD9w9bneJUkOFKR1yRjzUfTcOB/wXC+71Y7d
/agKaKIwAyjm0ahIIg9VuVuuAzTSvzNG5S4/IpkHNkvnUUjSyoMPMJSrlK4emM1O
HJ5lvndXrPzO9wl2/teFDxG+HIhcks3P7fvOEzfAn9tVquQU+wMEZyMlzls1MFsb
mybFu589iMFPRjavnRjxmn2IdpFhXGsuXnH741DyGBqvnvm0ubLr2jUg6u/QgeXh
0PuLcZMYtpC/964cvCDSzSDSSa/2i9qy8GAfvT8rh7Zk7aaxiSnZgmP752JSKROZ
DUnfwRakEac4aIx5k8f3tUE3JQ+hJ9MJzJ6alTbCkc1Zt/zKGekL+6y8OSn1SzcP
6hzpIEGIfJgIUISzBAQs2Zsxg1a9VP3hrbZBdm6TI35tLVR4Aq+eDRixFFF7O0ri
g7Qv1/07AVey4NP0CV5qDwVSGE7vFvuNAYAvCYivQL/P80ZWDv+PaTx6hbnySKCE
+v4tfsnjLIYk2KPIQqJ1cl6XC+7udzpPS2GFi0Z0LWpuFzl7sMYu/QrcYUtmO+vr
u/cBry3mHEMPhxihH1u7HzYWaanMpSIVVrgdBxf1g6CmxH/L7GzC+zRxrms3lVuy
XyjZQ7hb9q8A3bFctNfGBQqiQtT+u8QfrQ36yDktCCzOWtpc7tc9DaX1mtdsU1Wu
46sJg3TojH1qlY1ZQTM6f+mLCwHGREPRalGndNQ6owwvLsvndTB17uj2BglPbMc4
wF/S0txbjMVNHQLXC+ILum82mCo5wyshJN5do3yvD72qIzGjycj5IOI2V4XJ2taU
5OSB07zP7Rnt6eB/AIO9CGoukVRhxTgkZ6pW0Lw4oRSJb4tZq+plDxuNLA418lxm
/fcMv1H0nFrcWwrtN7h9STWbu2Y9q8NWCEs9lqyvK7q7cxOb6jk5CgmVu+Lzk4xe
qZpVs4jkeLz3cHDZyNmhqTXR/2H7yjxp2OC/cMvPy16hHwJFwL92SIw0xIEAGbj2
rV1y7Pf6RgJNTmSzrWty5vWb4eX6PGkNmP/mXPd3oXMEyqEThVk31/Lsd9DynNwh
4m1o8RY+/pgunPoQpiStE5mpnKan+epyrJaigQLkIDgg5E9LPPbMmFoAWxSPzfhN
n/a/u/+TmktTgW3tUDPGgFsS+EsnEAyI3K2Lgznv1yEs6vbwPpbR5EjlgiBdaqKU
61IPbqXdjoPDoOEUQh+A2UFe6OQSRFwYzBrhDASkJhV/aUwcfiC18c0DokLMBqnE
qPnN4M2GPnJcnVbtQqnEm1yIBDmSjPfEmuvd/z2eTSHT23PM1aRHW47FS5NevCKa
VaOFXwfLpQQqFah/SCu/C3iZPRdza5vRszs7Nqk49WWsBAhJQjJ/t4vxVpQGE8QF
X1Zg+V9EouOEE0ekFeg+BT1NIbPvILgruB4NnJSID287aoVi6M34HbFbeHE4HOVN
b1ZnqRBOcdm3Ym6Q0sE91rcPMr3Ii9gCeGVrECjkj6DQAcRyFC35bZ/aIO7/MPWF
Ma2mgM7EGIYNsOib9UhZYME1J6eeeyQzWVl2Q/4YPsO+tIBIA5t2B3yA1Tstukhr
T870b7fBe9no2fONKkj8GusYNk46wU8/EmUflLCdFOq6fN2mbEdL+HqQna+E9uUb
vkpRRo3VREZs49dAPskVq5WIVBzifgMCb10T3eCVet5KLGClzOYpvn0anbkfb4LM
CUQ2WEkQpsZftQSGsiGEtg/COx0O0tCUq59RNcOsOvPh1kcakMPzwwtOQ9WgJo7V
IF+NsPFtCZ76O/rAtCzZN2YfCkko6ZbuG++Aqbe3HXyrcbNX0vkXf45nXFC8PI2c
waSLBF0Jqm5/sFbuBrDSs05Ib4oorsbPx+pZvjy4uS7Z4vFqJLZOamq8ITcTgQ6t
Jz2eLuErNqB3E7bXjOHUwh80Pig4PvZ1rMgghGuOG+/K8E2KHxyuX2S+bC5UcaJi
NTV6WiFSF+R3bGzU8qBRCMnYK0TbOR3Zi3mQ6mQvQzsqOkIV735DqbcZJkofUftn
PV3FEBJZmDSXYW6u6xxTI2r6JudBMgxiyRK13bjzLAR2JougAt3c1ohXN/iGTjMQ
EuTXKy9BBDMul4qSNiyCz+rBm1ARrLVU7OydSKOJU9OmhcxLcbi4gHvn2h8S38tN
4VqWWpgNPILHBRXoNHuuZLiW2qXt5KOdbl8u0AbYn9PNUB8voxD6r/TBO9XZIwZM
eCSzjkw2yeHpyW65t+nKZjPUtCMyjqGQBfXtlem/waPe8hD0Pqn06yG4c0Yrgi9s
nXy8dZaDf6QdpSeNBVdoGmKopjiivbgBracJ8A6zq3nDe4cHFO8JcAsG8+RlufRl
TwI77Lyh/FGSFrgxFTV88EFgI1egs8lLv6E9pB0EQNusSWkTRxgXI9vtJoPIQ24g
uoqTTOWcyZgIbFb/ZkUESV0hq1w6/lb7ZpspmzPUsJt1MjmU+TU2XMQOM34Al/jp
zF07Kn31c+ZAyC6dse/AfbcMDAF+uKGcXcMsjlWU8VJ/O5Y81uXKD0xrOX3OvlcK
M7kc04x8VTRYvBeUG6lPQCzOylRE4U48sGHPEVJ/2Oo3nQ97S44fs3XYkdquN35q
X/0TxHkIoCxND+5pSgU2S+ZcjJ+d6L6JPxUV5fISJDB2PUl7jw7OGAkX8dZljarA
6rl2b1OYE5RJq4HV85N4lWgUfk6cFzR+FaqsmNiQGYF1wnhbvEAK/dnLhwfWL5Gy
0snrprl+kEg/Oq4E1knVqsljWPqsEqaQHsduNEUrc6X5mKkmCVfHPzykZNGCFZbK
DyNvPbo/0YWlIawSfY3jWKr5GaObiuk3G7r07+pR19gRqhuOhR8iFKBj1tlS/tMr
yFvs3aSTaorPAhJfpsM4FpXT2zRN7lPig9mdNMnGZ/Ft6DBRb1bnD58OFKmmMLtQ
`protect END_PROTECTED
