`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5P93dS5yZZh/u0OTelRYXciDOO3e+HJOxSIwkTX+tL2JKIRjYdy75RiKfaRhZRF8
8qx5Eji1DXmAKOMoqtlTgSrCwUmXrS4NsFNP+T48Ez70AevkX6Q/PlFC1ZMGbItq
7E6ZUnyb2XpCYirAZdL/frijkE6gYfg458R4Apl0X6JqjPi0breHHIin9eGB6OSw
qdxS8XK+UhKQokUf8XljLH+IglJPdSCQ4p5e+y5yL17XdVfS9EpqZiR5KZG5uGNa
/QDT8LQCk7HPlMwoEVeF4Co/nh8SfH73VgRrB+2+n/fS6B0xUijM0UO4chMkHaAs
GVJ+Xy/E/h9hUqv8b8IRcm0Ge3794DdUgH3iAXHOg3D7092vbgzEO+Org9rhWo/b
aWVOmuYCYRDsEtpwACqSTfkQfK2+7ES4ySuEaQF1/EFbj/lJD0PWiwZGjZF0BAp3
YNRP2Rf5RUlvrEVR1M1fARVXXcclAELy4DqmtunhgwmGz69DiOb9Z3gguYuB2tTB
piPizEXetmY9UhyFOo12JVzNlFjV7Bl4+sawDD6sCEaZR2vM2NGAAUH9INdcDfFZ
bVAWULD6Hc0LA1ulmli9RPkxqRiL7jwLZbQq6kTGaXisSrcEe4r1Vrjf+p/ri+c8
BUPGhcDdYMstjfSjUqEWlq4BEcu6WQN84B+L8bnJLs+bZJB1qB3n7QQi/ltypUej
fOwSvweXHAKRKdSnRbBO4ogH3zl/3WTS8qQFEEaZIkX8nybtwL2u35OaSlXXjg1e
eqRv/ajP0rRrJdB1AkILbpfmrGExiwIYo+Vo9436pQN6mOe8bD9swRUxpChK0gVB
6tgbRW7/ks/mwRFl105FSFVH+lXBGvVhuvypWB2KMUisjCJve1EKsXdxfrKhFc5A
/B9f5+H/+scGHlYayIsRIWUpMhJWub+S9/ZK/tSTjTW/Isito+Ju21GBznJT9dut
UeoTj9awZBbXG/EKHkKJSItvSblL6BMwiAsFB8RVor/dlxX4WCVgykoA2uvkxRy/
1bcIMH2IH/LgkAL7U70fAC25m6UethMiYqt/U2WGlk9JHd6zik6TCTZ/ZqL4N9DH
OToTCS+E1xRojGGEIotlSYSCvVHIvqdhekkqnQ7HdUSWTgO+G2ueFsNdEtakJJME
X1nBFHK1uAWVGvNeFmxjhnWW+LZd17os6r8lEmoMVPwX3z2Xr+VhyqrxtqiUXf1m
Hu5SbA5N3OCZkWLDGGhx6Y6NQzeLncpnqtAD3P8Xylam010OXc5Tb5nrN2blvoii
3CJ2iJwWHVvjNcxbDiQCpJ1MCiQemSrbGJy25GOZvqh5tcnA+nzEfdUxQEANP6dS
bSVEBKNhfOA9d8oRudl//A==
`protect END_PROTECTED
