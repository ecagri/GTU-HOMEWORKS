`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q9+e3m9lEMxRyg7QwXlAIhfCPh0VupPFs/NdRrJjf5zKYe/FLQnIGxeZaRCCvSl3
DhSJmv6Ub8FrfdpY9YDMO9DCVL8slel6UgocR8z3nGBId/QSUkwUf2Ue8IPr0lvN
XhLEjTXCJvnfv0MQQ+ss5FNjE72nyq35v31Dw9l0WZm4uSAmcno/AkiG8NSjuxHn
RSaOvz075Icbr8AmaxZ/A9UQGXCq++8AMEWidC3uqe9eweBu6MM+Tl6MjtFUuM7D
yHJX19feqIA4SscCUGr6NMtEYNoTrk0WP6fYP7TSzJgBmcnVwR1iJP42KrsqWl5U
+miEjFLkx9K1FnHa5LRhaKODL0yznX2VRvKWoo210g//H56U+iwNWtiCvJiocI/c
crlKvzqP4JHHGXLHW9RgUckgh79g2NAI67Qfi9ZgFb64bUECyFS9pLcA05IhEapj
f3eG/Q/jyDmbbIzxDM00hCZve2cdG/Nav6F/EgrLQPuksPQ7oOxDDrDc94wgg0w9
/UJD6oTAkrPawJrqnZtGCcsf8qtQ2Hrvr5AzM66vhaBHQbYCIq+KNQ10GoaaJfW0
`protect END_PROTECTED
