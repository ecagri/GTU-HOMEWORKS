`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zyFq1j3AwGSyVwpeTuni3ULsRTwit6uRipQVELbbthzzQuWe3i4RP+fCGyFdSWBa
cxTnrSKQhPP9YQ5RMl4NkZ6e61YTsPXRWBJUKBVrWrbvXne45LgsJeenvRoQXm+5
bhSYHGyl3mMbwC9wo6VQE3CR6/wqQ4vAIAf/DZtj79z6gwayRBlUSpEckEg3Jm9+
WMujI5eX5jRWI2QGEs9tkl7Yjj09Q8AXxuMlW5PUC/vof/t/aeyMWZ93enBTXWjH
WsxlH4lO/Seu9w8Sojge/x3OfmAS4ob5XL2whNExiEFhbfYU0GT/0Bkbd61oShGX
hgB9hY8jlG2coTiAYoxFFrbSfHgS1W9I267m/soFkBBDIhs9JjCgXB0BV84p2Upp
sDdZ0cR9RfNAGJlMcm43frfdRM3q94SM0BkOfs09s1lkMBji6DstKUSbsOvQdKmg
frNPd/9sem+TbM4pMRzugCTb/+T69nHNmHz6OllzpBxHov+iW/b1+upUpB5q2QnH
mqcKegz+o9401okxGhb8TyqwWGMny0zTxE2nSnSGpMfzengCpTdfgljNnVQjTvgS
v/qP2Qp4MuIsFbMScm7isPftjoKthesl7LNkSqY329YdRFPVTy+67RfjH3ydinn/
LFcVVEq7l2jfcMEsHxWO+9Y3ygtMZArTPqOYABg3KPFvEyHSxgSJwlob7tK6TKwO
oTEQkFIZbP79WgH0/jsQ2eFzdOnze8S8RXM6oI2q6XSbxZ7BmDwa220b4kxDQxXy
azNgE6uDH54T81u/NjjRflh174aW63WnwuVJGiTzjMsnj93uH+y7lOAX5FCcdMf/
pyq8JYxrOxKZUqFVIVE5UWzYjM9OueWEtlkyX2fuly2ukhbLpm2sExk5HsubtBFh
IUrLJ9rlwVNzD14m8atcmLIONRcdJ6kkp/8jYACMjxPqxbjviVBtcehKhuM8q81D
J2x9EDpx8zLRURGr59f7XYk4KODMC+RwH7wiw2DlcGcX9VQWFscunUB7RQGu1wkv
QG5NL+Cbb9euhbLa6p0GaV1Iu8kRJzq24NFXAK0yfxqIoW6r/DfKlEvq2tvQv8Jv
gzYQs26LWsnh4yrdfAC1N0ZVz4wGKorkSe5HOTAr+FjZehk3p2r/GqdgAB0laBpg
Onzcl1AimNT+3gmYmMHY/jjqqNP+Q6qHVgZMIf7kV/P3b0Pu15o8OrKP+kZ794A+
Txpd0SchZAVk7qzOuyzH997k0lPs8egJFRl+Ks2j3pSVseMXFNVUC4dSdCCEZS/Z
3AvLFgM1RzQ90nlGweOurJSYL0p5Z55CvdfTKvrGcSSp1Rx5Ic3wsTi1TKpG0SQk
HKbOXHZKVb5QHF2Se3Z1000GSR5JeNLuYk0eUOUUgN6YkPEV9hc0sde3rmXUAdEr
uqZADoDPs9jWpWgnPFheEsvn74yUTRvgtjl+uZ91VY9zemIPMg0akojjCy+1sRZl
+NFM31ohbzC1HWsyQ5Ci8sODnoOaXxRZDxXEuDvC67mRuYLizHp0Ea0BbSgVyumd
UeCWffz+RplTixsUnZnViVLVYlc520ZwP8INaBK5qvs1TiJk0gO3q7fcs1Unot0g
Q1lPnRlUQ/3zZlvQIQv9EIsGBwzzWL//oeQu2I2Eci/OQrehAUpySxUA/e6ZTHjD
GxQmANf7HoMvfRFSXRQh3LS4h6qKhTczocfojWHx9ptD6XuX9J5NueOMws/RAXbQ
vSA4Me5la6CEXcKrlcMpO03qIhCpEYdnRiV1VZGzDGmogGY7MNNfFPmyPviEwy7G
1lCGqlVSS/OU1VfkigXdqdhpK5sNwgSeCr/vlNobF53NLiQHisGd6HO8bGA4uYmC
xahnCkm3od9owKUPNOLO5x83mWx7ejzZeZrkI6D1N1N6HVDl/6W7j5osNxhIIYFf
Oj3H+W8ZFlBphpI0WA0PKeAV0P/E9CfUPWOZ1fG1yoLVooLoRHQYTpXApqQCB3sT
RYRE0fLidKuXtA2MyrURPy1QAOBjUKNWlxdVZwa1DBaeIQwH1aBr7l4r5PHVsQQQ
BNrU3/Ow5MucC7xH7+ovYV7wxBwdH5aQhN2z9XuymyutiwcEtyXr4A0SvX31ERAh
IHEEdIsT0nJH5b/l+sBZ7gAxoDInkGYx05xVG7LZ+bHGwZ2ckc8DgP90M5uSDhTr
p6HtZa+4uSDvYWOTZBr0RLuM5O/vycRNL3tlGTM7PUGoo+JgwFKOA+D2awB6fvwa
jliBT2AP1SLlVQYBMvH9MW6EKifI7eC4cz6UMvypxpDSfUbOQd05UTI6sWpRk+8r
f/GlFmRktyTuOiU6W5yV9JDlbEEA0/Ly0R0Ft/vIc6DY9LGjSF1n1UIf0GMioLNl
Wk8bc7BpKBrt7pX/RJlB8YWeX7dU9HQggQLyi1AeJZWKzRJiKNpV7c3tSs9x7XYJ
03Gs4K5V9F8pwG64JYRga3HBFkhCvayS/7HDPwfOFMgY2Pzby/x5en4FIZG/glHK
PFPvpEbsHO8Ae+5q++TBZv1S9beNnN7bkF9KcZexCu1hzx4rnxB9YY6I7KGc+mfV
Mfb5pPOJRVDW0OprKm47bEZHy+B3H2iLt7I92W26YEHD4xEoiWrtMHwhr0k7FeRh
N73dqCMvZqljYvX3q0rNrx0Lz1gVsqmX+vLigTYdgHvjodAb1rx8eoxFwB4VIi46
2z+7EQHlmjFeK5tK1KpdRVOBr/xGH5438vvfoiP72pnr9P5LAekbr9UCKMjYQ8bb
0PXCefenyZzlmiEZvs7Pq4ZDI29eBjLk4k5M4g12CQmD1fTy6nT6lCwKn5XwNzGG
Igg4tyg7zvI65S/f/pWqB+0dKLEho7qgq61gQSBEroDs4bq5mKk1hmYaoAALmIlS
43HqwtgO8/gxpmhat6Lq6GXaiB7LRLbQXeN2WoFKkCG6rp4HcKf/c9SR24sd6+n5
0K2jVl4MVW1Wm1raEhuctArTJdU5sH419SXDXxV4bcHQKazjNL4L4jm55LIN5C5e
RjbXTTHQcFNJqvtjMQXVCPrwsjUSYFPFvL9Q2wNoHHpX1S4puMtcNgJi1KM+OA1r
u2Z/OFkXSd9H4jRjvzSfz+lH2k9DZL2qTT/uY7aAeo33q9+eRrOIV74TnwTH6cTN
c7ab7KZ0s9Ze2j7eT//9pKmFT8a6VoTDv9nW6z5X1H78nkkw7MH0A4nxKxG95C6S
2KL0gDazsHIVwfmbaJvSF/JqPbjcJgrmJ35saIYQHVKyG91L7uROQZ7zSTv9Yoej
fzdgoa5VfbIcIR81naUs81CbgjMF1DxntB9GCCTU3Kha9OUgNT4bzuXh3U8m7jWF
xPo6gKjaCBnE6AZtfQ9xQTHOBRm0NyRh10dFrG9xF7MCM+6CiSl5cq+tTURarR4l
INKRGnb5xQSbSZd0+FheM/K34tOdfxIrHYrGCsPv5kklVIYEPkkICv5LzYLgGsG5
Pq7VVAbiesNrM5s8+KPj0kky42Mqzydm7pUfLRkCIEMqChWt9GrV6sTmGJgv3X63
aBdfndkdbzJbQPUiOHUwItMRYe4t7aTbxEfOt24say6TO6X2n02xPrOSji8Vcqkz
jlu3NADFuiB2yX6BhPuMsgRoO2ACFQkm7enSr5UBzIg=
`protect END_PROTECTED
