`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a61RjXxe6JUwLrlvAjRtY/qARXYsswbThwVKWR/mU6e/0GWrVaqj30f4zh21LmLy
u6mZmx9m05GeI7qHB00in/8e9OyJ3fPiRSrt4aGbgJe3dJc+PXCcVfv2HHqfj/zz
iEYTSjne6/Buj33L03N0EO43K+xD/PXmaBXjUpzXfLKC5nsTEPUvkiUOO6/SBtTx
TtK3wg1fgn+U9GExRca4w6GnTWGCTkgkvSRR2PWzaFb9Sd+FwzBk3Sc0GwPSg4Ag
8AJUwgrnl0a13f8JfZktNQa8UfqWJBQquqAMOEiBr0OQCFVldM3VxjTzPizsl9vR
9W2ozH22HvuVgr8RA7/XnKq5ZHB8kVpD37mC+ipOYp2JybQSUS7J/sI1nLAhXSGs
GbvNYUmEmmhr3ZLdz2pJcEFUlIM0SFYAYqpLW7uDFSeUKkbeCWbPxe0cjkDNVav7
owXzO69nrqljDlA4ydxEvHUYP2mNfs62JGyzGX70kh9CVrFgpYV8VsBewaxVcAms
TMbhosyOD6wC294CsDrLEblTt7haSkxFucyZxlw30olmDA4Oo8w7f/jM6N8JXOXI
0szmCKj6e1HzLGcL5z31zpvFukeqqJm/AL8Tm7h7buZ5k/NsKlqegukindQ6EKUX
bzA2TQeSgtto7CcabKpOfj7U0xFjB15qhZBS/Zam8EO2i75GbCE3FP3/jOYFaUoJ
U5pf3Lmq6dG3DdzYxmfDP70XrmuZvSrhu/Xc22rI2s9ZPRM5v1fuF33fooIUf6T4
g/4ZT/mFhhOUGDK9fBaPBHuJVBPHscReKdCBgLOfPQSrlWUEIVOGa8rin2fo0Fyh
s+Pz2ONepSQDc0iNgysfzB8rueoy2Aa5r+HtEHoEiL7eR02hoH+fSqdRXHcSzAKV
/8pEl+s7ueTlemp8muUP10fkqlEP8hfM8TjSDzM0dKT6H1mRlKrNOrOlJrBciupr
B+6AZ7wcpBoFNOtKQzYJjW55xP9KpAFTF9CNH/2OdMhChwjS6OIyTa2up7hU2uvz
/RXEwyfSEXkvLLtfZdIhxABPMfw0S9sDnJVqhc4N3bGleVzHrhYWr6NWfOZRushw
9lWr2OutH9y5OxhBwAqAylF4+jia6cyH5ZeYqWRuUI1x0+RPe61oOS3xSmgLp7wJ
I2GsgAXdqiayUEnfyLNL92YNb13AUInNAAiLvi3dsjWSskvR4iRZvosPodfcJemI
ekrzewlRXRwk9RiUm/I1TE5q2KB6ZWLBMxSxWLxh73mZ+9+B9XPL/7SrN2mBjCQF
1mlkI+y+2nbJd3LfB+95T8EVpY8qO9r6rX60wnQYkfAXJV/gw4wo8D8/lGxhl+Qz
7DZd+FizCAp1Asozw9JfpbFiGfnl+h56LEsXAtaMHmFbpHt2XlqU0cdkF5JR5AiQ
IQq3hfhQcvMSdnaHnk8nGJqZ6SKcsTaIpmh6n1JzIIKx5dGarJpdXa7cF5C5CaMg
B1cunlYtgxwK8CIz8LitDDYi9uDKM91HaWtCj3hu+zWC/ZrQYBx3NqHcBoi87K/F
UTyE9jY8iw/Q+/CFTueGUFWw9resoeBIZZ3IBqJ5p6N856oUPdeWAze2wzjb38lm
GyyLVNT/bsuOs8DeCWy2j8bnvGv8MlVanN9O/VAd6yWPMVXP12+/AV0HXEgHR9WS
8l3RlOGj5X9m7brwCes7MDpuPyMit1kUANoMGi6ukLM9S99YHK+oUO1/Z6jfvaba
w0pVG6AR4YsqlWhIHjDyPySX5buIgP6I520fIkjNgCIZKd5lSYSdjLp4fVtp5MjF
hSGHtvsYX3xsLkDGsmDFbzVOGCaNfLxO/NoaWw0R8UuC0aoyPBrh561D1HGv0AWa
`protect END_PROTECTED
