`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4JKjhkKqhT154/AeDP11F1IEGV8wsZ6a3FHl14bCc6Aqx/BNsYIbcuIKLsxPoqPO
7k1NJYv6MK69TlReE6c/XrfLVSghf821vgpHApRHHgTO7INCrBi1cBiru5pKbkg8
bQNIbxWuON4HpmE7t8MwsgJs0G346p+tG5zdP05vZN+iETsxnct/aoT1cU1jzQdB
1hDs0WeHR6stb1vy3mWZp2Yk2d6zip9P1pWZ6odzqi0+yTOMariIV708t3PAh5uM
ih7sYSoIFcQk1sGkv4UgMuBTI/hQcEopuRXGwZtdXo/qHOyscndhn9nZqYwfTVx1
8zsAL04X4vIerkf335K9A15zUKwAFVTW1Y+DWdVzyviM0YA/Lz8fDPkRvEDaDJvj
npHZGKoZDP5v08G6RrWqFKosV6WtSWGyiLC+/J2ncOkTgAOqFm5iCsFsdxS6CRyb
vxrybIgrjDFbG7Jun6ElaRr7xPRirhoytwZpZea5KTG3pDUyBQKJD4iAEjl3jcvq
OciGEXqdNaA/mjqU5ZPHCeV+0Nuf5VmtVQV0QALcOwXZW+7U9iLPlaQTRyawG3f+
tP3kYdMFrsXCPZHG6FX5SbwHv6w76RtmOEnpBekLTZABudO5o9T5FXCLk1q3SuSD
p68v5iU8ubNNT9m0Ty4UmAsclDUSd3gQJ/1Pe/6eePtU9pZH8AFA8YgfQcIzqjeW
cWwAruYgD4nRnNyzONcagULMqulUQ1q/vSQWbaktkQipZR8jf/r8YN1Dmz1DHy1e
D2Q+5VywRTPHS2tzj7V5PNC0BmderpcZyI6HvxKZ3uhhz3jwyVRTMJ3D6P7VFWK8
RZoLZPdP5AQ/NJ5bNGKr5fAkzMQ0QATWzzeIxcGR6LEK/WCrdKuvhsIccKKQEKKx
N6G5sJNUT+RWZv56lovJRiEyTGKogRLIWFdVTgXRAnQ4fQU5H+e1I5t58VY7csUu
bO1CCMgkJr2IE9b7zwtDvQElBVEkgEA+6Qr4YCkwWnGePTBAz4yO8JWjXwzmyLFM
3BMuVmXspi3/RuSru8dmroSkEZgw1LIrEN0Ja3be4usFvgdPlHHA4Xk6rKbFamaJ
x7ykmGFKB6sEoR1Q04EwGgHBbM0juET1G5NU21H9xDEmaOsiiFmTJfV6+UgzDPjN
51pqFJ9RNxG2acEVhVd3H7YPz+/2vuNfCOi3GzS1US5E4wyXQeAzg0TZMn0P8+8c
NGv1/pKx/GChDLtycdAXFlxRr4wZQrssDJOuN467jPoAGJXv9AuvArekYvwrGq2Y
eebTcHRJPO1Pmhp2MVcVLXnc14aQuAZ8tIgVBuI0WEVowzwVRDR6Z+qXIndVqO1l
QxZD2BXfraM6gP68bvXSjHlokvysE7ppFwTMqXxmlgYwxBSx9Zs860gRzObNpcdc
NxIIkGkzXw134AD0H7C8zxXzmFgDYKE0nMN25OWK3/9hGSLdqsNzL6VqPdKfTj+y
ju1EwZv4J/GiK2ntAxEL1Dn+TKOvIZ79ueuGC/RBlESGI+XFa0emxv/8pZAtnWIk
15zrGtmyGBIAmnJ/Oz2PKQDMFOpig28CIrf7LfKyqn58eVv02QQGxK0X4LksHcGh
i8SHi1TUDaGTopw/zifGh4xh7njfN3U7t3RxvDGuiWtszSQv9YDMLGASWDtqfDRh
X+E2hxF61XhrWjEZVzao8R9n4qju/iMJww68O4Otv37gYk0P6fQpT3alDpYXtsY+
Mpy7S0+hWylwt+WBYazbRM2dbn4pz/iBIv59ANnTZVMitOc3AZ6dy4Tl50zdDwxJ
+RCgsjcHymUtp1lAFsJLM/7XIcjZykZo4AQ7f5s+VEnHs02apByInHHv/Vw4pEvj
LCgyn17GZ6XOCySnri7xMYOm+Y/JPijjU9e8bNnrXeLx1pvCyf/9NxcwQ3fvvStG
yu9dAMwUea4Q5fe0thfjFViWtvW77w4AEyyREfaxN8UHmRt8HPemgmMp3xkNUHr2
taocGoy1okSOS+kkNx/diuFGBnqZT5piWhonnZf1HzMGI/wsgRI+7GH1/uBRJvuD
Qc3/fqAdQpLpNixCKt3sBrWebPzvCcqmp9g5T3+GIRie1L0P397hum57tVn5/cPY
Rj/VjBQE3qoa/jIzngDddQ==
`protect END_PROTECTED
