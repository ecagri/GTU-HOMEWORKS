`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CYnTqXCv2aGGLRtiETSQM7SvRyrxhwliqefNlpo4EmB8TJuMG6+pkGoHOINu3/al
QXEa7NjdnUiI0dEDLKVs3glG7pWsJrvGkD6H54RKhWro0GO+VCgFzEIuVgif2t/r
IVSLm79ipvNFdxWNXMPRgvL5PhPTWyn2pyPlKOu55sj/hGFIXSh75CaXBCmCV1hA
N1n9Jzr37ntoTgTAl9VN1GpAVfe7ilWqrlPqQ8UIVLHasxBebwBQ3MtqW+EsepGR
bhhrfTw/hZl2DxXbMd4eVBukqnHAfNlNujAGNmCG1k+05JrPB5cYrV+IKs3pl4ur
NxtrCJEICSAsRjr7JoQzKVd4eepPNtwvMDfqz11UxRnMqPRh7UBWA1kVhvjEbQFj
+MRa8nZ58mRneguugGhrI9S3Ca1fi+ett+1wy7H+VRcRNico71lpncqYFHPevqj6
mt2RF8AjqZG0ogs8BtCiwGo6quKoi1LMuhAHJP7IT8BhmAkk0oKaMhuSQOlOr69T
F+hZe+xqDwdPmciaUVRfzNFazeFpCMscu9fU9mMRmyWneYuWFyiSTvYdMXT+R7du
Gwx9LvnmgLOWaTpxggQelQVglZVd9cvtt5eX0H6T19F4y8Wil7LBxOOwnr9hm/PX
H6tanhQyY6l2sRUMujcXqIiX873uFE2CGvG0PClS1Y6XoOcdEtOBxVAKF/cTDfwS
8bkHvZAulzJK+J8+eLLMNWzk3y3ffJaPMD8QJNwnSKghuZ+EA76epDnbOgTb9iEg
CRc4/HIS1+cCvS5HnIZradQOn9EDbFnakTuJNkbXSalVkgQxhKa35XpAhodLY56s
wH3+DyBy27NeUGvGcO7AQUSkPijjt7Jcw10Xiqz4P47CJz+aVHg+pCsL8GD7lzkB
Q+23LMCS46NaB22syNQtSg1ReB30NdUdglt03LNUgzMiLT1j2A2UYFjwHIq9nRel
mgYHIHRN6UgOZvwicBSKBmT5litakHCJjTHp0dYwVs44fmCTATsiFhe/LDXBS3RH
+VliR2H6HbXTJb7RmMektrqd9oLUsCpniytAxoF9j6r3vEVDLBGBgJKuvelRcG7L
2ZH4aAdO6yWM0GIfC9oiADeKiAmZvCxp43BTpo+tJtUfO4dHWWx4MXD1KWYzrZnv
+vCHxARbUJ3LNyHNjPIG0xqR9yEWEWH0hSn0yWBdIt4WRO+IgqHQyqiM/OQQPIA2
IZXgmfbaHvrCxOP3D+FUWYN4byfKWcTv/0vsLFlAqv/fgo96Zsu6XIvv7m9DgiB7
6pBlW9EQlUwhdOpV9cL2YhJNPS3JwxyAZnTz0UH6KeV/IYnInQMwGw208CaNq9NB
kFH+NTLTihQW3IfZ5mI9o3bYk8D7eEpyXme0DmvLwWVZsB8PmNMoiMA4+RDK3VPk
Mp31PK+wfn7toTPCcpr6Kftwm+2HSo537H6lOjp7hEJRlSFecK+Lbo046QBuZG96
tXolNgWSR8wNtzRriOunyFmPapQ3Ann1r3rrd01nM0DRQJnhrc4oHWpWHTG+E+JU
3ZgSwHi5XUnZDlMSVpkmgGQDm0iSnuVu5zTz1Cs7pM3tx+H8MbIYiMK5wxK6NktU
dElcZ/keJcT/oT+zbDbolgrY7+x41oLcRORVvYT4BbsCqNo8XFRyc/2zflO88BKO
0jQ6PjAlQAZyMXbeLKg//7UIptsRceSWvoaen+Wshg0ECUuBC1WGg6jdzv5XSMVC
DDIGjQ1Og8QjMrewuhIt8MtClnaW//q1m64x56JOBIwI5deXHUIyoTlu/rjtSxZC
L1sD1B5IPOEHxAy2yAqLBhSlB4UhOFAIAI28+omEcJ/yeS4t4ztwn4pFESQJvKVK
UB3irXDqpIxKLn59sz1cik25kMyrXwGPlt+/IcjKYEkL0I2M8OVYg3KJybgt+f1D
lhpAJAyV1aXdeZZRGBW9uhO7acVPnWtCztC1Yy3djZUiN9mOlqTxhisgl5CcpFf3
5jySexvexYdMs4g234yYBs84LZg1Z1Ml2go8WZwMQEBH1mHnRlAKxjgCQaQDaQxg
HHD8vPfVeIOQ29IhV+xcu2KLjx59XMgOWRPCDK3hkv5bs53dEWa/4FGNaR0Tv7Cr
q+eMp4bjIUBpF8PPwFsWAQF7NiTRE+93zKcsBgITRr8jaXD+bPOnDLulgArWjePg
KmAIOnCtkLmfAJeYm81jo9PYkVKlV5dCKnREdWcqbCEZhCp1Dq4e5i7nRNpHli8O
hBRy77/sVU6FXKoikuW1irYd6WXosCS7iEueNMdc5J7Uu/Z2DzrCNbdRgFw72m8l
8x4idwCyJvHTCtucjUKAMxoHWwf3t9H73x67dvrxO9wnTzc0H4o0+iXwWnAUrxiF
lylqi5PqCWxWSFhz9HgaGloSZjD4MopGMaZHpuXJbc/v50HP9nSKqEXrh5nyaNaK
m7N9u9bQwcswb21LqzXalg6mAnywZoiiEK5C2B794lejQdGbVHudDwdkxUWPj5Sj
OWPEvCn7qsaabX2uXwgaKQdTdxcx9FAdof7qdpPXj7Y=
`protect END_PROTECTED
