`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C/8fUEuCm15jUbyrG5kp9c/IqoXneVF22qnhN5AjZaVgNU0lmEQ8RvfBZsFIKiy0
k528UcyGWAxI9Imxez3zdQ7F2c6tjIl8AGcXPKTrDsCmO/ODBnXdXBjMkJJ6lbTp
xFw/P3dbtC5gQQ5WCU6SMhGNYyH3OtYqmiUyxpRtCZ/KKPhbxv9UwusHj9VAcvWH
IM2n8OWcABXsKhqmwcaOfbdFFOvzZ8o+0d2SRwY4SOoTtltqjRCeTLZvvlPRuOu0
AT6xA6yfM+r2wjDvu3R/PjapuOC0NGV3WQJ/3YkJwf0iheNfHUTT7R38rWO0H+EP
Yimwcw8yF9Xf5y6utLINpSs2WFAt39qu8V2v4M/0twUil9BtvIMiVnQ2MvyXIPm3
02kNStQ9myJcFlZ2iqSK7u1GhZwlvI6cm7TjEr7DKQ93hUuYTYpIa7uZqou0JVKz
`protect END_PROTECTED
