`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0oBo8qONxiB8+CE6Hw4wYu0U78qQ7Z0nFNcTYKXZYC+ts3/Bl1m4fLgAcC09FZYw
FufX5UksKl07+XedRBdWJxdTC9Wbc/dyEuzaYNy84j965Ef2BDs1OUSRGHWZ+Di7
MRlyrgHVY5fYCGHmFy6BFWaqUyM1HVXIS5H6Tk6LANluTT+2lrlR+Rv9zB9ARxLn
DwEoi28SnfPx3bN1gdPqNOhOXQohQVcS0p1lp45afVqkKUQyKOWfAjIZmy0e/lU/
vj6Iyr84p8mRIjmV6eoQB2kTRbgIukFYfG6lbGf9O3TYeFNwmebUY+hwGx+Q/an7
WdJTm75fwryiWlnZopBuJ3i57gwfNCYKUrm1EwBce7Ojhee4GwrCWQ2g3q91uRyu
xufYuAfF4ZXg9epT9dV0q3v8rv9jDfO839UZ5Il0jy+X+kav9mOt1hcL9VU1miEh
4mb6psSwC4PzvMUTazvxCrAMiLrg8f6e8BVgHRf/G8hwZ5zS/jgPsG3U2XskbYx2
SnP2O0voB5oc20LalhzEaG2N80I8S7dpCR9bMeClc/Pg1Fw8SkCsKzgFXVPtP7fz
fDx9Y9QQ1IVx6TgkVBrWMbrJqdAJOoSdkQK8FFHcan8EQx1/+CfeBg/7E9nDLxxK
rUEF4P9SZEo5eekArzA7ysvXwsaguR//019qiDPW92ip7qjO5gjDaZC6BfFt+cKO
yD+R1WQ7gcC3/MhxyjDI2R5UJ34XR8xPI4ceDFE0QwxUyJhnzCGWNFv6nMRnTkqB
O9vkHhr6NJZjfY3f9MP8VLNIxZjJKcaR8FX7LXJYd7O9iWQ9ONdUg+AMKQSWYAzy
XQgDxyFiTgU/FnlFcgzReCnwwsxD2BqW+qZhdsuRNu4=
`protect END_PROTECTED
