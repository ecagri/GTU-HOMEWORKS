`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l+LJrglPSJTWPe9L5Iz5wsvxJsqoI4Umgo7pD11yUQWV1pGDmxwfwuMGkZBD4UIb
h/EhtSusN6wSAMEUERl6cv74OwT1a3vrfnb2Ms3POstBkIxXZ7b6hcgY02a2E+aJ
aT7xDJ4mtAF193+f0B9f+o2J1YltuXH8tId6a7Pz6oYbFkfZYKoF0VSiyZPCnTIj
w1BdzYEoiV3rVTe8b+XWNd3FbKUfSSNxg/iQnPX4IFxRqotRboK05SxpR8EnXAs0
zZCistS100ilrG3AvyEsFN0G8YUW7fnBbVwGK1gW4rxaPM2mg3jiUUzQbZfjzIbB
ahqtG50LLx4pW05mrf6mjV9FXO+nnibaLfrcM+bUCmgqyrJ6GG8T992ByBGtTOwM
+4jQ8hDfX/8qEBkoGZW5dB3hrI2jsmoTolWkQNbP9ZWbRxjj8QRUHvDmHdfiqMmp
2FicS2FMTdGz9TfW4m10NAEsZEYk0aJNMgYJV9TwV7tBzksvnKsz9iZR9W3scGLs
LL/Ab7I/zsqqD7Uq3LIMGR+2ELu0YSuAknTazNuVSAjWM2Y9vi6KHjQWo/DqN06Q
A+EQKGA0L8Lt735Q+m4gELaGUXei/k/konhfds1u5oF8KGVCcp5eeehnL5xpUfnU
scllCcYgehjhFUKK2FuUyiL8Ee1hbFoIprxul6TYoeFAHM+I4dewPGpGpLNfXn79
Z9a7fpaXf6tsD42k7qYF6PSe7cHxsywZHi4C3ewp17GkHMVaBh3xcgCenhdO17w1
b0Fx5hBSDq3FeVGKJHZmouuv5PsFu4o25gMDXVtLLmN/v7n6DMzAgVqx1npGBGNN
BdqEek2yTrOeH1nbUryckC4E9a2+n8Hi26lqjWmDDTY9lQRE0psaAzkU1eWEFhHj
w7oP48NkV/5DvJXRqcQliF2xV0pIuwuhvseXDadE9NCiyurcSPZ+ooAxzgHjq8De
Q2ODjoZ4m0WF8S9tGngYK6kNWWv+hLs/fMSaBQT3ixmEaJJHrpZD4nPnH5ejkpA5
2GHS8zojNxGkAPnk41JkpJX3YwE3h5NjjcHTMcmOVGeZKbTD+vFjIBwnAT0BOe4A
8mceWeNJrgZzDnB3wYq27tg361MjQXmmbXtKDO1k9Ojjp1D1OQuk2WAITTmsFeGk
aspSgmXxXBgR1EfXZglzL8EQeJ2LMbwGinH5aj1dJ7ciOoF00kOTjr5lW3BvQQ1z
uetojDXRhWO4hymoiYHqTcIt6jQWUnFc2VSVBZsMdCbQbKf3My6WzdzHcJcYAvAd
4RricbufIIBAyzSYIVdRINXHOzMFZISWWK5NuVedYDgUxYmxaS9tmBPENrBMsO9n
QacofpRhpiH4mJOs5UD0fStj2OYSe9YHdzAT3yBdPEWgsCwNNT+C9rD/5S4FbqIe
CkUZd2/m4hJVTr84fjKRDlemS7jaCKWdUfYi12G3shGOwdv4gA42Mr/Lt9IIWJBJ
Y3DBPMSv7OqBwZgQdFLKmK6AL4exJmPfZbnhkEt6SE2OfpRaCbmywQjyxrWyJATR
kuSGEnIZfovQNDYJ9dO/N+cGKNuEKuNbCceQ8eOzGKMxDAG2BsZZ/FkT2zQ+6WIh
22vfAmBFouER/rwBOq2IAWLT+07089tGDpMecsxHk4P4SKCI7gK2V9/jf/MR0zwk
hLAGbFs2faRCwd56h6BzJlJ53Rv9JEVTz/LAQUIMZHwT2LuTLN4P49x8W/4jBCcr
FKGhtX5QL7lbht3/ixBeJ9yKDcPxmT5bv9QLwHKxpYNjKMJPGSitD1NA5FgXek+h
v06b+HrtIWO2h5yk+CrQ4ZuUrAs6dw5dcG2L8spHxN+jFHIBRmlswNmMMsI35B4z
mES5qOvK2JBHNq0dIGCPCMWkEk5WIgR3n5nZvyFyjw0Tu3RfOIZbTu0a7ZwBQB84
eMKtgRGXO3A/iOzlf7SFmMaFBdHIuAkKXjXwhlv92wX/+yp4GWyt4wUgS45WDsFu
a82+JPQy0HZ9aNnIxJX5R/Tyq8MOnkyUYOMvGKOzDevd1q3BPsUvW0xHLQkm5+wF
Dc2v7TxiO88pFN4RnwPZKOkSQ7A/Gk82yHUQdy64Z9xzHgGNHxlLgMNccPWK/hhN
T5WMnSBjh7Jbr3VJWR+UZNRAZyS4ZQYZfyImZp4YHhsY4xjONjLTMB8BqLeECd7P
jamgEsM/8PkZAtLPTpp2eYdIX94rrNBNtamyDByAlNMzyn7EcyMTKubl5cpw7QcZ
z0/YKE85osVLV7HUv+BPOgEOZUnulTtwJRdLRiituoX89aTq3BkH1FKzxUjTc7x3
LV+3NILyLGxdE/FTDlk7gNBMFuCQySw54gz1AYjRJLk85NUiG/S5PTfQcWBSRvbo
jRDc7u3GVdZLE2fP2dFdzA==
`protect END_PROTECTED
