`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c1fM6ClO+b85ZeDa/NwC4BhURThSDKsQA1GY58MLoxYPflbfEz2E6kGPz4X4KTxp
YdZZmpfk2+b33p2hkB3momcl1q6rFo5GXx1t9UfaiWBNW3Qr83UVx31CJZx1ywJE
m4x7T9VcX1x4l+p3VqLs6UsFmsnuYISkpljdKECJTMqLGjl28oL8k9FktB1/p2u9
`protect END_PROTECTED
