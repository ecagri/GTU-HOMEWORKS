`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
euz1ieuZ8IzvC9F0bKM9gXTcrpgZj7RGvXZU8HKlOcHSOhGQRrFjrjEHHcAoTZRj
79lqivWh/4qE4jx8rBhvNhd/ZF6mQ1XTJVMUh+JCzQGOH5CaKwEL5cO1aHJs8uaN
yOcHg0mlejD1VXmKR7dA3Wh/UL9C8+JZNvUUhRYmUqSSLNSZoyBsc10KdOsyPoko
4zEP1e78YHztoSyOzc3LjlM5arAGP0giaS8hm4Sxy3Rj4PKnHen9ZPDv93vS1Qiq
gIangpWzUzghiau2EmwXq6QocaGyHmLwAqG+mB/S9nlygnH6j1uU8z0Yt4kPQ/vO
jX9VeuiGqyGLMCWgoN/vMhyiaOcDtxu+i6k7JiAwwAFjnml4+k+e4/RIjr/V0Xl6
+ytar+C9vxPe20PhWO46YyOekAUTbm9xfzouUVU8eYQXt3Roi1rOdmnRmnVdhtke
mWpSyidG73iKN7/miMbUmCfcFIzbSt/YGWmsSB2vYRu+5uAWD7NQ7JsGdbu2cWwo
/BiMUydgD8sVSnN/wwBmtMzz8QZ6p091BdWbmlw0yjKTt5IkarwaclxyC6FlbNFp
BA7l+gOnI06f4qwOzqWo8ysp3ErgDNqXB5EPYD8eYYpX9KTqKKPa1OuA9AW5Y9Z8
MkKUsB3DOIaUOHESIOK6THgfJNubYYioArv7DPpq0x9TGvH62hIlkHdsH3UCKjdv
KwYxFAULQtVT15Yqo0TC8tx6Oa26agIC8tXP2k1k2FraOO7Zc2ovfzMC9N+GVgmo
LGW4MsxSZmf0meepJ2ovUA==
`protect END_PROTECTED
