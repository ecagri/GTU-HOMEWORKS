`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vEsYHJUNz7Sgws5tmglMtJvboGNao/zfZEFo/aWEv/IiOpWheqrN/Zzl0q8Ewpzh
EGGXxErQPC4Z30n+FHZblRZjxcmFyQVgUIqcUsIS6dE3vlV/4E3YGc5/MKAr/SD0
O9LTxYhyH7mrbR5n1WYgigBws1Ra5uZfcSOndaQ8XY3fTUPTcokMhUBx0DCp0irg
mFQEBkTLYwHQRdBvcX/tCnUqc6lbcuC0FK1JWdWzpAKw5Z/RL8KiwNL+/l0K9QA0
kxUegZP0ahvo7Lsywck7QU5ghkN7mlqcHkU5V+pxKJGXEWt/1A1ytnXXyFr/nKxa
efbrT8Ra8R1UnT76iapFNSVfKD/jhYmoZGscRxWJ3WxRUpgmRF+LVbo61u0zJL77
hncDLHWOE71WLrxpo6S5GpLXmgXHig3RdttFCQxGlrASZrmtQaOBfPs/rUhmQPAa
MfdJGYQ53B4+KciI4ZSGTqGwwJZnewBh7VeUFO4ExpTMfypwXgJkmwibAj2a26VX
AzXgvfZLeFCK9DlyBCQfWoqdnmRUrFMGyKsKK+6wFc++XA0/vImEEjrEYNpgl1cV
vI8p8P1kFsbdWoI879sJOFeTAMkFe7esMMOyIs+NbTakDVTFfsEuPJRNfCmW+UEX
/BYJWyNvaaa9VAn5ymlxHcq72XMK+MIVAOryFwsuVI3i7gPPEx33eZSrdS6WzBBr
FKFGM+j8ktZbTKyFuWiKSBCpMJTYZ9rLNknPAer1odMw8p81NSk5tq5AiB8nBkCS
kp65YoW9FoWUrQx/BkQiyFXtut3nWQSjZD2ZPA5XfZHB6RDnWqUJFJqpNKO7hyaS
r9UsjZXK3SbR59h+471HeEleOaI7eDZbO4lYo0qy6DBX8fOp8IytF+4nRBB9BqJy
rHRpF5jHyY0UtNImfkRm9pz9xwyMLViGkNsnwnGnv9N7QSCZrrqtRqPD4BSiWFwV
I+yakc5/l6b0Rw8D42i4sImsA4bjthGdkFTghLHA6ahEXkD5umrm2mG9S30ciexE
WdxmtPrJ6617ot2yESXAsFW4AeqGthtCexOmY7JJ+hAdU7qhOPmjgVvLvf+KC/EH
erb/M48izKu37MUDrlJiQ5An6nDjjaZu7Fippphy5x0OH5h57AY478jMcKeo9qi0
CjhwjyWK6Aa06/Fw8Hqb3lDn6jQ6hhs2/DW7cs+OHPxouvE5Vb4ixpSVkVEAZZZ/
eMnH6spYfArJIWYOxdYjHHBUz2czql1ClZvbuRTyBCI=
`protect END_PROTECTED
