`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rE19D5mOH1HonyjI2ViaNzrgBJSONXEjIF9DFzWjUJdKC+x4kIjnc9lmHSmIjjkD
dwPOWKxUZSMUjFqdi8k39UvnwW8uRvWl9nynxpSxyusF5Rm68XgqG+idrJyJR06L
3Qpi+taWBYDp7TXHbd/yd/QZxTwTbERlv9p3D8exlyHwflVFaUZoOnE0Ef68ugGH
afa8npMuWUPbFwZxyQRfISTr5tPfmfCYDdjzeO+qyk2wTNwfea+zfG/xhyGxIPpa
NIylnuBewykJXg2TDsg+ApYCQGsI/As12/mw9qkDwcqUpWJJRGfeP+DYpUD16I5Y
vX0XEEgsKaHNMYV2NLf9P9jhmoBy6iB8OoSIaipi81tcOxNkUXimuXlPeVxICaf7
WmAZXSCJuEgKL7an7fdhQxgB7S/Fi+hMJYZ+2pJRXo+H9/Gkwv+Wf2CciO/aqC3y
dXa1T7IbEHIv/JWKDF78b3A0QbS/XuykG51SSskhT+/sNuEppa4/Ch1BgXkjPVf3
pX3AMW9dxFMxOpIF8+6xxrA4W6F669D0TPUL3PgY9muRn2cHyHtKNUgifvnO6FkK
ISykhRVuscSLRO9ZDK3QStffTRvP4Py3xlAqKhKd57zEtHJlPwNiiMqKUXehxHoD
3EmcP12q85fJYh1Ae64RAjAUL+N6dlqSKWIbDkqRpvZOxc+A2n0UbQXVUZAjzT29
g7GoKlQfI4zeuqIE4j4rsTdpmkmyTNRCEorkUWbgqusDV73g8RWPkvHUw99Ea0P6
kjdbgf+2lfJ5XFbYbh+vleGr4TPTdeY5yF5YMQjhiUoJMLy99ztd4kjLtLmQu14l
GLOi7aMoqpRf9PeTuAdV47Q6rxek+lKhLU4TUbqkB54RAOu6u9sHN8F3f/OmYULw
bUT0hUXQsFC0vzetasfnA6exV9sR+xbG0HbmOYvRAKL8UVkXbBoyRcNALbR7AbF7
qZ1FwfXNRcQvDCSVszMp8ZDwTPCAzJDS/XIJPV6lTfqCXKD/lcItyBN6IvrZenL5
f56tZxgHWGdGncIRaxWZAXkqN78sI75Vwp3ADarlnLOErvpF5DTo7ELTHUGcr9LC
MKJuvSmtYzAcI0eif5YQnHUy9/5Om82mShPytwdK+G4Rr4K9W0Ll/O9H5r07D44l
WEMu463AGMu8OubdZjFaD/+OR9t283+VR27ju6iyowTf06wS52bHqUAAK2GyXi1f
BWThQJLTGxKX5r3Cukivx8Th+l0nGIBF7PE6B3alG+tw7b407zFCBomRVGYLbL0b
rypVUomAXf/VeFjmnaN0H13Yq3NtQoG0xNU40GLyf6R9q/ySH8urZADdowRRNPIB
gbAW77CeFKSeDINJpxyARiL1EMr4LmTaqhLUrXascToLJ+Mjmt3bIos24ZRmI655
ZSHhrremiBoUdvAGCIZCBxguDEJrouYQvmybt1LHsMRVSagbUDVGiw9nTsk6OEeW
2CBM8qk1w+sQoBe4HZQxsU6J+4CTLztcGaH6TBLlI2h7LRKHrfKWAYSEq4JXsliX
dwI9UGzHNVJruDkeMRVW5ln6FSb6J75kFbUP5zPftlJfi4i5CmncEX7lsTPqhvvm
TLHlB++AZZZe9UGwE/prliaAA6jM5yJqDUv50ryc5DV1HPYBfxbhN+w8bfY5yk5c
lA5xkpC6cl03hu84Yjkit/CImrvW5mCyPQcK4cmhlz0nHdqegp8F+hVDKtVxK7Vj
YqnsSwB7YTKIZ2VC+y1TEB2zrfeiNs/Vua4+zYgJ3szITLaXrCKGzTKyvCpSKtLV
XukOd1CTLlZYarEQFsVcaRFfR1jaRMoXAPLqZVP3rrIemyu9GJKuivlFpPceS57n
jrBN2fgpQE8CnJv4sdvSd9eAFPZ/RxmafkzeZmV9JBxTgAuHEsTLGDuM3enfMiHQ
oAdZ2z+D/8uv5G2NKnMKp74p27YhSwgp2pjIp6J5eIUutlVRJONKC/BEOzZyZ3L4
sC0Lb+pLL1hxj86rMVEsHXDoZ7aw/8JehZjeGEuKDako9VI0zqyf6u394/t2UprT
1wuNgZrysIsXlhVGmTPETWZUoHiHrAKE2G6JvqCaFnAHBEMvM4oBp/ZQIAibhUeY
mET1k9ZNZ1TOkYSKOIMvHKX73ZKYYmc9d1cPbxCWX9kUltlNOXenhOFAVho7Qp3d
/ydA8LRMtqL4lZeo4JAk062vkiM7uhvFNc8AOUqy7k9pmFFpF/40IAIiOhowY1HF
mEnsSqz7aLvwzAcdkWyppKHKOGKxtESnA3AddLet9dcmrbe8ChJciLQ7d7mY1I6c
8PIEvFtv3C605YlaiXUneKeYTOJUNwzjai6s5Cz1hupda5wnUnsL5QY+ixbIzH3P
yfZSIr/gHGKULC+RP0oue+++k9pLkG3ys9Lh5Hv5MxDladBRMSmDO3DlBCLYFWdt
O8tm9U62weUhFPcF8wYosggm49cjRgHii2NxTj+IOvaHAyttLcuYmlEi3pztDoMa
iZFi4lT1Rntw5eoe3tFiagouAs+0rL+WYyrePWAGypSij5SX/uHu6rCnZmKMIOz+
Dx9ajj+DaQbiqHPehqvf9AtDD6fBwr1+iUlGip52LUQMOnM++uHDn/ys3TUrhAXQ
6XdZ9LbJcnqGX/INOf07Aaes28PMKOFYryVYkX5Nm0bLpvhGMYCuB1OukH+wAqNl
4YidKVodLrZAYMsP9ugu4fNgt3GiQH48jrk+k1LnhKTyj2yXBJmoL0lLRVx4nrgh
8xNobf2KC6Wruw+rbRJaTGsa1gyBD+FmN6Q2Ph0J/xD1nsbp2sYuDEmBkKIBFyf0
45kdmL8ViR+VSAHLHFk6F+Bfa7QeKVPbIe093QQBS0L5B5G3ngGvpXM3xiUcxhrp
6jh7stlTB2e0pypw0VyAYU6dHuJdwCIniGNTVD/eIW1cTyZbcBf+E7jH0qxzKstg
42/e2pqDikoRCkhC30aDqJkIJd/eqAZz4/dwszBHMGw1MmSNOo4WCOS3cBYexXK0
xyXT+TVDYoKSrr8ItA+mAhKNf4xMfKt1VENMrc23tcAzRCe/9+G8h2bxlLdoYTBu
D73A4C23ae+WPCZ/6xaTCWEtl7QIIvKvqA5wyLCSc/FMwtSlrXll3nBH8WUrjFyr
lvvFHKUn4QMRnHLgU/KM5Y09AteSPTv03Zs2Obt1UJXMzjbiAypp2/2nZpa3kRdU
m9gHQZLfMWlshMp7DYKqlVKHC6+XAryv9mW/rcxFR5mliQt43MGoYQeSJY9mNxrh
Ho0DR4GsmkZ0NaGLzqLOMy5rrrKLac0CeUlV43lRIKGNBifYym95OLaK6hbtQUXr
LkQPLVnPmlTfKF8wdBatNeq8JXH0GeSiTvFsdb047vX22WoN2w6kjXjLSdCi+UQ8
XsVovw4GxfUvBu48BKrjLL2y8sSgM8E72mTz5vZ2mtxT+AqazBTBT362o1hsoQxB
MR9I+9p6zXUJIRqKz3rLCehIUtZprcdqPt+HoIrqK9TxxW2Ubi3SeA3D+VI6+BDH
dM3cRPiKxvm6weU9F1vDZIP9QIefrMkjweq3AJTijJ2UQ7RkI9Okc4hnKfSB6ncD
AVJARcAfPzP6Vz8IM0a24omDyLpFRoBjY9qcrS3YvDvAi/T8XAklh7ORWkQl1rbB
Vdxxs2wC6rsFgyDkQ/2siDkoGO7xSzR679XnQ/PRPVxs9GTQytBo2TZpTUvhttbg
60O7ZHLz9v3tDyBFdNE5n6R2ZOouBcqUAQf5AombxWf85QRgyWMwCYUO9/7eZVJt
EepH2NWPeIHc0SJUnpWLz3zv++y1RB8VQq6Lc1tcUIuSowhb4kvujoVWy0E+GXeo
HYtnKN/dG8gCcguF+epjxPSrcLV4ipqNY+WIaTv6YRyKnLWWnpmVleYXsLA46q4q
d6yyHtvf9ucPcRelBLDHmW+dnX44rqGxsa2/r30ezEhItw0zKIJ2F+WsWHOnWona
sMxpUYtGFnXZg+1Xnjfo88d3U4N1zPA8kKbZ3KnCtw6KZBO9/xiuaqlR8J24jZlz
aQpB1NNQ0FKOD/5//dnaYW5KHWzVm7LbdidS5huAsT+DsuutJAmRnoJr+IUTDPRd
bd+IwVROQmdFAcxvrsOqC8d/HwQGvyp9RqRH5ntI9t0vZCFccQIuoFN205rYUiUy
rGNsQq6GNq7C7/USbxawmwsAYWfuyxuIpeE9NfooWRFnKbw2snPPvF177Cj1bA/0
TUJsM3jRWcBieNSzRJ+6gGiXY8tLTtch2to1dBXKIeLd4g2qJG9VQG0W3CXoA/h/
pBnYB1Zr2QyrTfee+kOBUaNvR6iqVdcTT5eAq3zCmyu6v4LXwgu+uiGHLrqv4V2N
DrMje22OZFfS/n7PZeaCBenZiROrpOHelO4+5lPHv/lZ6ygHJIy8oS70h0CElxeH
ZggBZv2RG50O+Y2OozxKOV1uZVwAWp3Ycsc6Zp1FbIGYGGe1a0cG5XR9/Gc2fn0R
tTCMvQ/lWLiVh/n7dszbCr6yrVa3u1KpDVLIRNmCHKX/DqvcodcPdgzMdJ+7v+tl
/RZjCDkSPw6WDZ9C0lqv6r/B7eou+gHvZentIplr8HiCtYNM4F1t0Got7qYqpZqG
S0Md7riQ6M+prfQgIHUkBusIloZbLAJyu3A3MlR31LyJ49mPNreoRY4rHiJZGWu2
LKqaVxRbEKECrKgBHBOAPxeG78MwggysikOF33bXSUAXmhQ6JNd6qXDlxSQ7S12H
yujnbggIOGtv1IUu/MyOQ+wdkrSAeHoK80Hj9OHCLiSi/bszOWlwqz9CF2Vcq3iv
SwOwLWjOFnUv4LilxircAp+5CrafqR/H3EhGEFiaAXrtVyiUPXlCJOSye+Ndzzxc
Y7msUp7izv1l6IQS6RE+hAdN77ENLQb/+HiurwH2ede2GJgpQ6KKEeQsgSRm9RpP
+PrPxxWsnpd3M5akeS1k0HkFe4vXeTQDZM1AebgwMeD/pKFr8YRXMI4Cf12fP/QO
vuTQIFWKrFDv+xEA08fLK0qpYL1+GzTDkXac8rZ2eKa/bhrh0OYyGIrQcnQP3SrW
Sx/mmHP4ruxkFC+CE9I5LF+hIMtDpO1BOAvm+y3T912Tmm347m/ISrpyL1cGxIC8
32X7CKo6nf5JQxXA8ZTIemCXNaZdJYQJEbwCVcreuTYay1aAbymFyH6ZOwVkxgoo
L2CLOwhNRVOOkwTHr/ykq9YWgMJu5+PhUZOHokbA1bTfEtqHRYHK7VowPDIgdSSR
w1R50ps+KkoGc/WBMsABvyzvBcopKi0AXkwDEL+nQQmaweE7CDyNYJ48waVp1DT2
Y5dsIBJPCTBV1KLZMtzC5M1w7XF1YogA//c1CxMhj5CnARiI8i/f1xxhcCi2FGcQ
3xKcVgaz38PyHZZFexstMImJYFixHhZecbsJNZRs9/ySAnYWwWM3x2fFnTQAbVdO
P5hCtsLTTIVTsDJyN4uwhCdWiLjsVDV9Vt8pRStFNnaUhsDEhMKs0FVQWCq2c5QT
2myLNm3Nr3Nj4bu4insdl7N6jL4wy0OAmxdfFJirE3aPXHVC63DfMoPKPh2d2MHH
/+tn1ZZarXmqAZLPP7UwHj/aNbeHbqsTOwzLCk14xQ/BklJ5BAw71wIW+e9wZyhz
ZNnHtWs/fPrRlj58vg0z0+y5CGfiZGMzh9F64Z8AYBON+SWwuTuYO14oqy2Ss0qT
SIbheUUMSPa3fzixXpiQ6/LavmiD58hHKrVanqfuxyWOKGJ+ZZOJpgawisNZ+oLQ
YpPHg31RliDcpgOJVI+84fqJ/6e/KbAoaCwYTO8zRUdQG6wuygGRHFvB0XHXjep6
RtxmFrFZ1/OQYflGRqEVhf4v2rJZoGrj6JBwabWf/PDnhbO5nrfgLOV5/kmP36Ik
+8/G/SJV40OfA8W3zUR8dgQXlbj1kqw/ya7KlG3DItNrILcMuhFf/FqtG8kXG4mC
oJQFbmJhd+jfaUAEwARWcxxrfP5IjQiA/eQhif5O9Xi8W/X4sL29pVqhkraH2zdM
p9yPAhSvbfrlajLg8z2D1+yamIANYneHn4JvX7IPmoe/sYillymNvgqQiHroXUUb
0q2BMrfMkzhwOsPsIRvdcZTQB5iFZZdliUSPPd1XAUVjk76FfOsjVPFNABmoksJF
+UX0uGAy+rhXPA+zYu/KJi7nMSL9WxmTbPejbYyMtmYzJGJtR8VXezTo1OaH8jRt
eh8M5ww13/Bf2TtMZxl6bMLlHpx46COByA2hx7EPbni7fP8yJAiTRvZK01AMLJlU
k+RBxfOUvqhdQWEWLiuXaltoLcq9QxtTox39WURsG+qIh9rrPTfNsE7KPzLI+cgP
VANfUOzSNoCxEIhtqAWbQDuwIpBFTWBrQF1suRBetgg2hqzR6ZFQ4HeRV0glBWMS
y14lDCVohBxJicJFLB+KupUM8M3ASEUpViZaWQvpdWNrui2HtC6hDPgZpMLCkhXT
Sp3udQFcqqrUClvaVhyHeslpD870j8dseVoTtxG0t2v6kZGeN37EW+zZrv4PrCo1
wlSwwqLniva7fx2tVxtyqtLMzzkG+ae/Tm4PTCWMyboaTRQDnVyMImmZLrkTjigX
FU0IAmLe7d8BruCSV/wT0ZPy65ion82TAvYv2K+Rs5B7k1Mt/0/tdrM1DOdO/Ygt
UYCVoEfmoD4wmOQM53Kq8Io9NLNxI4Nf4iAnjz4H/5gxn/frmXZlwjcIqHzcjyJW
laGi8F9sr2NcSnL2BrmOppmgoXF9SQ53IukRgZm2D9R3YtQFA8NzDQoigcfeqQEt
Brd4n+P4Y0yfHNX+/9AKV9XXcTu9GM0IZ3vtaW4eZx0jvhao2wJlNbkvlTxQZ1Qh
N4V2kWEMXhWjyc7xsydIXnxXtAK6JyY/20BgGr6xLzcxMxB+v28upFYyTrCy6/FW
AQVSQQbG9JTo4/v1JeBzdjffMWgjFjXyRAmSXMQ29CxSiQgiAAaksNem9LMJWqsw
oIkwl80SWTasI2eNJtozNgj44v6e2vC5cdzg3dIV5Hsjl6PPratEXByVQVCZr0Zs
fSj3YjgGaXgGn553KEXFQLicXSoUZa6cmv7UKLAa4asgnXjZ6SALWzBTYRnQWye/
Tg8cP676JUR0BXqmmrVMTw42qd7z110izp0J2yt1+hxx/rVlKNOoYsnG5WYiNwrU
f6XIhv6q7nn1YaqQAEBO5hyFTs+KwETUWjfscxPmvmykaJahLrtuMDkezBpqwsvo
2cq1JPm+CMO+YUalkawsZ9/bNqtzmo5hpExkxqbjtwzyhDSQhGRTqVbRzNcB3aY9
MNIXQ5KsTx0JnAYer2nDZGRWgvqfvqmXrE535F36hWU5zj2pMO0+qZrvevFLHhJ+
kbc0XwcV7UpPwIi1wZXJEf2T8ruCG263W5RzB4/3hhJgjJpZ4Ux+RnzSXVU/436P
LzopMN0jdy8Gd1fsyHwsZRFTQIGk+5qAT8dHTBNrEa/9tiTwx0UcHuzzzqgb662X
ZoqHzZPaJjtjsqonQueXpmmZ3ZesVkx+llIf7m0mKFaWbnxoH3Va8TkQ7rKaKlhg
CibdUhTP5hKciA1Cr9J7eKj4m5U6OYlo/I1DQG8vCt2vSChrlnsxgfAOkgPCAf33
Qd/EnnmRURFi5nej51BOd+DEEcxhwDw21wwgrm5icnR5qgzDxTYXrkHi5nNsakeu
TwPLfHHGxVbbHEmPcIp0v7OTmbKBuHiyNHh4CQ7RJEobJtgB0fDNVB8F7Z7T8RKq
nRNiLCvt2Wcl0ujGJ/+z1uIXhI4S/CiS0GrWR94IfmmdQxC4tF8BYxTrO2BIpEow
GYn4Z63fs84fgIBj++X/Jp8daEHGThPIU0jHJVIVuMJ6W+fO5RHOIxbVf6ndSWeD
bud9ShyfPWH8qWZpgduXjZWCuillUmRD9Er2eYAJ/GsnXXL5OE71S0cOCncpZh3i
udb39UmzLtWGBq975bLO1Z+wMKFw+hcvQg5nFLQ8bAYNbcK0mED9nLQCSIO8tNzq
aMOrqOBwVrONu7VCoks7DUuMI0j7H+RvNjWX8cOfH0B5/rK01tqsVWIo6UoZTzz/
Eg6K6BUJm6/VWZMH77yecDByKl5/+zKWU0IHI3mxnywMl7lW6tUJ/eCh+gxuChQX
t22Tw3WUphjjecHTaWVDkTVlxWsP7de26xFP00AbN9+ZhTRZEaFFhQ0eTjm8D/ux
A5+4elB5j6ZB3qZHhWyl+8D6kmUpP0kfWeFTkAvXfB86wcDfgfz+ybHI1vuGH2HR
czjanpDd326KQS8Y3J+UPquMdtV4N5sY3cvMVgFLlcQvdSc8bnJwTxs4a6S5RLZJ
1Al9PP+QHarNq4hMQ3C9l9yLv9VF8KuBxOFPrnEzdQLV/RKmz/SU+CX+OaySFSj3
0SQ2OZxkW3W0YPY/ky/B68FwAwoNK90BfDZjLg0NQK/Wlp9yWzn/hpQcIM1ypfpa
YZB2Y0QY8L1TxQyh33NUZef0DqWMVUkN99oMGLH0z2qHDTX65GIEnhRBpq16Wfp1
KTVomQUtZ2Fzm5X/gJSU6oLXb2yzSZCCjBtjQxrMvxk=
`protect END_PROTECTED
