`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DM3yM46iw0tuHxchY5+2BUE5NeN155ReunAotwqKuerEC27q6u48RQD0pUPGVjCl
iBJnG+d/ePh43RC40asO+84n83akpwZSnB3QNEcC8j1dyAplMBNoteNZ0mFrUjTG
aouEPCTW6TnBDi5Mq1iH7gEnwNmAlxeQxRItHqxZ1kLgBgwAVUVcqa6gphYos66t
EUU++oalBw6MR+pnDgnws+tJJ0NmVYv2cjAIiWnDnW0Hz0he+jo7W7tNY2wZhyOe
5pl+QLE62nFwFz3ZsVmuj9xGXSJtFk/t3NMytZoXwhnvIFMWvq9ydf/ghlQSY/jv
bzuMhLvwnHAeCCjwwDjhdSEk5r1ZTYfDbClF2iXqqeOAVE7VPeqitqbaFJyjv1VN
XrQfSMJjwa1YqmBaeqd7w1jmGkc1mb9ji1FIs909T3kBHXVVO/VdzuOYjKx7Ku9F
cU6MPWKQJjrkmBHYjQfFLze5XRKUW5rxi1QW6wjcNwzyVZZh2BfNcp3nrGHXLjD8
SmCsogfeZmSbslIUmzAi8XqAXrdVXSsdon8tigSGLPd9zGC2WeQDqR5mJNC2SLI7
KiFY9I9WuWD6MAaJlVzxML0FB3VbfhpmfsBrLOeEzZhc2QcTi/cTtexcwr/dlWfJ
aH5c90RlSPTOnvbCew+lomu2Q4NtWcByAJ3vGcBoImfOtANE3ckzxmMcuOR5V4Iz
NVWD1JMBzvNujY9V+eSN7vRaBCtaa3ViW86kBJSoZdL3YkhtXILds0ShDICHYm39
f+QIQWFW5urNtqLcTDc7jLtxYs2fm9broXdlSXg7U0XCTU1lqZr+rX0GnNFQnftY
k8+ERf/k4c7ENdR613TS+g93gDwrOQTPKHrBlbQR214ovUe5DzEosi5TbAmMv/wL
7AK9BdosTBHTpeW0dZsTZ/CQZLqt54JOHFxtkEtCQ4iwMOrE2dOirZ6ce8s26os3
Kh1fisZv1kEv+tnqocqzYCk5RHkQU+qfuYGgxnnOUuZfABT0WS6lOOBx82n4vv9V
U1UcEDEeCAKT5sL4YFRsEL6Y0E4JI7yPeifzAo8t4QbIeOEcKHkXip3pCj8fzHtw
P2qs4CfgSIxM84Zq5AquvCb59QsnvID4Nq6t4dvbUbkYaKEzt2BT4CZqKciG9syC
cWhgVw9eppsfQxQvDPeWLUJe6bu84pIQHIN5nh1yOfTX50d7cvAErL1dXMrZxMv0
T4Ly/hq4gH5RGQKYhenkzE/OWX7N5eMnnYR3JWYKRjOUjrYgj06mhugd1+iQgA7P
RNDI1ZqfFLv3KJV3bp2j2k9OyZoaeJ5gsvyQUGprjQpis+Kv1IMdcwkfrXdU7Nn5
lBFZYKHANzYhzFO4fpbkR1TzM/MXrTtgnKbqLJrOIzlsCnhd1/AmYJkib8mWgnFj
kRrepmk0xMzDAG5y9i/afYQUrb6nPasHTYJfXEcoWzHEgBbwtIG5z54kTmR9gOcm
KqwxmTel1Ib9JP6dEee3Jq9r2T1E2+qkySzhq+SYhdSbKBm8SPn8wsSq9MjsyJm8
CbGITxzRBw/ty+kxAFgv45N9lcVVO5Jrkbyu9HIxX5FTGBUsc6L5WZpRU7vziyTH
fcYwKsql5n3cFBzidQcBvT+U6YeaoI+XoYWCF5v0Ml32a1pokHNoCikB/+KsvQiW
W6srvP7FHhwJgy42EenV9rNGNqcFAiz1jXPyRhDb/tAW3lBOCSX2citWFMS9ffm4
c1LmJ+MVIhY2VhKznws9uZJlfTswhWCJ1N2ITkk3olcXX/4HJMay8vmrI/1dIOdP
VgztweT6z5JKuo4WTMMo5Ta/WjR0Ed0HQohU7z+efudiw160WFEPL4DQj5CloHLI
3DeGnK1S9ZJSzlTDKAwWnKJmSSXvURcIjsFMwNyXi3FIrkaCka177RnCK+PYWcWg
2SFS8CVfVmHxMZ4hAca6ME4Ho8fxjeKo6xdB8k5vUJe3VjHsjxgwmRavn/X1Qyus
8ZRQERQs7aCSflN6XlpxGG06ExhXeTBTX1c5KxV9cGZMtFjWZJ7pxTwRA/LPds+f
0GIrFzl7LOCiryIdbkaDBIOvoAjgQfqRkq5Ir0w8EsHn9nEPYhN1jGAVxRRh226P
VvcTwRVxJDAzvqhGifa+uLJU1xT8syGTiNY/wGoCb1LYRNFxP0J9h9MzB0aj2kOy
rTUnAt3UXMy3sXsG4zHDIA0ClvytyflJzx4YpWwkvGsVNs6kSQApJ4Aajt2bfRbW
Gs3tYVAk3B6CqSFurG5jCwYBRy398lSEtR/aOR1aUl7/KyN09AlJ0G+Yy8G2qzIt
LFPRgNtW0wTqSBGB0v0IPTzp7RoXLD6DcVKeAXXJphJiiRUl88aSCAcJL4OfzSSV
qc/AjKmesSsDeYRZSh3XoKWNACeXS6wO4WurHlpBcPHWRMltLPHIb1/YSUifWw8q
VCWWCJyriP9IClo8XkNRLCDT6YfcEQzLNsv7vJ+CUyV+7rRnVaC7+ObbQHPd8/B/
DZ14Ex2GQfsy+qLmLwHcefDHEOWH3fWi+bwlU33GYoi8RXC1wtPTUd1xeBy7Pm3v
A1vrr9cj3XlRwwza86q+YJKB6mu4uRUcTJt2dRv+4urhWVXqLwnuBsCt8BcSxd7b
KEkpkJLL+Y2b0eUL+cXjKR142iknTQ0udj6Hc6LlgHcdVujmqodcqOqcnbKPBu4p
UVZ9DWeWdk5qHL1kjho/i96ut/TrT5AhNUCz/yjcaFfW3BE9k9UppB6Ja3fzxHF8
aVeRexgeOrfovv/jhlAuSqdZmuhcuIuCSvr/b7kEunlzPhCL7Buee6oghU/H1/7C
uUbXkRnHRiFadBYEWy2b57wg0yOizdjfX8t4bJriu7+iurGqcnTI1EOH8C5UJR3b
7AVw3VPSYNOkIL9KBhd/N9HrYhmPGoaaddSvGwD4TUUhMTp26qoBT34rpamAfHH0
tZeEMyGi3c9ZcwvuSrOxoa7GBv4u6PMT+oHhXPgbMzNmMKBjYDy9hlMdRNothCKz
kCAr8BWdk0J5AZYkHW40aB/2aM/zEgDXqccd2iloFC8aZc2lrJ3S5Mp8uEMb1sKV
/IRtrs2QCPCrtorqww+7EH/RMfFJRcaU9mQFzWm+fyqgJj3RSqgYxhAoLN1KuZh7
Y2ES1Togjf1qYze2hCH4fDe9lOPcWSyP0m8jyGasO2rMxdxoPB71yUXrqEnJ/5yS
DuOM05psm84/5kzo4qo6lJO8HAWII3Z6oJM0WOTW8epx1dD9ocTZV7iMZN+Fsw8N
pqIAFsGHQtsA6Og2Et9sR8hq9iaXBWJ73QUHD08rfP3+7EoVOnpyBFAKloJ6Wdj4
EHzua4hUepwGKgfIV4ENQPaLWWLtnx8T4eBKVc+3PmX/RN1UjJaWj0fMJHm71ikh
LXTdhCiy5gCitwemQ/JdfdHl/G94gAGvE1eixmr1Y6vXPND1SDKawVJvGcFoYWvB
gk3dnjWvJS6+i3y3Z/Rc5+5vh/1vJ1PYciQnZjiff639SbgdxFckGHFHz0OFbSch
WYathvyNcDQ+UgXfVtsGzc5QxYolcDSu6IiNiVPA4kpTKG5jTerJu8U8dgSyeIIN
yzZWKoPinTV6TtIoPlYZekOFE4YG1Db2QbBOmveXAIjLy/Zm2Wbv+NGuh5rkNnqu
fyiYoQIvBFTmuEnocsjxSqQbvqNOi2rNwyYY5/rlv1oPaVppI2CAPPa24WlGwVkw
UgJLLUaDE7NXNWaw2VAHxdZM21pSPWHCMpGGDOVVeIqssdc/XAZaJ1dTm2asdihl
TMYopG3tgTaxF1s14/N8DNBfx/wRAY8ydOXnXHD5LlPHiyEZPgqpStl3bOAOlJ0F
Kj9CYo5VVVYKlstjI27Bi+xO0qzv+s5AdY4/f5t+u6ZLGoens5a6kejcUhVgHNvd
WJt71i3zhFv2fbFslZ+7Eg8deYPuFJV6mXroMp61iBOO3zr2yQY6voz3/WPKY5yC
G+en4BGB9Lfi64RFLoGUGj+61gl65I9wikPeczmaBXvnDR8bmMGP1Pm3IiDBFf5u
fqgBdYTFqHtHH67zD03U1LWcDEEZmc5rFNSBHs55y37jStJkQQV8KrlHyCUOmgy7
WyZuRf6sDXNH9b99NWQerY/iEAN1K/o1kNchmFVL8u3nN00wY9Mh4uwKV4v+C0Jz
EJaY6K65kXr/WdUWYt488hQtawtF+bYzyaKYv6gT/YCFF7kQZK/BUeC3d480Do+u
TzoV0vjiQ1GnmFxmAS1dSEFf8FZUK3MmqlL2pQ5xV4F1hBUZ1u89pybvnOgCOxAx
/i+4pc0JThlxxrQTmrF5t3S/H9otUC236IP/rs0/MIO33It9EkTLwlE7BWf72/3j
65KibLj4QF3dF//++g4RhDzhfOzn/2WH3sqwtTt4nM7xxRNX0inSjHphlXfYHqpF
55OFz1m4fdN0MjqpKubOjcvv337bosY2D+x4uDNoFWEQPcew0q5a1FCewkovB+e+
rDwG8A4TgC2fwUotpHHoSv3r7UqjlPlS5AQ8zEXorAznqUcfYtpIA8P91EfPqX0y
E7IKqOltwAaAPKBRUBNZUrmMmSTgpvwU8glEHS10Gwor4/NZkHfI8TdmvyD2ty3X
iawgDPpAu0TzS8pHe6uf7gjYMyn6DbY53qMkxtHF5xSf8nV/sL09zEy3fucCWg0x
EwXkBLjfO1XCQkwSSbWIMiHdLEgXpPZddaRDQ8TBhUwOUSHvq/VpscDZ2DLnpG9Q
D3ikHbEU6DXhlTEiTIQXNtnvmKZmXbO9Ln/NUuWI4ta9/bsS7VIHR7/+6/2I/Xky
tEd//q4mvcMagJ1s7c3qMGsPJMpGVALsQi6eRUj6cT1iN4+jt00z6As/DDhsFkb2
1thBLj+ts81rIVNMWmGDDiNoXZCbON6oS7qmLLbUUzrbKiJpUiPgxWpFnuEDz2Ty
A5G+NKE/eXlIyN53gTIruS7bY8RNLyp21s3FdIf0sAsruM3fyv3AKi5vTpkO4Hlf
+iRjJVTIM0DPnomO9oIT9pnHv1RlAi0ucR2mrG/DrN1rvOIC/bSbnxbqwj4AyRwR
5oIcNm2lswohvR12fTv7yM2wbUCy2YnhL+/WSRcSgvrC6UgHmrru2EdzYIFk4wpW
0HKo3+u7Tlclf3UnDM9aZD6+VxoL3FOF8UOCeijMt1+kj0imDry6LsKKwfjEyffd
Zaz0AndNpJisKMTEirgFIY/ewDYEUUSy6lGPhG0yCqxEcMgNmxlKWy2mBTR4EO9k
rBCbL39AYLnYzTyQZxIoWB0oOPTLfCV9hwoR4LW9KXYXuIHxLTaAV97oIqMvLoTw
ivH/4Bc9zT9Mp0T+iAxHQ178du6jaiwO7PYvQ0MqxP8xg2mcltvWwTRqGvKnXuYI
/+ITs/3my/9sN3sBL8MZE3bVaFMLyEesjgBtElUjnYzI7TeViHgK6nGwGHTcyo1w
Ll8CJkkxKzPH4eti07B4pXcz7OfOUGUoVJ7luCqnf6hypwcfb+NBfgYYFiEkSU9v
urd0UP65NuMqhK9YUzZAzLBdZEe/SlH1dASCFj0uYa48oOvN3Y8qoGxhsJXhhBfM
W1CnBuZ6DmI2NwGLBRuWuqv5gLiBeDS+0zwxH4t9Rl9YuqockZJ8Np1BXgzadW3+
09UCD00J3Y1d/IrdDpmF76Z7jLmeOmZtK+gYtz6iDTw4hrtvLjCjG0d+S4MsHoBl
HCLJPlECVP+lX/owykcwJ4JBCY6Z45JRJXr2PbsI8g9HDbecKGIh+447A9uQsywF
m/e1jjL79QHGCxpTBZOCyMN4KZx0JRvu8d9etYvCdOPxYP9q7b8KiJSv3zH+wa51
ITw+V6aUMMPGKTnZWfZOzjq4w969eErE7XOGusXFuXRgO6k/1Dv+TdtGilrUoZff
lNm3sj8jyCUnC3YDyzGBaWvZtHHceuL0IaLO72uFQlSD7ScQEUfdVktuuWJu1+SP
dNjDyu7W4EvRqYdtzIx3Ac6ixzzVdeqQSxNm4dxoTm92G8DF8Zdo3kdPYKV1zzzH
QBosgKL6KEe+M/yRuqJiVJD+X2L5jFwebjKj24XUGF0H7T+ngiu/XCAaBRRETDqp
cSyamTLDgMO6nOEYLfvxnBkMWW1Ukz9VwnWxCN6TfBPy3kUS6iYT98VUn0LQZkKA
kvXnPjf8A94Fy/zqJGu7MjRVcinDbfDgntV93BlX1NizaTJsAqvVEuqXAQCUA3M6
SwZfo7gd8cFZfPbJLDZO8rx2H0RKUPsKKN0Wc+JT4iVOVzyv5fJAd16n4i31+MCt
U3a1Na5gyfkx8WUg7SshqzkDRnSyKrDroJWUU155TRwtZox/BzbLzFBXb7AYqftQ
vKUfA6WHNBAn3nDGU9z/HGgeBNzC8L4jC6UZhFPY45RmN/RSnKoBbZTMKpJRxLtP
IRD0BafHbZf7Ix0KZKtAaBC3eIihKW0UawOFBz3DvrXkywo5df6r6/DTq8U/45JW
mVmGLIkZaaaLKMo3JHQCwy5fecoo8AUil08XXuS63aQYLNmx01ewBWNQRpdO7fcd
+F3UgkARfxvSzi9tiPOdXRvmDsZPPI2o8yVvLJBvXEkQn8jL/8yZDJQ0SvnaeAWh
nTVDYM3PzasAFPHC2KTYJxDa8NZ3GylsswxWkjEXUJ0dUArD+U3f2YyKaJW0cLGk
zO3ByrPXO9aRwQCu1DjmmUt4OY6+doqcNh1JhB/2qmB2QqtRDoh3gwytZthjS+uq
94YXpAlflazf0S4M1AyDytny2X1zKndYxf2jBUkhql2nLt1F7M9xoxhZWwphLjsq
0RLNWRt1uj8HVQGAtkXCzrsz+lMVc23Pt+v56qpqdRQ0HgLYND1wVluqD9Dd0BRs
9O7iRAymm939S3QEgH2WE8OVdCiIjn3kiLdAfVvk7mPIADgBO0jqeYuup362Zd0x
Pvh+wQFVcgmsL6oXPCXxv7nmyWCARJmMBljyW+3iRY+iBoVDlCiCZQmEN9CAjA/E
`protect END_PROTECTED
