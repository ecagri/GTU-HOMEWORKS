`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SGyiVjw2SnaLxqQ/g8nYAsyQ74sHSNp2D/zSXBYvxTrZwswzsVZ+EDgyMwsia7DW
1HJ94lJKfRrXWUpGiC86cLCFjgSBPNJP6WjYi8wMehDloKqDs1G4EUBVUmalEdqc
3LOiUv+mnpau2D6pZZ8gSRZodauPCUnzXIjseHJ+YGBLCrPoGLx/wEEG4D+KUUH9
Yp1ckuHGMD0ib8FOOf69RC0bCJA8EJ4EsO0oAWy8Ih2TRisLpYOP7l5PhWchrdHz
V5rwn5YXPkn/ux/jYb1Qj/+F1foP2IqRbDl4Ru73A7IPXQ9hXnpLCVqJdjYBa1v0
SeQtKNucPfeNuczEzVu4OsLhyDhrGYnYJLAXcQg4XUZf9DwyUpD/KkKu9yADXGVe
55/QmrvFZ9jMFd/2Th+w1bxHvfFrOGe8/Wk7LCr5C/z2nVN8AMPbvMDjgCvy4HwN
PdR6WUlWaOoGjaC6eCqqMpKk5Ve8HUW6gzUurInKcxS9qrnX3CEyaeaphZE7Hw2y
NdVA5MUbuRy+E4LveGMmnE27+Z9Y/dyYdAjCK5i97BZvAQWFT46M8caGblw5romB
qW0fJkuHVOIK1+XfHJ4maSLNHoRwndk+hfwuqDAJkGW6cq1lyZxSBh2q9Brpo7aP
pM7zJiHEr/bM2Qn38b++CTuTvxKi9UUIAW/OEF/7899QWsHhoghx6IwrEFdQ69PU
k5kJuvp/bTunJN30XMNqhrJlbWvJMssPv1xb1mCK+UuWRL5IqhwMd4RJM49uSUJY
x5sjm7N7OMpcOe5D6jQbfRebcjgFiA4NMVCRPFnek6TSX8CHK3oLu18RSrodqdBI
DKJW4ixDg0D+x36XiOP8EhzGKX82RJAz0l/SazzmQN8rRbqx68hMu36Hx+VSIG44
kyuNCr8sr7jcXwGA8ShF4ANtbC42K3RZL/m8u7ILM9DYD5Ff+RSsL5WmPn/xf8aY
4rIEn3uTtsZ0TyOK9BHWYoAd4qhQj9Cqp1bduUMTIuOd8m8YGU+YoB1s1TK3KSZB
b6dSlWeLRpmWzHLfyWIGu8LE/4S0gCPTO9CFyFRVgBhMmNtzgz5zjO+FCO0F/NR7
bgE6701Iw1BWTNf2Qi+fTlFG4MU9FlzNp879Wusq630jXkERxlN9PJQeZjDsiexY
0Hkvg3nap/JsGs2Oxro+4FSJx+UqV+gD1iqNypBjk6bd/Exg3j3kSKLsgOe/bvl3
gaIK9nk98mC0J3Njd7WgTkSub40Ic7oa2ZQ5OTffz0z+HylfWKkEaT799z0DsNvg
WbOzcf+kj+h/irlGl3lVb0fa32YTjGzqMcQFg5Le/gMGb4go/vJfn0w90wV0aoYH
rGG62dIpQldN+Eor/5kvmpdaVmKed0iYner77VE9sdVSQ+qDPd2blOcuTgnfDVoA
TWXPbC/5eq4v2jpsX9RKiZf3mGNNUpJUl+aVkTiVcFNMkz/5BicchKX9vQ456+7f
PxAnZDR9qpyjvMbJ/WvlZmGU3sSQCTKXMdO8Qi6XvsbSN0Ape8X3UYAL2cr4LVkf
0ELzKRK1gmFjJ5+rz5N5xHdqG+L9S8vtBCrpiqLHd3SV6YHfXUR0TICKijGrGZJe
OcGy+9cmM3MF7qPtqbhMxHVTYdynbMEv6lgyhSIlwBWi8RtULnStlrkHUscredjD
P3n+AkOi3+x+TYJptPUZa6VcIf6kmL285POljOebVYOjceX9aHjUxbDvLqp75SX/
1kBhpmPHepLziGNB+a37IMR85P5fULssjKQWeEHvxLWXqut84kDJqOf3vYAGKV5R
375Xs0w0LDqgND97p/pg+lbgmRBnDozw9vd3oLtEKmSIpY2GQNiUu7vJlZIakegz
AT+Rd8o1U/3KiJwNt2USZkk8DvwkQerQrGMZoJDJ1Fok1awOFCr3TtSRjZI7uWXm
WtNa+gcfWLjv0cdA7cynRdvCvW13cBMo8aW629uCUSsoEghATLUFe089z4E/cmCi
PXV1EYb5Xi+ma8zogQqj9BP0X6dxr1PmKCHITol11SmJ3FcZJyyQEfULJMD+NTOE
uN1ObrWgfnU7yt5NQhiQ5rhehyXYt7kUyZrqfSu1+KtadvvVOww7z4+Z22uduj53
OxBhPYmmx9mHgSLPjZaJ89016TZTLwjmOiQ3MmW9jXbbubXlM6cEOlCkudqdgMyB
BI/Kdh1m0GietVXMHpU8LyUnKLYJrsEYCpJdIBlFCHyZG86XtIp/Q9bgePGctCDw
uF8Kdlqc06U6aLAFp67TbRxlCbLH5YTmnsbKTivRYinE0Zz90m0FHVeMMgkUoTkg
rbIChDpVZkxA6kfvgduvHy7lYJOhv6sebB/uLtStfMAvjR8gAI9ljhcZoxNL3yco
0wPTrMZnnG7xoWYh1XE9PEL4xRcLYVtGF6faeZX48x57dlH11CtUeaMlZoO7J/s2
I327hO9Urzaaq2OKVYRTC1++icKEupORwy2II1X5OYM47kPdqEz08URBdO57X93K
FuB7LGCh5jh/wSaOfyZIwFoGrWmXMovx2YHXAG6qhnvgThVkKl6uuBCCkXV2xTYi
h5EmGtHAmRg91CLhpslfLeJzXhIKWBc0OYOYuCrV+sc7v2s+MfjXSFWJzWABFI/e
Av770aq8v1p8euH8Qex7B0+VxBg/WWpPiz45NlP1wMNIVox6FeqFTeoFeriVFdAN
nDc7nstMkuPYTHuQK2lD27k94rtL4xfmkPRSbubouV5N3ulAYEHCFh08MouLkMX6
Anvn6g8irNFTf+GYv7bUYEHl+vJmAzUpQQmvyXgM7ast/jhqDPdVG1qIRnquUZKL
mRSR+nKqJhA5FYYVXsVPeLpo+W9u7pm4Fr6v+Zrl9DzLyC8T+AJ39CiejISB2DJl
Lw0WTfFsFcqfOsg1HLjCXzo0l0mNeb8EG2e210Zs6D8ctgpsgUZb2u/k9j2uTvhe
sQ6hEGwc0xWcJLyZicuOrdRsrS1C+4dyN+4XC67qvov2IAU6a+kxd6zBhUtelQC6
TDPLJTWGzF7P7/4+TRUAIyrSZZ7wJwhacJO9N8JyPPCHtLuMm5IFvA80AvbvhXEr
UpHSkuZBBacAiVIPejxD/daRSPIQCZwChTGo4dxsGcEE5HBU9UA4EzYvgwqK6Feo
5KQTVi53/PSj9mvXfwHkuwJQdhl1n9FpCK47FdIh9iVwI/PZ4YmwrMrXZXMwyqZ6
92VcXuu8ifCmxpT7Z/r/IMT5dW/yXg3NZ9w9emyFpEeI1JCVVir5RH5MBJGaLMC6
92rjlohk31ocYCj/Kje13fE31F0CYC3iNUeAYy2xDMTMr37QlKNrDqkfopMVAD0Q
YCgF7CzGPq3aCzAKFPp8/4yRrykCUZAoMjPuuG7/VEXFHdluSCnD0VcMZQLpYwYx
t7TxUgmj81npImbd3Pl2yh2qApj9qqt9Sj+Y9TSVGqLosP/vY3bF/iq6CM9QskAG
cIiVo4yEeRvfsYgJRkIdm9jUh/nbvm7fB0keb9oxuCXcAQM7dy8DmEDVPhZY9aVY
O4br4Gi1XzimGtZzPZok0S0hRNsnWaoXY0OZiRHOs4oiFiaieOE/XslrT9D7p5kq
j3u+y3tGVLU2FdhAwUKzspydGulMmPSt78emxozGOEBTRmSv7y2tuPgegeYD9ecu
KdeeMS0ZlrpGaiL76oCQPOl9GReNaXXmNwRAVvHRZMLZPYl3gWJZSn7PV+wlzgGE
e7UgvMa7YyeaXeUB0e4T1R+gYVhVgxvR0f08g0UBfldLTqxT5cE+gdQZzbmPr+qH
JoH0XwV9ygCE01w9kLJHNJocA/jK+SS7wV+nYBEbzJ+YO4lINVQQk2kiKj7vOKoe
M4Y1s19ggvmmbJUvvPz0MoUxDA3AD6GW5qWv2UBPyEVIKfp9vjFH7Iw4KnRvRdT4
4naDDL5SJ+x/ObUpMR9hNPozyN292aNBk3avYhGNH04IhMLpADbclGgmdRePqVQH
SBwzEK6da+xrcf6uS20whoydFsxkeltCdlzHLHa2oMwH7zXBXQMwuCYpNgWC0Js5
CVOjPNXn7WCbLEif0fn9LjfvSqwz9CgRZZfGnvS7qKOO7Qvmob59yc2bdbv5fzQs
jkOqCtQ8ipkXeREk2h4OwZQ2K0DS2cn83amPZf8cdptWjqx5D5YD8lwdz+HSxGu1
Z5Mdftn/+aevt82/nivU44XriRLLx0jTsPtXtoeMf9UKDTW+cSIa3Ia1HhFlchX1
c99snwUK+6AZ+wzFwQKgel5IKaq85AY+uUKuu1OWgATRbmpmKHsC+hFmSlpXyBD9
PqIe75eTv6RxXSPY/8yhgfD0D6jpdaIgMLROWX2kg62GrZsEmgUJ8uDAK2/xGpE7
c+ukA4P4KYRGkU6/vetAgEu1uPwtfwTjhtxcwHYKcK+zkC7PgnmL+pQJ80szBYPm
nFqgNiqYpXaxZp+eS6S5AKWm5YCKJxHHK8/hLtPJmn6gKNDhlBU2BAFie06WFdwA
VEiko/QqKggWNt3voCNtz52J0cVw13gPtti0FnAnx1s27HYeT4BsXcRMmjqRqLoj
FS6Qd9YjA64EFIB0jXPt8aRlTu1a7Hi4WP6HvO0LUXNjmWa4UygRjqB/beByTu4i
ncUSRRRlYIXCI7hw9MkHU/fDJU2V7PQml2Wzs643u2x4JCtxrjW6N0lxzM/gsJXJ
hKdx6f4GNsBOYigsypwfxr9W+MCsvw0UvaFOFSc6ckF7FZJ+vcU8V3KiN4WoCdJ7
8cdRq+9FtOko9eHKBwTn3Y1kwHMmvwBc4TxFpfFEFJQoS0MxfgORpiLoMt6ebsGs
Z7SClmv93UNDfeyisvuuJw07m5pzFN32Qt1mI2228YjlitrV/z9O6LTQqq8vD/ZX
7DvPXKd2s0MX1YSUzQSRxWQ3OB3DZfoYhweGgxFzhyKNHzGmiWKYfnU5mUaTk8H+
bkTjkXdza907/8Jus3WVZPE5Rutlv/tUiciU4H/eCiJHj16nyl7NgrutHO0Chpxu
OwDfx8kA1Fu+JtqSAr0IJ/q/JID0XBqWJR0ruBOSStRG6+xhSdgcOEWcBn8CODqr
TkvsCDmL6ktd+R74GBNCwa/gYRX2pTJ1QIFxbcqgYQXpdRc6yb2GXlgJhqaL7rh+
QFhY5sIEqPHshWADrCnVwbbTme8RjZ8ONSyZHsQPkwNgbkbOmJJvGD9FAehJoEtK
DMLQLYwlsKvLJHCJVdoCT1XtLEqH//QKAzRiCCHSvfYPtKof573MwRVO760z8WbG
7WI+/TEToP83ot0bvaCwJtZZjayck9UP+hbBml7D5C1lzMPSdzsd117fszFdC5wd
iPOV1VZXJb7q7QqQy+JP1UcYa/tj6n3GXnhODKWMYAOf3NfcQzylQS9TiyjHWZAM
bXuAxuWCdc++T4cP90Bmt/T+x1VVintNrNZQvk+D/T3Mxl3WFOpshxEzkCqnEbdb
zuOVi83429AmFX7aQTOf3BMLAuXdR6e/9rTD37y57WqdRVT2M8GU2nC8u8cwRYN7
4U7R7IhMNHODD9L2DJoPiWZYKY2hILThOe1Lmh4GOeuvvIik4rl5tFOmgD/ENCDK
/NKaMLh9J49jVgG8mu2GB2JgsE+lCEuw0ZAX0ol6l8Br3X1KketpzbtU7+BgNq2U
djqzFRWUDn3QPqq5gv0QqtwGqO4ZnOpMyMGrt44Xkeg4xXUNsFdE/mey07eSEibW
/pCvf9gjjvN2XCRNc31ZsBcKvUg+593P1k54d6lFI1rs+PiIHKaDX0hM2NL2c6L2
FfKJLLkEWyQk1KvTV5fAjqN3O6WtJRk5Oa4MDlgM9dHlEpiJV8nDWa/Bg/uYdV8x
6bklps4JifSkKm2zclZRRmGF+wb6Q4ToN7BRFmTA4qWN86/1ESOCiu++QFAYViEr
jF2dWStyf5aWbqq5W7mmWI+RXA8jI9hLyEW6d9IoCSAPhX2Y/5ZeQr76CGehp31y
+GERApPrR4W7YlFbVjZgBbA9AiaC5Ul+/KWyaf61M8qbHATICzbe1Iv8zlS84nZ9
tGkMfAD57EiD/OSBvCtphqZXLmMcd4a6QjoAdD5pkUT9u0firHUtyp6W1GsQsWGj
ocPxwII6jSzsUhF7mV+zyj7t5Tq6qkJIeI34+PwxXpUEeH/qm6vh2ZAJBJgRXnEf
EZwDtdpAgEOAfxiFr4AFAhfjJ+jLfONYiNZ+R1JFFosbCfB2D0N3zDFzsGgXFKDG
A+YXw1wJzqisi0JJrOkUdeWyNFbfeyzG3nEL9ENzqCJUZwmBEi8dnCvIQ1JKTqKY
9FM25u0D4/cdZoEVESeNjaOz2CZaXO3hekyk0o/Jug5NmF5eBW+olEBf0AtE+fXg
rHUZrS+6iw8zozacARCBhxrh8rS0D2+dmidGM+mSUiOQ1Q7cENyzS62naZTtIKA0
PeRwQP/dDvjoV3+oPPRLyNCdMj0K1JMeD66ueQMvdgz/gFHm6WqBvZt/26mD3vJq
bd/Xt8SbAxBQ0NcmL8Wt2Dve4RfDjGO+xpB/jyYfH8auJc5ELXoBV5efmjpDyVCn
VrqD6/M2q1dJr7ZlLk/WayjzdhjgamOv4AxAzol9Oi21RmuYt+xNNIelVpRDPV0Z
vL7VsgQDK2AZpyESlE8GCWJjFAoYjefmWdvto9ydcG7dre6rJdixXFAVpYj8S2o7
uSOiOZulK1pcXGkgLuvTdEHxAEkRx7p8bmWEz1Ez84TREbFnLfNGQTMOQCenozwJ
x8oVd/u5mXl6toF7Yu2BAlmXA9Vz1PYAp+X98fkzHpbvRiyv5v0PyIuQfGSuNpdO
J5dXPfVN+tDWqlgW6ImUBUqicQdnlYY5vmzN4KWhxHIpLlaBcz6s+4X9ctHj39lH
/ajGQmaAIvS7IaF1dGASp8irgeNO2Aa0zKRlh19Cu86FmLqVgIlVjoB3hTdkUb/u
MbspMBSWwakkip4UFwwklIHbu/3wZ0fTdQJ8rnyIwZWnztwdyajkTpD4R56XGcsU
/+90JfIjrscTVZTzwv7dchT1u17HvjRjoWw+e67soQUoSfNUdWIKg8xH6LTfRQfJ
TuYPdDZ15qqAar8dv5484jP4LaloNYyhGJmDr5Q94J7Cm/KGpRHsW2IsHYJ60FJ4
YAgEtZj1GkN7AQB+N6Y/hVmGqSWjNEB3K5Nf6f2P2EOnLiOUaEl1hH8vfFNPSO61
Utz+Z33iqFKaBGdbVuYfrxNuZEOX9AyDW47t0fVYP+fu0vvwup7i66W/Xhv7FOBh
1JTa1yKvbMOrN/1DG7b413qqgYmXd2mXCQOKbYGAqTFaZS/SysW8oEKu/HjkrAJF
6iZY6STuaYrDe/L2Ay58GjD9o6Xoeiq34QZg2XOp+e7NL7MaR5wnKLNyDBKq1k5W
WRyBjZAHrqzV+YumBr6QfSRA8fifOWVmXJdm9dNp4JKHKbsR3Oll+tfFuubJ1Ya9
89/sISHCax0k41Lo0Sg46JlFyvwJ3B7fy5hnVuBQxTZCDFVTsFXHrvTSnyW4Jrpf
ikTJzmq9x36RVVjY0600WB8dIN+xkq/7FRXolTl9thQTzF7rC5ctcVd0NJYfB2of
CwHXjy4jkn0Z3yGJYZDSFsnblnDoSgwgDpcXTstVX16Ot+DinfVFo9Yz7e5Jtl6J
p/zTbyHEr5yHnIJTKcAxaSsXF+pwuXyK02whsvVhqiRz9Qd1fYI+PWWZwDnWupNo
+9SIiJqrn2H5N0SdtWWK+2E1TIaexpitk9/qs59mb4OMzpCZlK8TzKTJzXtog19l
PvUcKsbmq14tH207HYlsyPkqkXRpOvhytOm52EgdE3Ce3UnW8SDThhkEE90oWTMu
+4DvoyCDj4OZhrCp/8yQCHlcbjfs9POVXkYE26TAjCmqNp9MHiX1pBAj9Xc+3xCS
fkXvauip6qwh7Q1mnr98g+7Je4vgy818KHgCdqHJXolmSUmxYy+aK5z5GuC6QL/+
KzL9aThvgUUTWN+91eM3mRcQqvzSjq71cqVPLafgmeZ6LZ3vDuAvFwRYUg01Bo2Q
W1Fhs2pGbDM0oDh4ykUDHFRNec05G+6g3tzBZ5b6NXTvApfSrK8tsiOIrYFLOvvF
0ZeQIa0ORBwZIU5mR6zS+9imS7WdOCkUjrOrnAwZ2VgXGM+xIuMSP83kmmSDjaPJ
MhRLUICWKoVqW2jJoqxKPExO4nrVZVLmkcMrQ2IveIuTZwv4wjM0P8SZI7jxJiZ2
qftZcx4e6bXKTw9jst6YJyd6lchi/OjqcHg9W1qABvm7fB9pK1wa1/GTXrl+aPFQ
OM47c5jiVQ2RoI7eAPqEdurFD+PoR9jActtI2MrgHHUdSeSnv85z6W9SXrYBxRFs
HxZ26xkPSQ+XTbqRz3e2ROPwhFT3xJAm+R0/YamHl1nsDDDfUekj1HrfFWcc4t+y
VNa5TyDVSLfQACyJ6fbRyiid8s+9NeQWvGBhwm71hClSVGu4OSdNsVKIRaoapHkn
18P0cBX8LB3wFkPFmec/adqGpOZ8EGoaxWdWfoNr0E/A1W9SFwiP/1rDePFuO7h6
Yb9J3GwtOrMK18fkWlviAr6vC+dwmm755v1gFe5r7D3B2AXUAuGme+eQDrBoCW3b
oynR5Fb8AR/l+I513m4MSQ2p/fwvudgv+DobsKII1NsYhL1dC3uKgxIqO91T2HRs
02yfEgk30Js/xvZIrRMA5q2XSeL0op3lLtTLX3DfhsxpVr8m3xeZ8rbXe1MQ2Z+r
fw4QTKDd10OR6/ioARuZOkrS6QjOCBFj7bvassVXYff/cu7X8Y2Vz2x/B5PYEZZL
FGmtCqBJUw63o0E8GkOg0guBDVFzGhQ0wSPfDsPnvrbaN6BBsSt7NCLfE3w6C+ZP
4nxeGXSSkpd0NEQb91Rm9LNsUpdA10K97gX7zTTCUx3ESZzQYj+7ume8BB8cwF5P
LjNsbKRmN5K5jwK1vp4VMR69N3I9xkdyHPyhC/f2h+oQVHAzaTgWs7+6LNzJPoJo
Iio0Nse+dXYcrKvvRtj2g9GmjOOhD0IQVO8OnN8JoI4wvDys9BmR5AahHpelRQsy
tXLh6xwLj2nbacc7jbl2OqkUMeiBcqK/u6dW+5SYDOWsIPwcsmH/xI8knMfEbELz
o1x5UwCrv/WvHd0SUkIouqxnd1aEbV5M4p2m0lN963iA6JUFqmWCLvQmmm9jlmNN
6o529XyXP1r91wqKQXQEgPGKaToE+gB4mybJGcwiLw85CJECRWo13Xe+4gLfhmO1
zkT+kBaGiQzqm9zZwPBRczkSTLgQ3/+wEdejsx+KSDqhjyHGZ7+2tWMOHingHdUd
5s7po+Rxt8w3nreYP4giS/t/C0GLqt7B3TFNqityuM5H0xZ3AncnS5DEzigEOvLF
JcMw08VXtwpn6tFSR3rwRB7KPW1FVQYD0J6tGVy2euiCtUnqeVKAGPxXAbE7IC0a
Kk982d+2BQeM9+VJh8lE9p0lq4hZBkNKlbG0Pg9GPFn9Ewdvb+j1uQCfbHGlt/wT
MTFR/C/OeDUHcoyzNVMOXTiZHVM3dxuGBmw/LitkapV+Tstn0aPNOWH+NikwXmo5
QrVEi6ZCX1CaaXtMNNZ0iLxc6Y/CNPMRBZMB9ANhISxbBsd9DldWZpTOx6LyAF6h
45RA7N2Mz8xjG019tJ2tv7uxtLaC2qR3Mg/N0AYAMEy3sIJJxwqjGrJN4KMq+1ve
J7h3A3o5fC9Q0knUfN3oqCw3WPHkb8atqHEbJzoFHu/6VKaqc0ibkk73LL8kipFP
HIs2yk+midtFPpA5ez/cD7tvXZzsB7T3iK3H3eSWvkXZmndEzwiQZp/90oARcvA7
naunL7EpT5Mj/+7+qCtUk2v0gzBHC3JPDRJoOeiZVkRjwf7xWM1D2slDu1dK6sMD
la/iPNBiTjEjfVHasmBF1izRfHQCbAA380Bj1amMwToGO1oXvPIr9tIcPAoyiQLy
iogweOKUEDPvyTWB3lY6eGHWQMuilr7gCL6eQh91MwWei8wRSbWpN2+g5jpDv59p
tZa1e/TvJvbiEBFDOcNBl9JxsEFbvTVlfdM29FnMVBQ/KgwjowQB468PuypbrFSo
YRj+sOLUkraRhmCAQEbCSrnwR+k0yt1XZL+RDwsMFnQnkT5qZl/93KLKK4aAarcX
a+yLIRKVefEvhK+i7mBhLGGLx+73MhPE+61uyLnI7ECi789j0UJtFXWHqQb3qNIy
lCi1E0JydzmLKk0sITzGyynZc8C+x+OhP5j+Bk0/gXX5J6cV1G6DeMjVGhPXsQfm
Tdq3QczMJpTW4vUfHWhJz0t7CqhuO/RhDWMvJRSdYID7sQMmUeKsR4MYDVcGeySW
R3yklClrCDgKQnEv5wzx4gE1CWSgsA4h9SK1Z6Diwx+5KsK7hYiOz8lYEvGWZEte
h08wOI/4nj83DUU3KHDPg+umh40II/Myyp0ThWSAwWPKKOBEDQD9MHI/gzDFwdjG
ixzQlRnHayZ4qCGWwjr3sa1sXWBsfI3UD+JI7KnztVln8Bv3XbI6p6UJoRgQnnca
SY8fixsXQi85LA6J2QKhcPBQzLXAE98F8fPJiN6DUJXPdt35x3oKwGZIJVbV57II
Xo2ZGKLKsSSf5SBZ4htSwsxBHqJy5brCD1+te3bdng/UVovpUa/kltp45DgRaQFo
ROGR+gpIa9VK9o8uFWsHFUedgbHBno4Vh4MmmF9huF6PKch6fVFiujOlcsIelPP0
HZPdYTIR+6HfhtP9cbXamRygE80d//t8JG+9mV9b4TCNW764fnBTvf5XcF3QaeIx
t+VCFGRI4vCKabz6fzR3AM8ftSzoxwxEhPi+JpDOY+hu4FbczZqjQVWo0AumTTH3
pqmzUTG7W3ibwNiT6x8rGqOulovXasCcidUfS3JqkunEXkL0YnzQwVbZybzJ6yYi
6XyvkRkT4tTQTqnQgokxYMuzy55f51ytpKPl9H30kj646Jf0BMkdCHPyvgX6TX7c
37VV71W+YIMgH3jQZsIEv5Q3VSvius+LbjsHFC/tehgW2VumoH8GSbq3zXEBUFb6
9fVkwFqF2XJnxg4tJVwt6KTU+nkUmytAtidxCBbsQFRAcg4nDPV/28FqdyHVJNpd
RzTzYFr2B1nsgU1RWHglvyFKvmTGu/3OxpfAIJrVzfQyvmnWjS0Vto5EhAx9okXP
lNJh/grO/IbeivmP+5BtP2xcXaWuM2469w0dWumzd9RLokNEax0eJhntQbjLve/g
o1c65cm4MURXH0fkrnL3eFvMhyc+8qaqJsmz2P5h7dyKSO9E3j6UwQ9nxSiraO9T
CB413bJzjzSPAdNvqcF1upUj+9rgOAOboKU0Lj1jPHLp0vp8AljdH0lJidiZrZTH
VgPbEQz82+VnaBEnyZ4QjTWxGMnMSOpb8VM3K+EeT/xFpvxeBjkiF7l2xFJFjqrY
NFmiSoWRd3eduJgU79puaWCniqF8vUVoVNQwxOWu/hAi2H1wrV64cQkwrcBCLI4V
ZIIblzHjv2h7hK2jxxMMoudleDCUeZJQwPI+6arZGVnR0I7lNyRqzdgxqkzLStRV
0WLdAvzw3azf8NYl0UUWvGNx9zMtv6NcXrQV9S/DmJOWWxl4KhhhBkBUdIzDCZ6P
XLywUjLcBekfRtJlg0d+kNpQjG0N7HqCIykrMQvHfoDk8s8qtdeJrRBF/gF/ObHy
Mkmqjc0w3oIS+SMfTaslNj1RACjCTfDCMZtBKYzY/et3PpEk/JhOTPg+BD58EsIU
5/W+/rqWFYmjFPh56HfZxm6ILU+fA4dGBFUJ2abDLhlDdzeVguTX6G111a2etYnN
SWYmhVTYqMhbjomhziIUIOtRlsVOykDglOKEbzTIdZFAiWNhqm/pohhkd8bbdjzd
r8lyL23BmmAN9k6Xdb5XhP+XpFYsZo6/9iwALcPi67m6QvuWSHRWLa5jJKQr0O3n
0uISEB/4OIA3hGvzJfVgLF4CiibArmcrbmSMhBa7FJRtdFt0AqcwHShy0jV9umRC
RWTiQkeJ/Ehu/ozo/r4B774VcIjEwwQy/IrTs/rnaKr+Pt71ezUhRD+Xv5BRz3nH
OyQbERp687BPNL1By2qhBKRY34nIqGwOOiFqicwq+zumrPnTEiLSFpwYlNQP1aG/
fNNhTHMGFu6ROAQT4f+VAQdRv94+w1AhT6rYk0QLmHl+oCM4DuS9Pl8/nn9VO2gS
q7SLjgvWkBRXJ3O1hnP7r+Bz0FC1poCnPCkqeXFC85pV6g6xal1o+TKy9mXic89x
Qif1Y/XTWyhdHPPUqMehYZ9SxFRxFFSwh8+SJcIPaJHqbFq215w73IjnDUZQwh+F
WPLGYBQLswn/SRXXe5yVeedVKcnemztuJLqm8VfO9nPo34/WlgGLjLkSj3Ok89Mh
T4LQLbHHmwDBRi8Iw6ZmF6LVvGy055Cytgy3UHAwpcP4tBKh5uZK1Gf2MAN5rKIR
A/jdrM3mZr+P3Jv/dNPGTmApLZuzWeZH2ebc+FjKhwww136dpPU0/ygJU3DBtoYC
rn9+ftTDxAWVvnj/iqWoZkjOtabAyoZ7H9TncUCkuaumoD8FyamXuAzyE5alE1+k
F5ijtE77wCvh1+4b+y+Bmz3d/on/+7pcGnu9jK6FzTM1ehgub0yAlwu/+ZwrJqHD
sW2SoQXKC/1Zxekf/dLeoCB5Rw7a3NF+0uTCwUHr7bKm4f6SZoiY5zh9lTsb5DsH
PfcyuIZGdG3tOuYq+tyrUg+oYRx3aPrYJJrsi8mXFE3oRqR2pAfkN4FmxUZa+QC0
+0hWr4kJw5c3EFyWtXKWfNhlBVJ/v/svLapGYIgrF4pf/3LAvIkFcPB9M9Ym3yjx
dl4K3eOz8s/1VLhLQgpsspriy+onzU36pQ+mD2v69Xah7C7iDfSU10KEYsdyn04B
eD4MO8Zm3SzdARR3pWbNFWfNBFbngECY+VMLa/tSVpfro+RsswKXyQJENTh5hGXU
hRagOK/8bxhHYq/PPD7J8rO8xr1PiVSFmp0qKb42vM+wPReywAV8f3T3QkMIJZus
lypmAaT4WF8vWZihxYqQaLlKGYbaZfW6EwOnV8tiH4eCOS/erQxSfeOKrheFqC72
gQ1i1URcZ8fz3n6rN//IHK+nhNX83862qzLLaGXK/u0UnahvT7A/xHJAtLwq4QRM
4OZB/3CGvvixpD36FbsywnRDPF4aKBI8zWXpEoc6iIqzZOKDSLd7NgTxo7dOCtlZ
ljFEX9TFPHHQj2bJd8iUO72rm5vsDxfDSEsMEGOgztOCiybTj1hAV2b5paKsZ+ZR
f44+fzHcrmvia2H+QOc6NIX1zlZK8O7kog7ixj+Q/fE=
`protect END_PROTECTED
