`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bYk1jzLca3YzWRwMjDCwkKi4HN9PNHDK9CX6AbdNG1RPzJ64MS6BKIbuOQkdzRN7
UM0+wurba6UCuEKqRfQXXyf+aiYgpmJJFgpK4+mffV8ADNO8cuS8q8Cc+avRRQdF
OtK8LAsAkLqUQbklzcK38JcVAPPhqETjnnM3JR6KY5zfmPEaIUBflr20BQmM2NyM
FSeOGJGHfWZMCn9Ygxf1WzbrW/etGwP9vqOj9Saohiu4WQunynP+4Yfd2N9ZtwGg
5FITPOhjoH/dzPGOTX5TwcA83StdJKeR0LXAbnusZd3YttJE3sgpcKsirLvINAyE
LBCaQNK3I5BibAG0EJ51VNncSSJotXT1JZhGDX1OSZ2lSbdMj9WzvoLfS8EEeTAo
nmygc5klZ1KebyUecVD8uQ6Hk0XbT1eDPkGllmwhQ4HJHoTIzXV9eLMCqGpBzuAe
l6a8MQluOOd7AG5WAZxIZLs6xsb2jAvJVoflbJ1lpOR4g4Jetuc/cazZ/wJUuzX9
nBOy2mSB/lAt4nlXkS/Lw7hlpDdtImNlg8wrI4VNfqPCjlQXn6w7n3094uv7vXt2
MdNDKIVa2czdadM2S3Rx+70g02kn8gfrFZmxQpfPI9erXrWKXoeu2U9QjCvMK6zE
TUYvTXG7S5xQRWA7yq+RNpcr/e9i2j43oojXqPoEyyohIv43FvUV/hL5upj0YlM4
rrvdqDdFAD24FzuA+oX9sirov6EDRPnAkS+16doylg5wacy4lu47LEmV7u2ElAmB
3THd9hm9JRTeZVCyGMh/nmW4csKWa6J84rQbW0b3rjzCskKBnbH3P7AI0UQ2+s+k
DrzEHH3cLshX6UxNSwiQMJ6ZGTn+jQm90Ea/nyDq18wF/78dygTbQEOKmvnrE6F0
zKbuD/Jp4Spk/CUm81vH2v7ON+DOqxRpFFINfAFyFA/EsissvhRuBhUwlW6V9oa6
B8DAHd0HYDZfWmN/bfh+5bYrgthb13biihGd6EsbPkxjfQqqN2usbYAVbf3kyaod
hAmiJzLH21hAmLZoSE+pzPPL3BNBRYOKbPI1NhfSv6d3AWYP52B8k8iW7M8qkrj6
R7pimA2C8VoVLPPGTDeMHw5dBbo3CY1WQoL5oiTIItydR1XhvRPMh2T0zDbw1vPg
LeIoHg5vLVEOt7nXoQFw9Byu6gIIRr5d+Ke4Ex8WPu2cHJTG6Hl5XUjVxN0kdus7
WloIXUtlq/7Tt7eiH9ZU7Ykltv2K04BIVCgYJ/xOyXQ39WyqA0vsa5nXVc/ka+MH
/LyZ1ko3jpnYBRWfD7wDC8Q5hoXWzKRHaOuFGFzBISQNZxeqjqU7P3+MhvsFtS+K
VyYH7W84JBc2GDYxAWQUdA==
`protect END_PROTECTED
