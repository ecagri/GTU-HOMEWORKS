`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bT/bYra71FpGfAuQWPUyZ3hg2+0cl37Je3krDpQyCLNQ/FDVsKkOcm5fhf0Og65t
LRRJM2imi8Mns/58q9j6DkkflTJMraQI4rGBJgR13xhOFYlpgYlzRcTlO9eLF5eH
kZRivZ3bWQ2krf6tN8ON88mge/DeZNlEerrEZ5nyewb3V0E7toAf0m1zqTCAOyJv
OcT2+lA/DqNCImI++NWSlRsGZ3aiBERoCFozQ4+8lsYgO9+PS681CZpiSCue9uHo
WU8IVBtkB2Z8pslGlRPCnnhbjBJ7i0TgAXJ3Z+h3lCO+brbSvwF1EMFKP74Owe7L
bKVbjqcWASSp3QGucaXvxZ+QsHSqhr23sQZdgVaEdArRt/erga/hKQcGLkgToFp5
CeevnbHtPPyIyPyLrOc7evfjdibbftbuGzOKCrE1jfTAjAcJK/2G13zWXeasfpnw
mHykHJbZndD4wfh0KdL74qtiPG8V6y2/w50AntFp1rkjSlrZwEMvBEf7ylFug9/+
3nWPBNqK1b2N9UtoCnOmTkOhFUpcPCS1BwK0L2Q0VlD2JPVFICDBA1T9Oak+TBOv
7Sx9NmQFUnBpGFp3JmcaKhgtOkvShQEF4EK+TL5IaZ4BXDveW1KYx1yEc+UeGLds
`protect END_PROTECTED
