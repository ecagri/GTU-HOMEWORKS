`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jRF4jya8d52T3PeaUwUvWZAmNjR0mT4sfLC1dzTWU9vchWdB8Xsin4HkmPMWYPX+
Qmj0n2mNuiR0iCxUbhpOvBUku2EhKKMtwjRPO0VVQYPHIBJTzTlENp0rGqr6F34M
C0QBNHJHnnfaI73Bmr+Myggm5q5ADWHIIkiEROtjXF6/IeItUnfHgs2vz4nIpDN4
ljjvfUva7aKDCEfuQwIU62yoqEzHAyPBfgaVfp4YJoKZgkkdRJKmzwsx4hgD2iIA
4zdm/SC19RFjF2Ep4PpmvN12eJ4iYykQgu5Wo8Z1/lIjBrYH+fso11ubssL1vyHi
lf+EFa/0m9UzCozSjvrIPjQpUty6lXRk07XKZ33ZBH7zI1RGETGGU6UIIPh/BI9x
aWP1qlddWLOvDSQy8xVdN3jsb/eipkfQSY8uOVoYp+is0Ch7rHKFiHGOPQrIWRYa
xvy322lfdOVr8gI79D8tThkbeJ7hNqFpeZ1depO6w1Sjmvka0n0jmlyXHSfFw/iS
wzmUFKHRsH1oRwLbjr0mUmKQflsv1NaS6AOQfjm5JNv1O4+rrAB130tdNq8obzjL
6mE++7kV5r1HWjQNJR9ltawzbabQmWPmKRUXxF22dfWSEKw0lPGEhOxupIVzePG9
TD5F07DyI84htFsqCt1lL7YXUuNAKkRk91jjHBdSPQ09LAbuQxoQgVXz0K2UR2Wl
3BqV6+8oU01ROck/8pFBHAumJ4yP4mtOHDh2ccIwnIzdGz1uzacI5IH2SP6tSea0
xMpGa5eIll/0mPPfUXDgwNATDmU9+B9aRqb8ceRpvgSfLBqJ4tVFYENZaJOC2F+A
ioQRtJZlOeVMWRYUpPa7BXjQ5mR4bGFMjgKZUJXWFg1+RGIZMBrozZWYM+cycGa/
9TpVYfbDNZRy5kJIt+RluoPhOK+8QE4vbIZtscNNGbEOVEzsyMUH835POUQ5IkjH
kvUu0rx/jceB4GaaiSQvI1Bw97yyKg+sGwKHgN8LeVfrbtKynMfkhevE9JMn5Bq+
`protect END_PROTECTED
