`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cW6dT3TM5vxvjpJ8pdHNVaX6Ej7oCBsp4oxHjXMO9GkggP5jUUs1WGL0+iO7UUX+
ifo92qhAZGVzpyXHKetr/C2Elkvmx6MTh/Thng3QgQAx+q07W7oFqrT3T9fwUvmG
79Tw/a/nWtS4MrBAcgXzj67NtYRCgATcCYRZze6NHIYMJ029Jy9ECf/YPsWA4lqT
OtMQsiIAcsbgvdWyZXN0I3+ReNad2q3kHhXn+VQn7Gihi7wURciO0daBdwqJ5oSl
cFRD8z0sq/PAoWdDWXbv1788tpw1+cPUPAdlszFZJRSwBcW7dGWqL/skyn2k5bDk
bnzWJb+xkooPqCsWMYYdqg0nay8TQK9Fgq5deH0cF29MwG//qsTAnqQ1MX6OJCHB
r80zdYSPnUoRlj84xj0WUNv+JP7OSZzRbMRVdcaYpQBjy/S53rqXYnoGC+A6VxWH
sTTAKFGwJw/xbwSpY55El88S15xml1Ubuw1FIG//N+N5x4gCoYjNIspJCmyqtAlY
/Somurbk8Db1mbgyWvlxmlvAq0KoDK+5VxLbMRIttHj3w3k6nNWFQ+NmGI0K0B0t
QzgSh8RivCAf/FPyv6BLNMTUdzvdpTTsZlfYL2jlDR26PE6olmWN49hyGicA0lur
Qa0TJ28GICjNy11Ufjfjmvag5TUng9W0kEHhLV//YnwPTwzYoIWxHEHDpbz4wm3o
0z3NVlrTu+/XrxoJbzk6OdTeQLeRzranFcOdKrKNFQkr/lCHo2KNUytnaZYhMyj9
M6AxqzCAxA92qAJQ2x8/bVsM5Lvnoa57EK9K62bhPFzXCT4s9A4WVt5Ue1BlSx+C
T+4xB46nk8KDh41GxW+BjfprNMopG6AlSd5PIWYwKMT9UZZPC+QzGfiEusEklqKd
OzoT7BwfymAaVqnBlkSeOicMPcZ9UTGYuJFQss9OYbizO31d9ujxXIQ72hqeKEV7
M/NPBunK3DOovobw3CatYny+8sgz8GzyTEThmgfcSLfg4CeP7mG1xSbFG8qFDhx+
UceQtw/9PY+ZQPz8kFeSqI2DRW99SJOwinVhY9wmzBsR7KW2v2M9UL1LVOcSRdgl
yPFFwLWwyU2xvxutF8TwCK4b/pczaMhq8wpKAByU7bLJwCkjOFE03gz7YZkhcWvI
uIbFiA8lOnzXGJqKDtMoEVccM1BgaRKznq3CSnTDcyPFSlIl2sES8z/uD2k03xws
kMt9mv2qwuFdXzCMUhk9qM2TfRYU4Pokdv/T+C1u2BfBdIcr6rSQKFJEK7czgMww
cIY/5QzFZIxdZtbFUuijlo7ELPygfIih9LUhDfX/jCQ+VL7eWjTgFKYh9icUz9Jp
Xz8oxxxH/PIlqheVSc+qSqEFTn4ncFS84fP0OdVVUgqXpbWxPie3icdm/x5iPjNz
oPBGRSL3UaybPKjRwAvjMILPp1hNmi4nQHVd1wWTvpnakyUsQDLkSLF0oKkgdRUH
JufQWdLmwCgeZQu/tmB+4oAvacJvgY/fMI85gDxOPaXwlQgHyP6lLHYp4lE+elKw
uPjTK61S6Ir0YAQJqOc754jfcMXnhHTFM96cKSnErLo/IZqepM66gsKzWqXXRRGD
NHS/IIpKdq8JRxZGuhs4nZHcMdtLltbXcIwiGqupnhslDWqthGcLUyTFpkec7V9j
Kximiq1FbPCemJH500M9Xb44NT9pVUTi6a1LFZytnKuLofiCtYk1lbuTA9Oxp4gE
2H7pAaRnGSNFkTqYUGTagkCtA/kfRCtX45a28KjnS+K5getH7nsR9/BNqwwz3KRG
+8zZKodlAcfYwmi1+MqXHvrJxAhUgCXmmW30BUpqncG3CMLPq1ni7ihfGk0nrxua
GUosx8VPoPDG3qdg7bVCm58JWX3FRlWvTv8zbwwrxZZJw5Ea1g6c4mmtK1Mrc0jV
ehLJTYVRyLSB/hjov9UmddeOm+j7wQMRIgk8+5Kdvbej0efAMPwefwRHqQnTr58O
iuh6StRs326UfCy4qD4DIPpEbcFZkm4j9zZFErKr9gSdWmjuHswBBnqn7VI6z58r
UR/APxh7gCvQKuJ1ER/vVYh0njVEtQTt/je88beJzPnu5EnqbGK+llkkXnNqYk0o
fzSIoTPV+54I2z5KxHiL3Okx+3qpwNpZOATzQh0FEu3AdhIeWWj9T4XH3DAF25bk
Zj5hG34ZvhywQidkFiG0nfePHL1gctywSHN8I2+wc0z/QRE756BaYHDGUJ/Gt+DU
Ifndr9fpWQBgtl2d4JT/d0IsB5BSguZKRnjQEbFSSAmmvZlZ/ks3YLbYWHFN0ux5
rj2XspGT918oeg4quFOn45lz3Sg2H0x3tzpkC6C+z/VP0vb38HlrIaZJVdwvNxHN
v/vT8++sOre/Fmp8BIC3PSW4rs0PSHX9w99gJpySA2Q7DHmKwtZeE/Nel+FB6gRB
BgRL+roRim4LyNP2i86m6KzA835R9TJoZp+f3xGvqwxuYiPSt0Si30yS6z+Knm0V
zbT0P5TS5DIFBD0cSiH/ALJe6FHEt2tgnWApJutlghSXwu40aLqup/BMTBv93rXC
CSN0JYSsj6MtThu9QH51mO81XZj4YK9L1SwPkps9BChilJDZb4PV0ZrOJPsdf4rw
0F/5Twp9S+4bM6f1ekxVmmH75IMrymTDdV4iluFG0YvJOUpRKa6ag4Jr0ZFv+Jne
cxXqdrWSdSSIirbeXfWFlCmcdZol2gwL6AjFdBSk2k/lRbgpLP+W2S7/RhT3L8IL
n17hAljKTp71qhKaURPwbZ0hDeYa2ILZ0uKz1FKmyBwXz+X03m3DgBfRfp6tLfzL
oF2GGQip3BccP9Qyxh5N19FMoCJEM36rnViqdz/LXYGUxIeeZ8OPMwkm+skQEFH2
JbC4CH0G5TOsUZLhREYYzERPxS/aiLnYEjfComR8ZSgqGuwe4Z4oTSHGQHin8A04
uLfDJkVDVRveRHvbTKCLZ21ttOE9wKRJI9GwowL2nSq5lfPoJP98Rgmca3HaY44f
+zwJvoLjWh1A0X/aaEEXA5BsFY+koogkXRshh5r+ZOQe6N/OWXJkICIfp0LyrE9r
n3gOapBTYLd4TAOhZQ5bYHGbQM83PP+QpYYkCAQtJHbjnDdwSDZW5m25uxdS9/xI
qbBun7Aod4f9sliJeZCoUGLpGh7AcJ/OVX/qVyXABeICwUWKAacsA9jFqBd69xzF
0mvO7MGc0+SB6IOAw7GisP6tFrryJC6RpmGOsbMPBJsp90+JlPx5O/j62ZQGFtxD
F51KySCdJEjNdW9OUqT0Uwn4o+hUjWArikZzLShF5UUCy5ODrM09l635gri/6pub
37Kb3fLBIErSRHU1O4D7QC7WeofLQ/q7gO+D4Hecw1HH8daymefKtYAWE/eHhaR9
YRVY5Q62RE9AZ3uPBfs9cXs718cl52SLjX0UF/W55N0hUbeXQ2fvsYMFO5CwAyCq
SUUfXHojiYgnaADve3XN6p7ClYYDy6m49kAXmnEfdKpJzmFK/5zN5m/tygrN/fYL
KU6HIdRqcwW2Zy+rxE45G0dL/UVB5i7gcsebPyUism4SPLuwthYnzgb5QjgpcekT
PNe0wBayGcjjo24lHY3WEPg98tM0dEYWn4VK6XMZa39DoPYsfwjheCRrKx2gUBtD
qZtT48hhwDSC+u/MIIa2prp9nIpPIBv7puFv4Sgaao3NNl71orATMpbYs8+2n0nX
W8k3C5gKiPQXl7BwmfJn5SALd4690NseO5Zv7jBFqltuYYLd1ljUcuRhX1ImE0vS
5fqkLH1VtrucG/nZDxuGcYuheBHfU+BsfH1MsNcdyb3Byhv99/5yVuwO8tuK7nRq
cXnz+92IludDIqAd+enBlZ2BUqUVf2dlVkIUnyq+ftP7FrwXFcpUa8bSRNVFQHUv
twg9D3puLrYb9vJRdQEJgRaI8xQA22w749V+ThxXFyZnnOTqv4j+mrwFTrQfhUXj
tZYpH3ydT4qgmuu4HOozjA2qidrOYbyuX5j22B7hP+34Gnga2i3Clsjy0j9iEa0d
ux21W1TnYoMZdst2cDGIbu3uSRtSo+vtSTLkIkXnfk2QkNn7t+k7RKuGsCneszmP
jwmtg5iCMBnN1v2+rXU3YxtmVrVCxLQ0ERnzRKtPKS5Ffgug2hQNJwP4BxiiVdaH
dQlUkbLYQSwk3coPExnAgYEp/3kCJT79/pohhcZXQ2HG7akZ6lhLZ/QOuAUrj3aI
zAeunSPHb+ccvoKZ2S6HcFQPfOPyXtbpr8W+x/wRjiAzF/KaSiiqy7ALOoxKDDeB
NME5mlURMEq5br5kAQwmMwnQsdNrPDtT9RJhlXJSOLVF3UpPPO9F/SyMeuOHPzo3
ulOUp1mVUmOtZwztyWwUOxF8Kcx1j25PkTLSS/5iaYl1RXiXSBkAqHRwHlh7mRON
Zqo3BP40iz0237os7BluaeEvfc1zXFTg+AOjhbW99CPSTm8YdqQQWGOV+Ux4p2ZH
86sCimsXcHDkgY1b+0eJ6W+pDJjxtrO2azx0YiQy+WaP/PXFcFcZK+fPcc6bxG2c
e3ohtxehRNiwBhVB0bMNRiusAawkPjBVYeIQ8AkVM9FLaBJd5AH3PsM4JRCeUTQ/
CdVABpc0iUXis22aEhaD1O0YzXY74+JuDJ32B/2qyo+b8jTzPk10l/S6u+xIcDjT
S55l1kJS6WlRmHxYn1SQqIGVVhXQHbJdTmeNEg/Cq6i/hM8xzuSs5f30pVzlosCR
3P31J+RZC/wHRCtuBW/byk2ZWuEkGZ7ar63voqyhZwbHAvU7gucjZBHlnXtzfqI0
psb/U9e67YlII8MTs5E8RkOeIIeRNsR+4jvx0qgOz4HDNA0cEhzZE8T/LUFCYJQs
X3kRrvJrKnyA7PFDJeNbK4dOKzRm1dGpTdEIErzY++6yD1lPH5G8okiEf36DjNi0
dCA8qrACYlsst2rt2b3qiYCr5Wp4ZDH9ziuMtuH6J0SXmr8sJ40TdXXttUc/ek00
NB/c0kTIccD8u+o6WpxNnt8c+hxcKiB9Aa5jYuJ/Yv3JfyrMppEP+Cjw5i9l5tb6
l6q8Buciz+TLvQ3jR5zjM6pqYq6hgXESNbFFc2WB1hbJz5ZoQHqfT4DO7aSBHcRN
EpDcA25S40QzKx8UX13O408RsYtassjuT5rJ1hGo2WH3FAX536Hm3kh3PFdP1rUI
rUsr9x5JjQAtcjoc548zTQRQ8+0q4qlYwcheXKepEvmMkk0IS1nbT010TdBZWsCi
ERyYRRYXwGR3QSH4HIo8oiuxllSyB/hMHkckaVmEdTWQYE/JpX74b/bTrgPMs/ob
huWFEgdYFCm13POL0hU8oZxlsWUF0dtu/ndKf4MiRkNa94BVlS0dVwQxgdsisP/5
7QfduFO7LZQ3oihDCaY8nZeakyXL7mBwvmiYxlhmUboRI5T9APgfdt5Z4CpXh/dZ
NPAYVJkORO4yNBCQ8y/nt9o2jGi++TTB19BXJIsoFyutSIx5N6PN5UUAFEArqwpF
OOPjbtgRnymXQwp3+X4/WD1O5ttLfEILg4mIHmDLpA6yXOzPmJP0oX6AhjnO3UT2
e0dlYcxN2CUDgYPoPb/p4V152wnelvDd3q7FR0GsiYCaGxdSIvs9aDMnvUABCi4y
DrO6EqAQCF1rZQ5XAzp/DFpgaMSo9oCTJzGEjHdoy+Gj5xqzhr5ar0OlF5hTk7Fe
GcIyeCe0wRcGmF2r1Vv5MBffsTXXRXdiJsBFdybNiQF30+TmEBwUAqCJVhpEua3f
ggX6kvz44wDgMJ1OwtBSHlYTFMT/4c8T2U/9F2wrEdLkmfJ/DSguU0DNCH6qfo16
KzMqLP4wMm4KCbR2fk7E0PLW0gzSLGY7VFwJ0bz+MzZeznXGJvIJbnlrHTZdTWik
hqLwY37WV9K/3YYUOXT38CacZwo//oG5oGHpPDVa0o+QbY6cyWLTbgOql5NiK8tY
Ow28d/mMPyYn9KfCcu6DyYP/FI7TwcdeVZ1gkxJeQxVq7Ng50dDFQaeBIZSBYhx4
DvHfxO52r7nl9tdHUia1a7fbEyQcBzU/jaLnZTaM7nTwvaBzmlBH+zvf6xdtm1re
ENpcffShDJSvUYWuPRs71jO8gHy85cPo4Qppk2O+meJHRUs6hW74CxJ0Fqyp0PQl
QxMQQjBiE1KN0BXO0wid2epaMQC4+HmTjCtAIJ3mkZ86iilmh0JOlm1zxnywz5KF
SCBe7NDkZjQI34a3J9HeYWgmURw1mggUTQsIizDDE+S/nDqQ2vZE316oXTSS2W/b
ZqzPT4v1EwM5+kBNn5MoUy37zBuO4YFk5QNvuCbNvuQWxyZekgONZN0uZuNXQalv
`protect END_PROTECTED
