`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gacW2keuxXDwZpeJVBB7xat8lbzM5mjS5pwYv25QJjqjQJaTXSShojAKMyTFy47S
0B/bCd3NT8AfI6ggJ7sn6GZvIV8SnDYoI9D6hrFHx4QocTigON53nK+zttcqK4IT
3uTyzqj4k9yhVeC7cn5zDoVLVMjbO6c6S482iOkzvxQf+shnNuiWMOfGLhLI/PCs
N3mH1Ui3D2dBxqf8If13t9doKyFGD1iKJ+eQkI4FlMVRGJyk0qKXOmIaI9S2QO6X
+Q+g6+rOF2Jhffs4+MGPHLelJBLnHKXvd9sRHq6tJQEzGewu6AH7WGTZfHYRS+Vt
05xwV54V6iXCKsJhVYtrmqJ3A3dFlTinrvwRew0bF3im5e6Jd2fDJlbpWx5r9Yll
PevZ4kXogsKZiaoJTjjlxsFiSsTrugWeLDc62ii+nfSKWiKWVSpNgc4sOW5yZM7v
92x8mAOmJtPXOYw17NN/yJWQlQF0+5kr8e5YxzC3ukr7KiWU1VYlDEqWdKp6Ty5S
954/yuHbUDYCJEKBS6bPxAXCb/FhnODBPgtnrl4CzmW3nposG4uW/aqkdkFgd3t1
NlIZoleRcF5j0Nu9x0kxwpP0jB1PAknmDDbIYvUe22hPQUmvVFO1LoBoTZuIf4O8
1qZolmli4J2QZ6s6JeCKSJW8ewLbcrMHtK9FRcz3d3ZqRTxYtACe/P2p/sq5tRVK
6eehqx8obnljlgVPIXcxGEM3aTDzw9dq0dZM9A8+Ov3MFBlPjjJYlPpFD4is/Vto
hi8S73gVPi3rkXZSY3Kbq+MzhLcUbx/Lu1kWGTWEXbizzcqYQPaRTCf2cREfGT0W
b0Men/lV5jjtdYOKOTLJt9yTH1+kzQ4ZVWa2FsF6maFD6HGkbw3ktkFHRHNNnen+
9ao6EL30+KXD7RfD5Qqli9hUQyw9CxQQFi/cqNUHDsFBivaC3EZ1CtHDYX5LuY7Z
zKcSJKQnQEMXWTpDO/H0ZeFyyZCjigfQjzhoFgo7EftagFOilt7v/ODCPTBuA0ua
QVRsORUCDPjuX/T3uxUNGcEdZFoL7n1Nt724xz32K57euwGf2LbVd3x1+aFNsQ4U
M6BcOAaw/XTJDhhCrtYK5SNr+EVQl7hKlqqc6oEDuJzzsxOIz+E89jhQMlJ308aD
z6h/lUIouP+c3ozuRGpYgHaJtHWievNPZtAPk3ssRPeuEYvFV8tqVTGMAwaTdLLI
LvVcRp+7tC4Epb8flPGEwQYQrkaa4B+6Oa8FyVDchvs6gMU7z3RxxBbAAygcTWVH
YPIgJBBc2V3NKlw6+ZnrH9gE6lfB4B1qUW+dW/bB87S2eFmBCA0gud7gGX96TzM+
cXJ8L0U2adjWSrTSZpl7NkfaPo5QaaNMEkEVk2fJ66W+Ck1x04Syi5qugRG63+fk
0WE9gIP0lWvspqbJIgzyUEIuyUlsLvKOeLr6DMHrnsCQvSHvlaATtQjQQ96WKX2i
BCPzlJ9HGQ4ToVssfd5SlWvIu7PqJ6rvzGRsLHRCroMTiH9gyYhhQMnGmWjg8PO1
J5KeDXOJBPG64gSMxfQPcUWziXvrZWlaG1xp6C/Ytkn7hG3ut9Xs6Kg/iRgwS3X7
k0gv572wD4cyVpbDeIC0tpYB29JxYF1v8HxZ+0ezKai6FgAx9Vo2HZBBH2kHkwAS
Md8Y1M95dKlYncQU5Wo7+RmEVaXp/xOoarEqvyj2+LS1mdOPNhXr2RpEFwXqfsP8
EHQHs209uIS/sSRgRWqxDQ==
`protect END_PROTECTED
