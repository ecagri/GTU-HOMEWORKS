`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8MLd+XI29+YAraRughA0LglzD4eiSnv00XoJ0hHcgWez4xuNvTDYA9jmopOYPnFO
W40yTDaFAmoiKhcu+cRkzGys3y3MgCVL/rToqqpfCoKwTD2f4S/hv+IzPkJQRggn
xDUV/06YsHcr4U9EuWOAPbXUvI9WsxYSLqyc37w+KoUmRlU2q0KnT1LWsn/5CV5w
MUTLRCz+ii8mhxmKu4I4Wi7sLpTppLOpcivtJsbIlQtZbTia6UCMAiy0lhWa7Z6g
yk3ENMIkR4HdpChRj4Qr0CG6B2WVCq55N/69OprjpS4Sm7F8k9QOJtHq8plJmf5P
H9gzGKIWezPTknaOKf7YwTnwdzyON4MQhOAIkwnpdvdBUMo9CX1Am31lBUnbvFpB
MUUcChIyv3aTx4MaD8MbkTPybfAtTpq0rO4SD7aufA5TyaXxmMcb2fxp/qGmBY93
tvSBjcR8iSdu2VLrvKH7E2O5LxyDSGk7L5ShrgtLhpIpf6HlHjABJvfq3B1yD8GO
5Y0ain80I20NPwRLe/Jg7lUB1fJTVBiqSHF2CRcDHN1wuMtoY9AO8uuCe2dUfwRl
k64OdxW3tLJ/VLn8GcXdkTuyw10BqTlQBEga3/kxYZ3eLFKUkdelPtjetAHljZIu
aPNdjXe7vig6ftcOss86U7MgZ1xcDMzBV6aJEWZRq2YwpK1hUXNbxvs9sFJoTE1V
MZYkNQ37XQUlAoay832ev/xeMNQ8MdtlOKptFfZDI7Am2ZB4VwTZP8584Qe9s7UX
3Jn3kWOm/UxI3OhKGTYZ31x+3m9Dt8O4U458e0j2gAK8wwOIWCJ01fe9G5E5ph1/
xDQ1obapkLERf2tMpUDPpMJ6FAm2CMW925DCAteRbNWQFd0KLQFuCr9NqK0FM1NK
15jybjpkGXwunXEupAVkSziDKnYNNvjueZc+iOzj/lSw0T2OQcn/Mg7lb4z3Q1D3
QFmAc1JgWOHlmM28Vp8Qlc7w4i3Ue/ME4RYvnkp/m2/a2iwley3XKIwIDjLNrVnT
Se5HhfqhIuTONvIqPxZLl5oQjsqqZCps/ymZhhgPOk57Am9N4oO9rWd+UO6OD25M
99lXqT7lXa34Di1yzk2L4jC7Jmn5/vKCcMqhuC6Z8a1Y2AwUZBFLJAG+XcwauApH
UdhRqtC93xy08BzLn/AnXQ==
`protect END_PROTECTED
