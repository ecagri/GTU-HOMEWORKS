`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6d1/1bD41bqbZtx/iuqRfB8HXudutVGTsIQugZObk6IS+MdlXvWevQbZeULj3P5g
1AoPIn3rVK6o/1aV7mubkS/wu/eTx+LsA/XHaldzd2Vcmh+jMNuC4h6Plvx4frEK
/SejqMtZXiqKoiKPgmYrbjCj9N25xISdKc15oASRJ5+r2ro/5reH8SC15BH4vZLD
3XMlRUAJ1OfxyLDq1StlkHhoB7U4cs0K2uT9N5BrKH3c/uFWyRJaRsPrIobf9SBu
j/20tADSrKsVcADWvRmtB5s/TDNMIY9aoAqnifes9KRaCaevo4ZWHBk/kTNiWKRW
aiV9/KWCc/jXGX8rbc+NSdQ6foJP9ib9fxq17lOLoKUXJCK0biSNBi8WmTbriq91
m+GC9wogf2+sr42wqyyK8exqR86Byo+N+SxKB+XM6+4Pc5f0mY5h4zVuQ2fOlRrO
YJTWzK1lGSSMWAkDKwKnLaWMKz2V0K5K0O1zfGbGGjnteyq0kTbAhb0bkvYyxFei
lE5ylv0jOD58KSWRzI1wYImKFa6DrmWwKJ8/HZplo9qclMRK2y+7jbWPKTcmj0Dt
yOLL74FBoJuRLTe6VrNAn9DcDWyR6W/G/BCKrj+esrxQuUI8TDlhG+L+fewjcpeZ
mNiF3YCOuSiSIpldG2b1coDJ8fX1vHy8LH/RIi7VS19moGLzSN2euvFssNj4avFB
LqBS2BTsOc6lxCWSxAlyxBiXRh8lIEc2Z/cFfpYDKpFYsVVxfdjPjZ56Tkcxhqc1
yNXdiQ+7Es3PWAGearGZp7GH2jYhcawYSxtPXeNHUSbxXEi1jBToFOR+b2XgxfVt
gdF6tHW2H1VM50770ObH9ennLCGFTEbuMF1ztCn5mMRHSbEsEwXVj1uNYkGYV3Rx
8MV2oQctI+IuRRKEIKDZrOJowzPs15EXBk7FFMIfXZf2C/Py/wWBr+CUO4yCKB/L
bF2E52+efi/eif3yLULcRZ+G1HYGgALrS1ohiZHetVMFK6sTNfhwJuvZVxx98KoE
P3QFsyTyu7ExW7PMWIvaLp4ml0JgpqLb1p+rx2JzZn8R/PsmKkLHIlKtSP0UqMdc
HaxvY9FbvAeo5SikOQ8egGNglTQL2+x/b+ZmJTAVqekEqEBjcTimqy8po6rfQpyw
wFFhLMHSNuLgPo4WnfbkhxZerESBbp2ejX+2ifqwEksJMvfO0gXdwHHWEbCRMcBm
V5m0j150tGYy/YO7mDev3O+bHEQpmYq5FQ4qVCvIOgkLgPxmAJe2gJjS4/69ecPg
OijOAjzhsx7QczZIiZ5TeVG88SZgS10JqGaJAHL3swuruw49oMgFh29rpzQWeahO
3cLMdxKlQkZ2fJVOOFsrpqVb4uqDJF1Fk/tu1qXOUNalAmbGWv58T/4cm61ReCml
NDJw56ccp7VkDE2LH18nbtmeZ0w3fCXNn/T7HQcgO2LULRBv3m9fUz0dzfgeGdlQ
ath9+RNY1Sdvv6l0lk9SZoxpEDTcEyDPNxC1PbErHMxc4VU/RUbsj0nLtwHW/Oa+
IGLGv+Vo2a6WzmZdDr+/Yimax0feI31BUUP3U9yK8dDZFuQg25GIsrIvXRBWiRuz
CdLx3ijRXUaUQT8HdpauOQ==
`protect END_PROTECTED
