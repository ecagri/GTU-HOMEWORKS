`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mTF7teblKLgBxKJ0JAmnABiKdaDF565T1k6Rj8KWQPslo9bvjJBvkgSw3uB6oWSx
OOwPwGtA+LTwM//nKz80k6Aw4eMfkM6iZv0JVqrBafH/DIryaLmv8HKBZzvd4uaY
ZkeJVyHlCGHXDAPth9IuVYdvIrmdlh4PzNiD1lCopjInjNLypxpmCEETm4i2NnbI
aWDgim1erzfxnUrXlNNyVMgZqoTDFWQktVXVy2ByCkWLDB3fpZQPFnyfVzTNEBeT
JpYOMZ93v6niDA9SqHxVWvlX768jxpY2GpvksP9Jojkh4cDPrr9hObb48XOZhRAF
ADFAH/l8LKRLsf+58XUd9Km+djhSB8/Ik8e+7l7dfP6PyBqo115Hy78DLFLiQzKu
4/v7qD5mvhOB+bqp2weXAsEzy8olOgSPdKBzdA386TxhTo77SPGf/6UpgyPi3LFJ
dgABVTGBn+BTQetVZvtm+ZOJ6ATJvyzXs0CbDysPQFfmjnHUNpMn8Ym+Q7vNhanw
`protect END_PROTECTED
