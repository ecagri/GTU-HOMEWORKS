`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MhhKj9bRZNIPxvmcW4q26wjQIh3yygQ0jhMI6hIrLQ5SAcccEQtZsrs+GnT2rhPJ
vokzg09GC/MNUJ5Ug/rUqopTb7ueeUmA5NRyOY2SGBIxStUp7CMDxbQOZFtIxom+
DOsvQJwQg6nvq87SA4spYxI0A5+r3rshNlSvm8FlsxvTT1iQgK86uZaEfZJp/A/2
CGIVueGKOaMtZQLZn7OECsKOfKgHRWYWOTAqCp2qn3dD70pOPo6C8ZB807/hlRUy
VtNdzhWbaEJL2nMckZTF2njaxBUBRAa8bxTER2GlPw7SedsA08pNswmf3clPtd1d
ldaKwU1gUlvYC5eaAx18jqZLgy4iA9cn7Le9wQL+Gq+wQKGk9JPhjagE5Tm95d4i
iZGYb95/JYVQgEqyJ5IXw8QyajctZml0UIhNH4mXrahT4ErtppZ0nicmtPwOg5xB
wmyZgPv6eXo+wQrf2sYYMaIXhVH8KgxAvxNBrmQqwMWyI+ld+VI6NbD/KWmP02fO
pV8tE1vBonDJ/lUl9k5c1hal3dPvKjV+K0ZQWZiFfoXchJLT3QiENV/GSHqSOa6+
Io9B1ooKmZKJBNAhXIklO/PFiZVSr5hxrJBppqwr9xu+s6KsMIzDY/gh5c79W6eX
V1eNP0svB7LfjmW9NUBZtze1CU2Cqog37GZPfT68Gl5j9yXrIHZNeIVM4RaY5XkW
Zk4I/FIJazorCTNGkzixU9YVShDxp8YafT4fks7xYO2JHY1uGBzb8kf1FmM/yfaO
gnzPIV4CA2ijn7+qTP9G6lKalSMvPI3GnJVKDbi/cSxyeY81xXingG/8wJQC0OvC
DpfkIuQG7XiFFT162bZHrF2JaBKHePA+lWxggDH/Y6i1u5heeb6R7mc7Y9wXZhUr
peDc5/KZlr3xaxYzTroALAP+Ls5aZA2ezYjjAvrcV0G9q5PRBnybvN8vBGcu4EZS
`protect END_PROTECTED
