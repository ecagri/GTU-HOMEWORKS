`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0Vd6VIN5sJ6ZLGAOtOonNyAXv9ZtM02n7u//avngRUTDEBWOiK9WEOPdd2OUGqmV
D/OEUM8BkfqjhHCy/EJ3GEXjgId6+OPbKfdvYWr9hCRyVFbPdt5C6OLoLWN2Zm+9
tgd4n7UOrMlUN8xA2bNKcGcPMgmoqpUp4U7g4hY+uRZ61UIssI/5YaLQzQXFs1K/
UmJQSNAx7Y16/kOcTjYF1LtSk5eI7kti3hq5TFY57D8GmjY8GcZJ5eAj2ZCuoSoo
EH85jkm9FpbtD6UNYnadzsA9CuCm9cT4fwO63RIAp5tCQb5oyI/h99N/T5Yu9P5I
4xfe31ODMDPbtiKWsB18lLAcH+oZBFyBmODyBo+11ZBN+To+zlQCgNqOAoXDK+IJ
+MIU7x0FJv1DDehc7dHAUjfxuGtmcXTLS744YA1rauBIpSc3WkXlg2XFK1rxKgWx
ZfG+PN54F1Q0qpuCgqnF/OHnvu8D6a8RsId12qE8O5jeYnC28+baCSxtwUijQPgN
LD+cYpeKgl1jOtwYQX480yHcvopLgNXQmLCme/nW7AQR748EUMgYKIq7Fg/mTOPF
1YYLiQO3aip+n8tkgFtQQKJjHUnavYVqEMM3G139ngRzCkKj/bZmaAAdFURs4OSd
CFs7FY9JO1cM/OL90cJzlVBbQorxa6eUToh9M8xyM8hbSRFKY/6xAWFe+X1HkjNm
6C7VInmTllnqtJm8Rt1A0ZnRmlX3jFJJnO1/2s6Mt9B+6aQjkVoY58FmY7LUDsow
H+CEtNsNiryr2hpkN+g2Yg/ye4qOslB3eW/U/s3CawJzjbYf+ZK8RoFRgFNXPz+p
jd33ZYfPrbSiJeANH+dDs6Fn1UEZjsyKsCzEONSqMBiPm1yhYXDkg5yDWCKB3hFH
FYzs3EdZoU5xqXQDsK3wSNN+5zlYKgFKan12ffQhxx7J7eRCtB56iZMZna+KdbJX
VyB41QIjR2BmBzIUbQCjWRItmxVKKQ7qk3CaodZJmID73Y91qjEpqx3Z65ROWiU9
+BCtcKjSlat+xzkurz1e1w==
`protect END_PROTECTED
