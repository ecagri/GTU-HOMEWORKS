`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wOT8DBRve5PJ0kH45BnxCPmIZGl4egGfdT6HPgxsHmlet+0FlSoi08I80RO75hHO
uGQ0OIZ4EwkUSJGTpLnAexEhdvvFYt6USExCJgepUL7Q8RpznYR6CK4I1X9fs1i+
BonHpqkuTXpWCR0+iZ1X8PcVROgGslE9LDa5uA0T7bykC/VvvpK7Nz2yYY9hN/fF
No8VxGKflwV9esRGAIKFEWC1gSRPFTK2Obx/zGLnsCtl4gidKwJhtmjFeqPVbwbk
vu7+5coUeJ09/6VgfO4tBbLMVm2+IAKiMIsq9m1pV6/u8qV3qSCupOHw1Yt/Y7n7
uVVtCW5p7fIvvL0hMlNoE7M08Ncdz2rJKq9VKX0Q1pMJhhf1dOvOLoK54z3nkR8I
BEF+UNKVTvKqcfQorJtqqvZ6zpHfhOVkqngS0l40aGh00EggFcGkRVpyd+xo3wVH
jVepz0WCReCPKyY1mTdShDjqB7q6OGGJFVpmOlm9+A0L1359WTX9qpLRAw+fp7M7
tPI5mGQkfsabltGUOny/rAOaQ6Gk6bf9hv4WWFYU+ZXX0u/xy8k9h1BvrvoU8HOC
r7ZFGxp6tqgUqBdQLpoeGVQs3M4jmSCafHctIIbd3grHQA7oNrzur+B8nKWZZ/w9
Ruae7LleWxowb6Ii16JNvEyq4CRviZIYQ57HhDgRuvXxMC1hiKCpRkOVLgUlCxW9
tPYgP/qRtQtmXUilHYBRA+9eP9RSgUDJ7pzYi9jN2JNDmZsYaA3aREK4v54gDCQo
FTTFBmM6Rj5+ME8wXE+4fbWMTge+h0Gb60ppzfWGmZKfTLlgw44DcVC6x9aZ4k5b
t3KlY1CW9JJW+j66qJ+cL4bxMId0rQvTClPpyYGh7s5Yjq7Hoj3Wdpapy+j68PXQ
V5dGV7L2zFWjOMAoZcEq6Yhooy2BW6wtf4e1NLlGSmU08rJFRnu2x+hnp3XLqe7Q
UU4iGSvAFCTV6BbpzUa8R3TqgA8CFqmASan1Y6dxnJFEDyES4sI1WK8L7rQPvyEU
Hc6d8OiZL1rD6gLCocpGlRhfqd5zA+IOHRw3JTSM+uCmEVzk6qaJMXLbmSpuJRrJ
YIrDD2BDaVl8FUtmHmd9xK5DA+WdZT3iNKpM0siGnOP2orVFk4X+vFKU/xcw17if
phc6VoMzrUjX9s897INZDh6CYNShm5qezixWoOqc10a+VI0LdsY452Ue29uO55+h
o0txS/wWspnpiqzwgHrp7XvypFO9u0PCtZAtHwt5XkKerppqrWuGlGjsil/IVJsY
n1LE/UG2k78hU298y/5AfZNSXXsQkBWwWszf/pBJQ13Im3IY6M6sChIOixaUjBOE
J3pCvQ0QiKV15JiiQ1G8UPeW+P3GSawLUGnMBR5oHPYXaIuxs1+W9/ohhxDS/6Er
ZGOZwMd3sE5x1tpwBA5rGX2vcfltO7GhYJqIghp1ySGeFdV64e5bYYLcUkUziNol
3vZJOGjgHqfOHgJnlOOg4S9dl/XzrH9bOkHncx3XgTe1zEd71fLbWX25xIcK2ukY
DxG61yCXzZSuVloL+07utmidyQCri25Yv7fwda+JyM1WVBUA5ExMQsmCeUfISWzi
yAwCYIvswEzkKIA4fWw2PLE4PbbM+tvG+y/BA2PUVjMKzouZWCBCQB0kYsoD0RM0
kvcuNHtqftF9sNcJoiR5/7nlYkVbRjlST7uDkdBaiwrWVzRm1xDMlCHVXp19ePCb
9xBRTllobAdAC6bXMLsfMrI022qqWy+083KBxT5JPHJwa9v6g1HRopJHByUP6D/R
JD4kST42kRAammRGXhYQ5/CsK1/TSXgDG0x69LXxkuMxrMos85BtOop6sm8fdG4o
76qg4OvgWgt6KcLIvnvMC/qtVvt8GzuUvQO5HpUENteQ4DV1er0oIo0U4intsOpr
+0PyiikepeENsFIE+mz3yI959b20O8Izhy8/BRXH7ezOUV0L9KvAkwygJirK3kxA
yddu9NG2P6ZS1QbDBGE5jSGgpHxsldpP+vnQSogcOEBRsYMpLHcYFBfTmy2UcYzE
a1scDKclnOe/1zPDSALxbZrDp0i/yxy6XgN2qGb8FksZooauVHatdouRqkhwbcsr
T69YLLNQ7HBM4gP2cJMjA8ylE2JuAZK8Rs84ZzO9i+B/xB/3aht4FWNExzc8j7IS
7j/EL59CCjH6l8gEzsDRMtv6GgfNqGYtAHhwd9tccjlrbpcvZmRrD6Gg/FwUHpez
HpAFXd6VmlfzcJ5zPkPGIiCmnVhYuAspPcsFt83TAEWQeF4dPESSUsIjlrURftk/
DZ97mL32wZd+9fE3Ey1DyY6tpWdQRHES3XEYTtT8siVfJlaUNM4GGbMAD5v6DJH3
xYxeaG5C8I6xwtG57x0cZzBb4wZ4zoofWKJ5+tgzYymi2hKUQXCslSPAUy7DGP1H
qhq237y6w3cHrTUy1d2FB8jPcjdHeMZC/f75E1GMQ2GYTtLelnFfZN0T/UaHvjf1
BBymoOGIacyEYFK3bIA9lXRNBJIjGfhNbIsG5YkNL5vk8tQvPdOdfXVLEuIlKtZj
3xRBAsRaMBu70o4RdyTHXzi9MQ+N/VPeG67Z5eFBDGa3rZhenFw2DQJzkpLqysNi
K2co3oVPBcZcPOO652I21WXi13PV1qLh9Xdt+tVLNj/Nr5xAn6/gwDPZ8JAJGd4v
YikxdhtN9j+JzbDiedipokyytXtk/NDJHd+259AI5zhajOdYCxrFFt6bvrbb9T11
/J1cRBFWcVGo/ynn1o78hQt4HBKRTVzZMSbOjzzDSNdcuUOgVt3lpQ3dwzmjUNiC
PfMsCc8wMiEwn9ngpS6NLmp1D16nJOeMg1G82kYUZ1DC+UiJ6lZfvOAatWEVgc3/
ghUhF6+ZksZ7yGMR4eEX64lDm5Aa95kammkibX9ct4phl0iZ5WdITBkfWauDQMzn
cMSrCwNt820Ozl+bXU+zXTSXNWE87oN9VXpEiOh9zeqImUnbqV76VM8YOkib7BA8
HbeJmWRkCU39Jg+SPQs11Ug9ndHVPI8n5MVgKY7bgkOQo/4lrZsxO8TwJGsJHfkI
qdKcvkpM+AUx/nPyvCRnzh1GRhLcl0g7xuwodsRdoo2ZUWoiRCH0EiQ6CT3jRHXo
et0/aGc6OQh2hUnjfO3hLRQSRWDIcx6dqfQ0oblZQX18uHBcI+ryTsswZOhoUuzi
YmaDDCZp4q2Y35rz38qV87XpXZtkmxDvHfCuo6oIGmw4yeAsJdS0cmYyvYD47BVh
cOhEdH2vc9OOIFWxf8Ft4ToVHcSHB+YjxrKMaMv6EDz78kgWksdCY5mjGdooYIL/
ZU0mxBr6n7n2BfKhMXk/9x1V/w7IrvAOHObYO1cws4FJAI9yciXoksl8qL4iVft/
Mos85ep/daHu9JdgF0/oIITpJc/Um6cTSewK5/ridZAj06NGaPg8FDY7ikE1ELC2
z0CNhW0NqkRbGLNhArDWRGJ+cPt3Kt54M4NDRo73hBMO6xvOLIqQjFdnaTGvMGzW
nl+8vdekrxw2Q8DZoM8Lr2Lxk8CpLsRMnmquLZnB3sXH9dMnTfbResKqodUaTuce
XpWsWOWS/S2Hn1zUI7NlyjxF7MqvKlp48radSrVDRYRMsklLBpJBdRxbxQ3buJJM
4NwUBgaxkuBNBD04PeFz/cx4BrWrSN21EsdkJUbQ0xKb5eeq3nvWIhWD/gRUG2s9
YvkwxQtnWZGQvuImuom9a/pqmH79U7QMjH6nfrI+jdC5p/dUfFIE6iKF4gy6UB5m
x8O7ORzAPs9blrXpaJnLcepmrmx4i9k8jaKyR0e78oNKAxj+d5o9DLg2eLTXJ2wz
dj8L/aLyxvVcgRgwvW53vn6oVSNQva90JJjeb1qWMltjg1vo1nKyh7/gbPRfMrmM
U/3hZShHJ3UCAU5qj952eSQo8f7U5o/Ve3sFdVDY/8d2UubjqzuZNgrbhjpYn/zF
anKGqt/zsB1v0cJ3X9etKgfUJpmg5wmeAZEPqFWpQD2FZlR0kFly99E3aDgNqjUx
D+R3trkhbTvEnOo89i0XGpSippGbpW6SzE+lD52fRsbzxEGIaaDXFtzpz0s5kFMC
DNj0qPBX8MalNgtKuV5l4E71CvutQod5bnnbzJNTZzKZewmUh5dllNnG5vuNj5pk
VCXbnV5Rn9ygSeGqnnLLKoNdzU0BPxb8V8LGqv4o4mvmSBTHe1Qpb/lAhSphVE5i
PRKMRbs7vmS8A0HDdhK0y8abXnOrNjcxj8lSG2UOLyg2sWimvso46x5mBK8+UmNH
21hgQhEz6UpNm/7tdSBFvbpyL2Oo53kxo6dLfdtI5tXeHtgDafeMLI7kwn1t0/iz
R2Uw9kKbUx4KFy/Ggbla8YVVQDvk2nKxpAoWL6UD/JujI3z0nhpqG08MHUUCwDM3
/ncxszyNLXMB3xEbE1lbcJcCM5eCOYJOvumJeMXC/6RCjuNBOkGcW6gOhgBwhGh6
4Gvkj97E6lYDepMwFwYfGyG9VrpCBmc6HiSRyuUf4i2tBTpbo53yc1AwVt4Bxd4b
IRhthQLaK7bIYWZ1h7lmJ5kyu7YCBxLZSpMXeqMf7IdHjbmnTvyhwKIT7K5bM3qh
6qgD0AqsyZZ7KlCAxy3GE3+p55QLvaOQH1whNlHx0ogYp10JFsfGseVvrgy9vU0K
5P/Ns1rpdXOARyUn3jLQm8qyPoWYckaHdVQFXcIcgYjewO0efUezY8jHoAPN8vdZ
yEDhU5PcOVGun68qjBKESzowt7Z7btpcuR01Mca5x9AoAwtsaYtGRPbLtHH2lD9e
j4iy11XUkEH9lDWDexr16F4f0r9JWa8qlTJ0NSTeu2vDCN33L/Yc/zw4Cz/HFK7k
Ake4i4yfuF0qc711IE1iW6ElEiVVyL1tu+rNe0HlzVuYXRDru24gT3d+9p7GG991
96V7P3pvSt8m+W0dgV5FIicNP7kjYMf+3MzuYwaLawcf+7r16XYuKo4/53Cnzqto
VijylRly4CmGE/Y+MSH7zsnuYi22cev/iWAP0zyLAwq/gMuqcUJt6iyuPq7vhFIA
mDjgjiQwKt+zt9VMvoGFHUbvkEff4lGEPFLBX0ZI69gaCJMs1A2BbG/BEPU4sKZ9
9TVFFnaveE8bWNRV+QfnpCGVNuOc9JKRKpzM6wU1a9sMhvCShN39Bftt59F1ITJG
9bTJ0PMiN07sskC78yizjdN8Xbghtgwuz/7rGY+yzE/DAj8IqHt2+Qp7GiQH0VWj
aYzeef1si5BfApxrQv3Fl+GT+nl4ffamKIJO4HClh30X5zye/0PZBFPT0zzVECaV
ETC6msJW9XvNU/ZGgOGBl6FOg3yZbxvI7TkMJjxtDNZiZs474MfruqbDLPnsh7Ug
Fz02yPl76H2+J5hyy9GsEmpRrod4EyM5aoADlNkwpjUnrmBN5sHH6Slt7mCTmA3Q
hkxk74imD5XMpX3WlUZNr1RlYFR7q77LB56k4harEM/dDN8+nE+xUIFr8W3RLz02
UQqm2hJtpgOuBb04Ho/8IpzWUe96RvLHgRUtqaH9lvQ1YK8NPohcyod7ApuY0Des
ri+0d4niEqTN6My9acgErwscoE3Z3uSRC6CSlHlJUy87VmQ4YaAZCvXx6BxTKR+5
DK38YPtm/QtMxg0oA6xxC4CRm4faRK+sALH1Fd5f/1L7lwcMFAB1Ql6qzWI3vxjj
cFJxgbYsZE8Rq3L8jagnrVh8wKRFbeXx8A+RPzc0qwnmouBa32PsnThpRuFslkOC
lpSWSEwJrmxx3rZotREF6Q6vjccM5a7SOm8xN0KSp/s7vC2d10CIZxOEisGswa6D
JZjxYld6mO4FXDvyXEOVXleWrH32at0oTjcE703Y4nFFWpK+Jdmp1m3voCyUNdob
tMLbl26LN2HjVQBhRoF1ZjhgjBkd0Qlu1FTabfHJpgKMiXIWx/Z6URi3lw0FAGZ3
D0NpwMabwuvpUUZXvyXASjftC+b0ghAESJi2nnilYWK+T9t0AbXuSmMnFBNHL78e
dxTKsG8MLDU08AvogvqU6eOqk+og/cHnADkELNZvpG52a+6z4jLkIS42uNYYikkg
cn5cCps3ED1cQg7qEcGJ9TLWDgdSNQOeLlk8uODTrAtQprzGY14tD6bj/ILPulXw
VI1iT994cJ+H3XhGkfkMS85N++TgIuwYEtuMZlgB4mUPSKY5E96i2e2rgi8ONpjw
TUpys2W7HkVmNKh7SzhLpOhspZlu4F2NQu+EGRw3DoRpwvIHqCLmMxvH7IPlLqar
2w3RR8/ZYLuOfcx1wsXQViN7Pc3XYviic1s3rPSNLFyujTNxerYL6ORfrqwE0m4D
StmF+8D52iJiAKyyEZhqcDAparZdO5HjyzqfKASkhQtDU9Bhi0+0zx47FEoJV5kK
SADjMc+OUGPAreGw6CZkujTqoODQDI77yWZo9+m81IE4MSIsmuKyk2WiBFKHgUcH
IK22N2aTcuSj8HVyvO0SUfUfKy8RiBkMrVobA258RuVUexQLPrLucl8+emF/Vqsx
S86fN2I1biOWsbTSh9HDsM5idZ/omJM7r0epno4BkAd5EwjtUAvyQKCbE/1WtISG
xek8eSweC6PvDpzMD8j5rSkFTCXv/UYvz8ZR1q3JxKYlVdnd8B4WfMmxQXmha31T
e+SHF0NW7k2C7ITrhAbmcB5G3j+Q0aKp2CXyOvCR1sw/oX+4qzhqlMgLvvYgZ211
mU4O+5hri8IFGRmGZen+0tO+m+CR7HzMO5/qFBvqqyTJtQOriST1VXtby+xbd+/z
zL553cq6CQcdb/eCPvRKEoKfyueq39AxweZMpIjcu+k0cWZeI+VWLUU/0t1pY7Uk
naQxjs4dzxIAETxewX10bsWivSByyfHRHkpWZSSqSZ4=
`protect END_PROTECTED
