`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VbuLWuOD8SRQgP02dXrZsSupIYLgwv7zocu1r9YcWPizAaj7rSgFmU4QKOv0/b3s
vsEtJ6CiZKr27Efx5L5Lb5ZOvHDRHpjer7ygDnVCjIm81IwTn8ZG4KoQi8gjzUJv
PCDvZopHMIyLkcY7lyMUTloH4DVGiLd0HETJiqjctiD3nlgZqONbUIeLmjrIjuPa
EE5ZfWj4feEaP+pmIxfmOwV+qejBZOTBDaNfx6epMd5ZjthTTpVUx7gueyGNKpu9
iwFxWi9HhNRgPT2Sl6oQpK2JGjgO0OrihZU+V24AEyNf3KA00/s2MdLN7AY9MVQM
k0vhNcmg0CWVQrmcXrGxeL5qR73K/N4IaMTJVR9x3jpwhS47+OCD4qTpPOBJaqrB
EZmEG1FETSS3czDj2hGGzHkcLU7pH40D4lREOr5n4G0uATG9NS1Cc5BpZMLQu8Gl
Bmg+NiaTi4h4YOEVe5I5srNJrU7imPQ31tJ/5OzsebfDTfwjzkuHa5FKc9yWCAtD
sW5r795JcJ2dSRkKQHZ9gTmIBfHOpyytpRYquZ7INed6EWAfb42pQN+3Y8WOb3WX
YrlvDbZNP9mF5ouMYOkgVpSX8hEaNbEiHsIS+SeTRgIUu2Jdq2smVlJRan/MaeoK
uNWfTB8Oy6lVScc7ubPIZbgkEBhnD712fmUyoN1C/QM/PBGnmOjCxV/q+F1q0hLs
0TY9cQAjCq66gqCw39t/ITfnTQpt78ZOKoq2uOzt1Jmi3QZEV3XVTKr05SEetVKf
519IWWwjyWrmUMs2MCKX1k3F5uyJplXp4to56oQxblLZ/QvEzP8XaXDznVQDnMJD
HIR6pniJUEt7SgFdJADegXQkCwiGKIzd00BjkeK3KLknGtBF/RYEnhdke7a4/rYp
a+SCzklEiatDGvZVOIoAMscKqZcnChYl5sAieviJ5gEjvbtDFJqsa60FVXrsoL6I
pCbT+mMkWnD54LY5CBFY0kWnxsjFoAypzl6JaT3XKbb0JlgTO7D4zWW84EWTcdKl
ZDsZZT9yE91H/xCM/WcFICvpj6I6dUtoUv4ifFfBVdkXmZ8xBUo2P8EotUPyDdqj
rAonUs1lHaTUT0qoZ1ofFn9axRED8wfc+oIXGZeUXLIU4FzezD24GR/K+3JVt8g/
blxOGrcCgqS4xHBULaRrrlfzRbuP0WEgRuPN13Y6A8bgHIZ5a6vJVw3zw0JsQ40l
oiNdzDfO6S3rm4S8F8X2VIYpj+LdaZGLpvwEQRF7porj6xk0o6/eb18Ikjro/K8i
4d7HcCQrROC/8YBV73DoywY1Sg/MMimpv5KtbefWW6Kv5sDBVfz/q8gfMifYHbvJ
ZszW2UopKJG3t86irY7kfHRcfoxCTtr+HMoltyvQqJr7dWYfz/iqqSljEZSfTF4w
1mjLKu9B59iQGSscIU1TDv6l6wwOZLs0Ax9ejfr5CCckzSGXuQ5mA/UdF2NyoI7h
y4qkpC9TE3aEaZ5ad+1ETxKSswnmWabyNWtG09aAkQVRofGmJsB3Qd3VnHp4QbrX
yJYmC5eFQjXH9/iZeFQjQ4hD1yEfolHfOrFPvzFqPq2q+Rs5zEL2Qx4wvs1A2tkZ
2Pn0Iv+z+17SVSAvVBsIVOXipVB9dKKKzO3a3Pa7Whg7rAhdfbInrg8+aqMwjlcf
TRAYfowd0CClAfCZkW36gtVRf2O7FnqfwVKhYaeuqqYB/o47CHYiacX3qnVSsgOq
0jlyxVt2Tq+WCUCKmAiV0YhwM97jqK7kh2i9KVx+v3KSiOTAXZGSNWo9H9frkTM9
76XCZlwwSss0ei1uNa/NzDRL+eSwFA5qWIWTd6jbI1hdG/eZsmZzS7lfOUTPFWLd
WHdeyAK/LP+nuJHOe3cH2nHgrDr4lQHAs4n5KoNQ7z+GZaQTddKUEsRdmn7sNIas
7YwO83gLjklu3THd7ABzKvCO2aDP9jOIsngg3+AB02UdwKUJdPZFo0E71IrV76Bs
wXli5dCx1UkuTx95Wt4qxrWSLz+Eyq80dZ6VY6AfGhg5Zi1J+qyeQHQSdmq1AmEZ
6V76cIKHMouhGbXKU2sIHR5emOb292ePiGGdrv25GoT6FnqvUH9KRXXiuBZswG3K
g4BPd7/9XKHxKnx2JSIBvX/L6SeYUYowKo1rjq1K+6BFKOUEic/exQXgqwNbwNPU
FGyNNGiqtXO9yA/I3xiOWyhIRmPK5kPeULCc9sCRbHpQiKeVz0jfsTf1pzoZKjbI
bYV96dRgFHRtOBTX1Fk3HJ6myLq4/TKorrtHj4sAdfSoREpwSBFaHUyAwt+/5Flx
tDNAgPLkEsXC1KqrvhkmR2WbrxvjryNDOfLAx7PuKmsl5lT/WUL4eWYpxRfiLLAU
45cWvQL4aOHHPE8R6wMbqWq0Tfe98dMtrPuJlo0kxKeiX/+2Zrz9KTk+lIHZem7D
gAEZfyHeX1yWGPNYPHgqF9ixJ89m8OhEqxQcEeiGK6Fqj0nrBKo3Yt9IcEW9oIs8
BxwcGJo/5tiKxghZoKoeeeWxw/pp0N4cZ8UYgqE8LUX/yO94QXjg7RwvBJsjSzRr
F4OPPy4sfJWBDEE6SiLJpMWSoo+DWNcSoKWE/029/kmvkfIi9Qk3oThGBLXXSUOs
+XaWDSLi+phszs9hhslvz6tLDxnjKUpkTRsDg+AhaCPuA2xoWXfIsonQyUURtFep
bZPmAMDXGcNvTdFXnnitc3aQ5k2MJmzcEUAgo/nAOBBZ3UdHWm762Xw8V3K45HM7
Iz5pxwa5wZCS3+NU3EOq3YJBHbJ42b9xmds2ZzKsx5/PxC/KgJUB2SuVpd0PHKQs
pnaXSV7I3SvQt7Zm2pvn+mceR71J4NQPNdmpCf1FfScIE02k1rfGlVmUpRIlPXSn
5jhgjDFqAoYcXP3bpsq4PL2xMCy7i4dxNiiV3AMMu0nrAlEIDGdTZeWuIZIB155+
w2/Klt7daHsOZDiPqsYMvbRjSjP+LsxQYVI8JAoXpkzz3Awvmv2Hgf/ngiMwRlby
1XQNk1M87xPsSUGfGt3SOb65ZdKsLzp47s8ud+uST+tWa9Y2WJuDXGclSQuf3bhb
EB2QGp/UAEj+FRcSjRpOiABGQZP+wR6IAKdJLuFYQNIyOxQmuOcfTvgqCOkXzDV/
HLBZQphWoXe53mv42FAGpf88Y5VQrd5i3e2upZFt3IxlEymmph1eKG+qtTOY8zGI
0fFNXzyZxHC6uHYBD3aWWuklLGlP11nnS4jpl7ExNpWc4PrnSaSV+dFNYQhwSRvm
yWYcK5F9QorbN9BA0Eq544FBM1JHExuK96fAnz4iGMGVcuvxv7FkW9nS9C12FtGE
1j6TRS61+/r+TzzplgAyVKGY6VTLs75JkUNoVV6tj7YhFxE5gVcl4KsiQ3ronNHn
SbK7GgnRpVClLn6ISiJN5I4OV89bdYeTEXEKsu0aAIaaCglfKauV1CwYKf2M9Evf
3W1mudTxNd2zRDKwO4D62fZmF1IR93HwPPz8B6ZfcRwnchy4Wxqba7KcYOBucinL
uiNjznc5YtljBOx7b/e5GNHPxkK2RG0AERlYIkFT03zrKSolji8YmnBF6wcm3Db6
QLCN28LSvAuDUpHNYVGx313tuSZlWKnFZia7wvNQYQXV9qWwe79hMhootMD1cCuG
Q1WsCttO3QsFRv2WE7fsQb/5LCzNvfx0TzSSyOFKRM180V6CveSRUKIkmzIDibQQ
wfu7+EE8XU/HyGbcJns9dQ==
`protect END_PROTECTED
