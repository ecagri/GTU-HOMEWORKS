`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ANJXBizhiuA7ZILFXZOuwbhtQvXfQ/GmcGYHrH/woATUktaADljdhDNRZiiJS745
/+B6xXs14Lk/EgCa54jZ/gMav7oM9SEVLTeUwj7vDgKf3B0fRLSmUfSqzxmkXybh
5/+zTKtVFobs99bu/KblXqqfhmnnAGBXokbsdYxu1cR6ptU1maKfZ5qCg5GNw/Mh
ELIGELMRtL8qd5oeX1uoVxcaRhmlOT/W1BpgGI9QTb9daBWKK4F7bM4HsRjLLd6o
0V/m6zV50BH7OVLU6nEytRQ133MQf1/9F5rYGPVx23/u6BB1zU7rmmXqMdgJ355a
jTVgt11uywt010C6Z5I7V5ZVsavVfC8Unsro969C+WEYtEO48Gw/LM5VzRi4akjJ
ezhbXSP+lRB/1qD5DmXLbNxgguWGNJQnLA5dSc/wRN+el4Ne2YZuDp625k1gpg5a
4upWgnlb3Imp3SANFWcelUZT2lQs+3wuRQkWzWg4+2Xo5+mbR6sXNQgz+DTACmEL
0ZuUnRhDxuVmdXhopp01YHtsBrlvNYQBQ5oI7rKDEq7ux0HsBt+wGYazQGtwork4
nO6PXIEeZLO5kg38xXeaduPYiEJU4BCA13/vb+FV4wp9S4kuywa24q8kkmbykeA9
6FaeUFaivrRljZ1TEc87QKpy0tbQ3IHyD2QDVZU+/Sr3f09VYSHdj9r7NT4XWtzT
UtrGTfypS3WA2z7K3FJwLlCzNavtARoG345+XUnztbPUkRmt7AlAbl4eiSrwrpwA
d5Vr8eDryZlhusTGgpjPEvsxOy/WdAfQRnVLH34Hq3kj5qAmp+hzuoSucnZXm7I5
j4Ip8d0qe8o0vy73Fn/TAYyTtkzVV80EhX/wv5PAdl8qKOYgDDqWVK39Dqdm7pk9
93zWBejL63gFQihEwzXNEYjkmhcENfavEfsLnlqnMln+lVsN+eawRBkn2a/Vx7Z9
BGsXQh/XYXFLygTtSyUPniKAr2rWJd6E48+VdC9DPQ65kZlM0DAPDfX4Zs28JibH
MLVcqJVA2IyHlU1nl3EAAuhhvyazfr+x9gFPx+t7yW6xc0DbW0XJeDIrM79R2tyF
83rx5QfjBgB9xP6ubJwiAF3FX74cBVrfRoyKWQtEmlhGKfMs+zJ0h+iMdwRt806l
vCsp9uy3aA9Zj1/m+DDmIgzruNIRoi8N/1Ry0oXe+BR0MeEjGOEPjsSA3xtzc6OS
joWWjxscWeJ2PAG/kqf6Myj01OiZF62fmiPhfWW+Lh92fPrLIyc6aiVi+WIys9KM
PaY7uR/lOYw4pbeYijv4GVc2PdvbQzHRHD/2EWe6yozWWEJ5g1fwxUcokgV4Zpm/
+AMANw+dZIIuvsdcfZ5vae3S80a/KtroenVapP2H8L0Nl8bqhgsGERQs2mBjtSFr
i48b3nY2NxdXIqMmfhB2rvHC7ha5TKrAE5UX1Bl1NGgfr2ggFNWnoVJj7AyRr84i
`protect END_PROTECTED
