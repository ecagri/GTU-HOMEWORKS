`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bYFWWK6WT2ikv3gFKNcqrjiKwwqBgZGKyP/pXk6aRalaZ/AhORLOP6DLVBUkhwuA
R/xUihVnozd/AS+D7KwW04EEQ0bLfxRBHZcqAYkuQxGV3UbOLvnRTcsMCGCoERbi
1bzXiK7TKFEpE9xiNsrTZz6yBfO7XBEiSokTUzb+huAMQwOt/1iQRdue15+BX46b
xOKNxN4apuG56fmgwPw9Euxe7xumbq1rC2QntOGNSQ6TklM2eyehQjh0I0u3nuF6
qRA00ZlN6o2BkUxV06Cs58P4V53lLNWaioz7IAG3eyC9VUNv/6n+56+CZ37x4/JA
svUldIvIWIFyqnaurq3pwB4jw/Q+9M0l7pmBuXPMN3Z6ICjX+cPTzGcjLkq3MVFr
FXvpIbYKA87IOolMWfcybXT/A2zwBuntvArGU5qh/PtzuuFPeZSi/EuemIk2jE9p
ga31Kfim+tVjvH1beIenebNkfmWi2TpiOZPrOB2nfuFYhTAYzMD0WaBoRS4bR5qa
UUw5ieMaCyefiwC6eeiZ5jRtScvIviPqCXeQtelmUhngBWRy7EgTUPscj5Yr4z1j
tm4eK7X6sq7D8PpZkaEAEeBpXhftO+Aqb2P3/QTfvByyHHKf5FjZ/go742uncm5M
m4AGOH2EZ48uleo/SieOyTxZb+z4vhGXjNWrg8EqJlv94ZamWlbBaeOdksW3Nosz
XG6WpbEHWx7MruLHgHONsk5dv+ljbfO29TG4ApmEd+6reuDrYeHUqeNwzivY4Msn
2iYkcfYPxVlvjynTsulrN+v2Q0pVNF01Tr8zt/IoWqE3LbiZpL9jXY+D0aF/3aP8
ciLZnWpSGPvmxV9Rv35c5ToKRFRGGeu8sjnNtGzQucLHWr85k+fo5P7eboNT/e+x
ObkcwSsGD9zcjWtkjiQ/Ii5PG5UZDh0LKSPzA31KWPixnqNCsx7UfnpCO5lTQT0c
2taF8aOahDFntkYRkUDc7D8Rw6vQg0lRA8c30vSjH0Y7ef5mclwCawot7Dl14ha3
VQPhsRVMHivv3aiRUF9/n2U2q4ojtPVpNHj6gxo6Z8ksIKeDgsn949n1cj/QlLay
g9xo/a9SKZWSkZpemGp3VdjvQEHhyLtlhIHC3+cSMHW98HOHKqTLiLaSO3PtyG0p
rZ4q4zBSHU6FPqWnr7S9MmLD1aalKY/dz5TbHDUq6tlxNaEM5ZOgeM3FyLC50t0G
WMI+DKPuzLZ+IkZxL5jVUFNrj8K3fq9l+KuCCHUuUnacYjngnmd5QUBl94AhzxbR
++tL+HatzfPDUvDt0KhE+aoqgQQ9qRY4SYyjjVowJmz4wD+lR+/bnXEVTT/C5LGj
WN8F/xrOGb0R570F5SyB+VetZt9QwXn8jfFClbz6jM1LJMWkp+qmn2sAo/f33oBE
BjTHW5dolm9dMJLcyIrUgpzoZEYPDh+xMYydyv0sKWM+eusrWGoD9TVfKtPmUp0x
F/ktJZ0wwYmz4CFQBsg1ZZ+0wMGAg1orxmLi4SfRS9UrJw7MkF62sDDggbIgDnLt
j3D6yR8K8Yvr9N0KgqkJgeWMt83SI6Md96L1OULXKjCpr+tubxd9Yjyr8rO6yG9Z
ui4biylBQNQIgixmiWDddKBOVU0MaNveD9B6MqwyjMycIuqhy+mTiiwRpJvArTK+
saDJWOyVP4AdFpqYskbkGupN74S02SNy83fgV969G3InXizV/SfDT7vAz+4NvzQS
LyzCH/YmMGyOucHL7Esh1G4IhwzdXEZKhDWGQ/qaO8H5sMMIGKjRk3BIQCckyOMh
OCYPVXzElZSHUdT1DYei+JMMACKQQSEDRsw3BehPzGACivxuPYxCdvH5iCOUYHrs
zTMRJI2D52otBHa/6P5n8AZIRZn8Iv+SvUcDOBeh4xdSEunn9DwtO59kEATKynva
9yWhHNy+oVYK95XY0o3JOEiGGn/NzpqbuprrGA4ESY6ywQwCOL09vXHAV9+cnKL0
X7nVBBVmjHWPqFHiLCI9fw3MmTg5p8Qc2pBJ+TB3aXvtZxB9LC6fTMjFBD8hVR8n
P4XAp+PC/zJ1gXYZeMiwABH5x3OKbWlImCLwV+mvmv3V7ycd1MsaGtqGQgJfu/Gj
`protect END_PROTECTED
