`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sUrVOhV8fTinDpiH2VwbKq1eXIKJII8AkrIR5YetRgRthApeGdn0XOD8CL7vZ7Ns
vvR5ugAQaMq/jjpO/ffbA2acu30CZSST3pUf9JW+HhpHg1r+6rVY7Cfqo/6hJhqk
7JYflgJBWb8N0/K8mMdq8xr2IRXlm93l6tWzPWzOyD0S9Db59iuEmxxi6lJvLDw/
wy5DSva1ALkvI1EYF+lXxkUNnZt0fcepIvjmuD5/u1zRt2a5wfrardZwSUPysYsy
6CWeyKaVZRFiFlG/IX/bNragnp7Rk7CIVCb9Eaj97V9ULyBFOGHG+kOvwuAqAUm/
RaGw3Mcm+s4RImfsj/xp2gBU5yZe2rwTWujZxx9YDapd6c21uoKDOfGn23n/j7Bz
nu4E1GSFHgPT1rL57o6i1yb2wAg10W99C2x7E5bnIbLM7zUlUnAkGZ2guc5kt1Tt
vdO1JSkLIH7jWEzROg2WP7JyLMzmsW6Zbz1GnC88oy/YOlf2WA2jS7IDywynfW5/
WAmA/BDnvamAJSD5zQB0zzhOb0RUN4Kt+x9+blA9g9tTRn5cblLAOOFOOC4hWHO9
i1Ml3RdwEoNmQRjrXKF3WVACc9ANyBA2mazg4xeXP6cI0Fk147nrY9JLTDdkVVbg
WhVG5qyvqGxnTBIPxzvCyz++mVuTUAb3WzgU/C0Q3HVh/RJwVkFkZdknow4elsVr
jK8nUFpHWW4yVA7wK/qcBR+0HgeFShMUb8h7kv3yZ5BQNIaBJm1bQ0cE2dg56lUH
/8olYCAfoA87cbMzBY5cIyvYwgrZ/rsTplZEhcrOhj47TGKWByYW3UnX10oMEGNA
O5x6dtZXmhZhfH6vyMaUNenj074/AlXSsRi9UJFuMVUocbsCdUfvFC4tjID/5xNo
uGNbXffxPl4rpnj419VDYK3YNcxvqj9M7wF+9D+0E5ZmcttM4yrZzP00rcl0HJFI
JKpRlkN6MsZNecWxxPahrbr/wuoev28nOto4ASFaBwQWEDkrU2sORSJRko3SsQb4
u7YtQOp/onkmytg0/+Uuk6F7FH1JSCIYBYGD7L81+S/rZdpB8LdKyRO5xtMnqN2N
udk8xPrLFFPAxLcljj6qTT0c1SRgI6Tmj6JB70x09fxR7S2cdDtYdex8Ue+qFjF2
BPg4MAz5ws6aXFqyFm0vK/5Jq0C/znz1QLAww1SiZs03HCSJntFFNrU1DNs79PHu
17idBNq9ITRVSNPehrRG9Qx9vmJwu3n0LO1Za5XO9nH+dAA9Rv1UCxIsV5zm49eN
Oy2yoZFdtyVRvOrjZnyDdf+jLu77rYIQicqPviGW/4UPNbGw+xlti49h1AoCNsGR
cuwoc4JndgoUfqSPLWbFjxTzdTlPznMm7B63sHMoKoEn3OKM9VrV+imJBESSLJx7
2/6Hb30gnVeSEQGdizdKspkknO5INKk4Pv5oy4h9FeZlVziUJxuhE0oRFYKHMOUy
ek2B046Oq9NaJrQa/rul/+lHSTnx9098j4r79JRIOYVdqcHZHRBBH/3nWuFsnFxx
0h/yn/eRjcsS1FACT6qmNjZak1m1Dzk6p1LzZsfpssEC3n0nPnht9EzbTgkeRumb
d35HB+m+ahfSGKecl6FGaAs6nslYvFA7OZx+aw0GQIczAFNxws+QYWqStVeK/tLb
FFFC9rUsDN6Uk36aOrq5E0lJpHOAMo6Lxyk5UvXrXIX4hGgtD4Txu2l0RMJG+0D2
nfXyJhkKqy7gO8a3OYaIPeU7cbmSXN53+d2/hafAFOr0CW1rQcB4jL1DSBFyNEYh
kvGIUuxDKHZS9ElQbHBEJyuTkVXKJ+sUX9Bwhz8DM8MSFsWXAeAVOj9HIYU/37OT
rUwNrg2GPy/cfy2d+CvCvmRA/bQHCI63uaeXrK0CcvL4XpjmYOKwt9Ex6IGM9wlX
cKSmsZk0r4NgqNAJW/OUDzcMhAwnnpzHlO11tVoleuChhAlvPteD5bGSMSNgUDdy
fcowbMMD4630v+Gkb6IdkoQQSzb42AFs0P0SxjkJYhE/6SqqVvS+/mVMYL69DWCN
gTPKjJ4D0zDJmY82LGmBUmyMymrPVvsFDXfhpaK2gEo2VasEt6Af6fmZhLuVHEDw
4dvDK95Kf6w1Pc+Y2GevWl7HU5L6nEIgDCk9NWrfCwlxFRe+b36F3oNPa+uPVDzV
fIPnHj93RP0zDdmlNxLQpgh1KMm05rck+6hTCK+jRitHeCFHqX7ychjmWcZZ8TAj
5fUbJ8/YGv5M+UATMdynk1oiMql4Aeh/7vVf6CXjzSl4PMT8i3yiGdFCCrtw6tn0
lH1oZxcxHedYSP15bew3GvZS7UvjuUlNcrNlll32nZDn4qzgoMckHKY9naBTnH6V
RWQh2tCgOWau8a+dagXZIY7sVKGiq3wdzh7Lu65wGjB93SoNzMA7TwW/TZFV/FQf
+rRvY7p48/aNATpHPalJXy3poHA1rWmJzTdJKWtepcXV62ZXtDxjWHGSu/6rjvvT
HqpRZID+d3+3Jhr8sf5dL5XCSkSVmtTSWHU+om/TR9W5t4XGT8ckS6H3ebiLjQLC
YhzzO0KULEdUaQA7xO+JUrXp1mrrzTmvQo26B4zAz53PSBaWulS91T4wzQASU75c
IcX6N+2YxGKAhARACa+HkAbLSQNX3MITX4nWcDd/9vE3TFAPQgrTO1hIjGAPqdr2
KKd9uD/7cH8XNu/VgBXHHg+DlaMeeNLjKi27HYtQUJ2IFoW1MiRKKZHljiIwJMsA
`protect END_PROTECTED
