`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nqzHdRQVdwRg9QvAyDjpmGPvNgr0SbG6jgDa0Lphx/lNqLZzb60Z6fgk+AjI/o1h
+ov0JkWgXUENWAf9m1Qt5lYtCd+wdIdcqQR5RtOW2HpPPeeOfE7/OCxqhSESahtg
sIbjZR6OaemfCwJd8PQCWQ5xGrw501C9EUXKAJcu86v4zUUD3/9uMDmhQ1p3g3SO
kkMwz5TJPK9IZPEUe4LsqgPCdHSgJ7cL6fn/ugkdPQxfXLJ0S2e6P1CR33fS+sBJ
wTxx3EDNnPQsSLLtYJh3Ve03mw6ETM9IrOoJWzjXflXttyFx77tM11Rc4USNshR4
/03Vecx18Gl8U/SAzviiX5nCrYrZjfbNIRkmVR68ln27RDCDtnHtZNiwWdXlMqkJ
TjGyekAAbV2M+7/W6nwsEL14YewmpIgyfIeZaRv884ebj/cLQQcnLrs5uknv0SZn
mOGy2r3U8MgpJGggHNHnai3XW47ZHEe359u3DfngcGceHA5OhoZWLnAT7j5132SJ
iCXTbZf+CMIZAcHNeYXe2NibUoZtdhXQtMZgXnH9CvmgcVUOR6eDa9+su4vj8+zR
rZrRlV+UlcXTbrxAqzLyTEJf6Komr7yMq636SnsD9gCug/NF3OWbAuh56ApIH3Ue
zSv1n9e4iRzU5b5IqAzAoUPsnPtS+H2tbH3H6A8dVdJeP8BkHDj90mjgQi0XW6X1
CRy0MDTcPIRzFpnfb+O2u7gS5FT2XQz1csoZvQH6acrPnGjSOtmxOyc8mk4HBK4G
4LZf757Dz2UxHQ8dcLpWgA==
`protect END_PROTECTED
