`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
efCHAMe4aDLUM6jt5HVYeCxl022VQcMuMH+3Kxv/gFMM3gz381agSrU8ur9KHs41
WZpVeKxkkGhk2wntTzN0H/pLALr/v8LiHhs7rllu+Z1J4O3pU9mGDazgnSRO6fCB
6xMl8GPWKHu4UNKM2Ecjiwe3VMBpa+0vG2z98359dkwKz658Gfysw/qg/WXICaJ0
5nq7Rx0KXwgCdhM34XZPabgCBFz/nm1jYiEe4p6EfXpFJ4HX6CXQY/YYY5vuFd65
lEvjL5ZpqQBvq6YPgMKXREQGF+YxBY5SYBLlPPaNYIhCbUS77sUAEc5EmGL+nmT+
jPnV8ocvsiajMxZMYPy251pQ63LY36zDl25n8M1aRpaPLcM6A9LE0NwPcbjWs/0L
oXDi54zc5Yy8fnRfUMCZEg==
`protect END_PROTECTED
