`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uTMfTtMwzA6wLbwK0CGy8OQHDBKGgCDGs9WrtA5Spx+UdRzuKuHWobar5p/9Bk+r
nmedPXOXj23UXZVqgY44uWOBsGKSWGhAcS+TPO1W3fMHYL6YsHaOrf9d7rbrAxZs
0bM6/7FuOwJ+77Y7JsPhQkuiUUKCZMcAwon7IJ+d0YAmfbLBKNY53JMLZF2fJF0E
lc4sNTFlikBoICrN4x1KpLoNU35+gRi9OkLW8s4jPB3T9yclOovTtIRkHPEXZ4UY
BF2cL4EVOB+h6swEixjjQe5m2GvbBjrhKP7dRdYpO2teEV4TXEq/qFPDbGrj0PSV
lOiKhF8J6QzxfGWZkAEqnW6Hu7tuMH3ManKR2LaxSCHl4vDSv+It9scWEvP+SHxu
C5vVs/QWZTWe5cQs83vHAOgYTTn8ZaKUbfGq69PM0+Ea+tMYHnz4H1Cqc/y2a8XF
9fxWSeitZqCu9Z6ms75ypFh59gaj5psAmZqaJN62+i6pXwPIgUrriJkkzYd3A6BN
iJmlQZ8TkT7vqKqZihJ3wS4XvY2D4bvOuaDXK311n1bLlMwPzHmdShnPr6LIDQwu
B81n95UPVaLMdx2yF4mHHNSPjs3PmQj0a1qpxTfkh+iziqPecqRoObtcAr7rJ+4/
TIEqtMHO8x/eU3Ei61oRMbH975UoBlekmbAhfvTPbul51WOso00wrygrYlZ9e2y5
bNg35ZrdpxvdvKrkxgsBUVoICFg637IVVp4Bue8YNwIICvzgheVjoEKb2JZRtwVk
K++xkPX/tf5ENNDKm1PsdZe6nKjpylZ+idprz6qtNMNw4HF1p0H7CbzDVHwWrVIW
`protect END_PROTECTED
