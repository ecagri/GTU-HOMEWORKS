`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gYPBlaTMNAbT1OHCHwH2QVhbYUGbRhxQWzkx0M0EHbf04eWNjyZsnfe/ofFi5Ehb
AUZa8yKnvi4SXi68YpG9XKxiveY9nPwqgQBUsvY34kgXOkt0reBPoq0TlWwkCi74
uP/jt6+zsUaijSB3HWdLTVQaB3Urf45neYwnnr9b2EOwCPj5V9oMieO5UU0vt3Me
I141b8jZH4kcNVW2x206dudpHOKpVYzvn6KnbY+0xrLI9p/W36h2QYT3e/Y71L8z
5mMK8JbkyZDX4FsILRHP5NXMKBUiAKu3wKBsgyCVgH9f0Z8yNp67IzcxUQQwFaUp
p7wX3+OeqB/2bfYPruFjzjgy/cbr3+SLOdThSt1aboMpKIYLfLcdOtyr3CRT/O5q
88EeON0aiQT3ijFW8TrFWsyzFlpEK2sHsWEegcx5gleM/ISJUJtYV7A1UpXCCjHy
d4nr31aT9eTmUERe4C6ccLUWaDOzOvpWDuuhU0OCMmobj7DUq22hsJkjdicxUfVb
3XwyYo0meMHhwcB2IOtpFuHdBQs6yqZbif/kmW3u1wgyBeg9egoFggUIgNCFY017
KdZCyryNS2uA1Hu0ZUJ9QlZW0rSV5h89N6ecuiQndN1Ep1hi4boHdui9hOTj80IX
f4WdCAO/eUlwUYNf/1jiXIND3vJLYNHkosNKl85Ics/ix6ORo0o0nBDJfPND77HH
bTZRGNkvoGRFJy06x4Swwy+f+/biBlrGBsfHo9OrA2wBzeDsZFe1lfYGnXk3NAy5
2N3eTAOtnexuCu6xChMRf90Ctog+RBuRmMfptdMo2+l3NQGqVIxp8lt5oFzAb1Dt
zoIlmFPjNCGVTlh/Q1hEn0tM5efETpN5p5r58JF9PYo7VmQAP524FJJjMDGs+kK+
aViwOOXMIwjZmub7CB/86xojKJXFoIgj7yqXOivB3XDH9khb1otbRrNoF/hHaA6L
YMtRBHS32V8jR7TqCRk+j7ZQFYvt2EDk6bTDWLcDHJAa4+7Kxb+2goAcDZ0zfbrV
f7AYd5K7rhk9CZzz8vvYaFMFWQ2u6DEzZ9cKUJO9iokdFuc5ibR8Of4syztFIknO
4oHouSRqGrCQHjW6kekzDDpO5HX7Fv6fBIW8uVQZkbyEi74+gdz9EAHnvcMce/W+
c1TFuFf9oIWSRGHRdyyoKs1i3jn3P6kPzWLAQlaxFzZ5fvgroeOYkSxqgzn3EYFK
J8LodVrN5FKk+BNr5fyK+xKOvD/7sy0EfQP3sHFpUiAccxJndu3LHs7eUH0wA9Jn
tKDQnGATOz0gUHGnsA6fgmaiCEsEzygjYCnboQKim/SSQgx3gSW0D1NXBCzyUAuH
WaLb7SleOE3TJkfGG23X9KGkhnNY5FV7DDycaBA+/Q3cjWi/DbgccYemvpSsB0Rt
xhyxBvzOv4AUEOIFkuRnjZBXUtGupEfOTMDYrCo7zdwFlb1bYt9F3Req/bl77Nje
wjUC4xTQMbMjjTA5dI7plQEi7TbCf3dj7AuwykfylVd6KbkVotKTxkODL/GjC7qu
DEsMNDUHGqMetnKhj4si+lfOZA63VJVctGuKqBlm2EgXa8FMfXrLq4DJLEJNfq1p
2TGHCW4A2Wx9zZcYSbMjC6wF4dd6MyZuFb5aDOdgZdI5Pt0YWAtvQ2I/LAV6KMrm
MQoWRy5olH+mV6eEtNSvWZ2NmTtc10J3hMbIqBnaFIbp3VmyFv03/BtT/F7+OnuG
pecK9Ilyt4fgtRzcCo2Wy07kps8HgS7Ne3RbL9t4JqX/RfDF4ShAnc91r+qGdhpR
PZr0kpzvJ0pgi5ESEY+ehYT9zX7cPGkudquIqnK9lR1tBZTtonvV4XKOpQvxkDLO
1ICPB4rQw7f4XQIdOGvCV/sTpPo01PZ5sKNO3mMXU7XJAX2ghB4YDyRCs4OhcID2
FjW692hSdoFbLN9ZEa6QdAamhCizeqv/e+sxC1Lab+5NDB8b2HXlIm4i0weQaNiR
KbQYJUByyLlNUGSQdyEKRG7p1BLFUK4xd1tMAw56HYWp5ulfZdkE4E+Zwn4tClnB
Rh8u6/G4bjxWnLUX24h3vvPlHnXaac4vbmXxJX/MjR9M2XN9ldrd0JCIEU8dReik
hwe7DnvCe/vfzF/au0lb0hwZ35vveZYTfPpIJ+DyaLoq38phnj06LvwxEXRLLUYh
fzqu0OoHLUS3r8v6mWR0tyIJfxrCus+sHGEKc0x1CZwPLcgu5TgaBqcbVY3gDpbP
8QQ0HNNDTAzmCnQtye5KiC/tFrarucemjLHYwk585GiRTQA93F8ClweOJb49I7yi
whEXymNYWdZDKTYiNObOBGAhrD9pKSyUrZkefPDQA0Vby3JY4PTlPh2j3S5nO7Xc
hm3fwtuiIDYGHYGv7iTcCdHJD+JeOtYPyRf1ZqNjx46hWBqYDnNc8uzp7K9h7UcP
MxKABjg3Z6+F5I0loxck8H/9rmvTrQ79N6CMIGfmtNpZxPOn1EyETKbZRdGHHcit
ba15ZWTbMCpKFolGwwWYCpFTFW7SXdkN7gVprPa+JRBlS0ca9IAqCkffNoFI9HPA
v973IXorVK2evnjavFfqTWNcZmUdMqYIR2Hk+yrU6SbAOzt21vVHwDBjQYjWYM0W
SghHLM7wXg8TKyiDbaAe2S63SJhZRBT+pz65MAIvOaR3uIMsgDwbF4ZkeBIQE46J
YMOg/3HD94C050RnqLh2DBxwjLeVkKYXWidb1er3//Xk6Tols1rr/2BT9xFIT9Dk
b8KoMvWuvzjy+fSvJ5lmietCnw0EN01f6BFLxnA1iY61zsu/mkBnwLxhMZOVPBQS
207JpO8m8kZrAleOePJbvjH6O+ww/v6wRAaCfb7G4DDWc4Yl9iML+FB2CspiEf71
iip5agij79jT0iWYcjYIix+gfbrjiez3V27diJI/+iVAqJmCNVgAKaeGImEaVN38
cDE6ugSuKzZJO7NOxseQ/Kfj+v22UGbtoCLrH7Q5PBtN00rE8bF/i1BE47ewW2FV
wia35zrP6ej7Ylbmi+uIG6DzTCs2uDUgGBagPIkPYExiAKLmHA8wt41YiOuH1lxg
D3IStD44uRWFZuB/xhEEwp7mVbHRATYBdrYILzzf6eVn2nROX1V5qD/uO3KmbKQm
fwYWikU9XEiCrO9qUqsx3CFPjhELDt+Mkbi76XAT2AYorm/udgnG/PXAcKmRyJA0
mZXYhZqn1jakHWKszUiwN6XinMNz+2090tdMdBEx1a2lSQkk7uds/iEZcM226MY1
lurrY8cVG3xUunJ2HDKViL88Awpj4tuem8bR4NDEcjb+5B86DH+yCX+mqQZnoLm9
yGHE3ZvWJDW2gYsDePaLTHJGxYZmBWM62GepizZg5YSoBjvtn3OZohoT7pvK2KtL
Gw6+OaWhqBguVn24c/+azKWxDQGF9OSUral/Qo8qx+IJkaKk9ax5Qd7j2nu3rPdC
3VJchm8qmqC9V2wnL3E5Rxgl6YBTSWtMWI+LO0VvzLiaeOaZNU3bDJaMg846+zw/
i83NvIoQhQ2FetNDs8JaGiarRmKvM0ybUZkhmY9IvVDu3Ho2KDJDiN+YaenDtrxk
+VuYaDuABvYRt3JT0fiJP+Hm8EAvskwQTsZyjmn88ycJ3ND/Zt8eHi+keuH1LX4Q
nosNcWYk/sP5ERpJlXU9XebCfLiHONrZhYj+Xc9AxBJ+eXQc8TFOoeIZC/ANdJVM
DP378AO4XPNu98VxKgBHJ0wyDLE4mhNS1oysPlAPflSM63T7ik+eX+CqQCfpCO1N
qTkrhkudpYf1KwiVYRPeoeprepIRYt0bfzkBoTXmZ04kBcbfozaDRzvgjWvGqZLC
54+OrJ1N52o+rog1Fkj32E8SCov2ouLdEfm9Lnjpd1aQmakwXdS5+ampnpmBuobv
MZawny/vNM6OLnzcWFfXuqnUspfH4gWGt+h+mwlXIlNKxMjkSBhKVE8UCFh41evj
BvQQW2lLvI7zJq7Mzk+ik1HCHrz2rFgt26FHFxDrO/+uPcMLQuJZOeHVWTBxBbpR
SfxeRgPgulRHrd6d6Hez4A9tON12zzaPb0NYiEZoWstglcqRUvzw6wQxHdXd51FE
kZIbi4zOt/XbTXbxbDXX9Vsuy8U3Kc2/D6W+1np3tOJ8M/RDPZ7biM1nQS4j0WDP
jadB7W+40+U4530SUUDH02IuYFguvN3NJsYBrfVlLjP4gAivK/AuHailo4Se4171
YQ2VJj87gPrfUhBhv2BW97CWgo5Mjpxs8x5XSAB3AJAuy9c7S7AkkREPX/M9KM0w
lccgodHSqHNM3ay0w1WLzVcx4M7gfgmC5/KiTRq8nfP262hYeBNK0xrlvOg9OeVm
Y1ur5zhbi82qjHOI3HgQhsI7Dy8l3wv0UXXoGVoNPkehHQhAKWuIJeo8MheCwbXw
hRMtsh+MyZU38qDaVJTjQl/hKAFjKqxxXAJ/6KRVQVfBQCWoXiBYp7jAUxazwICF
gJ8Cck2b+jHdEsDdELFsOfuDK3e80bHc4xzKbeHJkoEmPhPKkxm42HMWJ5sEAx3R
RAyvRNmRf8SqcwRfKlIxM1ROjB/XCQTkonQcuyiK2UJFiLjfJXDnI0CXzz7KfNdR
+wY1ewdGKj/JFcHSVAhsw6jQoLzWuwYU3s17DHL1SJwb+Daup8qV5Y6OB1Do9HV6
7o2smXaZSGQUhAt7iRDHVjOAbZE0PM2KavJqBfI3YIQBpmLa79z75wdghtQe4l1b
MOnbLewPSL8fGGzUv45eLhCoC9sbChWVEgP63/45s8W3aUT8F+7CRLNRXsCuXgJS
Rcfy+MAf24I6ZvZ/ig5hyHn5httsdY6dXC4LmcIXkeDCg19QmAlY9WKjKUXRyVwb
M+5yf4/bIOvU1WOMYmNLdy99PrIp0qZjmqi3G5+uXk8erXkb84iUky54QH9jVu8I
x+Aamy6h+/rKM3tlJ/eiLJUxSRYqmdw/A9NKv552yb8uQ2UVysCUsWAKEcHJZWF2
D3WQn71sjc2afDyH5akul88HaEN9epQ57XUyb8Mei9f17Npd28WHlF5Yrlw/YHI5
h95dUZ1P1kLyS9okrg3zeTDcXvDZESiRkX/WDWMwt77xEji6L4jE3aLYjw687jKL
cQeDpimkQ4kHssrM++XuFn8xEt4pV/UnYxOUZ6rRT6NBMH7/asMJPZTF8fcOauHG
77afVKcxWAs/yU4TtRjEMvl7dKEz7ypb28pVLA2ymH3dHeX1lDccDSGP/j4AZdL1
xif1BLkmN4c6FL1kZtVezXFN5bs5BgWfUKaZmJkUYO9b7VCnW4pUS/BVbFjHplo8
m281ATPSUWTbR1cYdA0qXCEo2SiBN20rpzcGdXZUC9QGVD/IItVxPXUJnZtoMdIu
Om/9D1u8b4A7+XFzSkzst7i+Ewj/54Mv8lRCJQx7uQvXVRr3mlXBA3wV+29/NLBC
fN/1iJMx9dHRcwDkk8dTFA==
`protect END_PROTECTED
