`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vkdZkLkEKL7jkuJuZeTEAi5XE09cIHJZXWUzYVFs3vgnES793oyVaubgX4BsdMYw
WCbFySGldIx7ZrdQ1JnOVLM26CZwFP0lfqtXPrt/bJxOYeh5JLh7tZvD3FLdQG8P
G9k6Yt7sQtnRrf1czDId/rsvZdHLU0FYGoWqCfJqbNkdsPTDl0bEgFDc9XqpN0Df
TtHX4GV1uYNPTIMtTYS+fZUzXd8lVNmh71Gk2JSr4aDZbtsCSq8jUJC2eFcFomGo
kQjJzlJFd/liNGDpeA8Zpqck0gITP31aJrWPKDa6kZNP7Y4/RuwdtAE4qDdj2dtn
4t0iZjSfSs2/5yVIta1L47kQp8PFmgda2WuhFzqva2sh/lxMe3oBU1Uyp0s7QcEQ
1CwgWAiRDwYLDsHnQiltJD+x+ms6AYH0flJ+tnOyBs5Qo5X6zsK2FE1QhA7Givac
DSVmswPU7YMTVuhbzRKxtVP/iVoWXs223HfF5XP6x1GAW/45llFt2y0CAGqpjGLA
gnFKc+k1MfjzaDF6SOlZR6BQkC7x7Y0etidP6kT1cehnJEjOfiyUvYU/okZHR5Ls
k7Ee1L2oYo7IjL+thR6OWg+vCxgtu992duzqeQbWEH91RS3OOD5R1fTYWBqryf6B
04URCO/IlSqov4uxzqJ8DkWPA361OyR9uJ4tJn+oT/hhgVThbByQPhP/KTa9Juh0
RpFI7or1mUZxKOnNDRYUhZpS4H7RUDIuXm1OREgWGeZtKSTS0tWMwHS2N6R8xLq6
s+R5EV/qTkYk9P9ilZus1IW7UICW6zQgzVOmkhOs8s16ujQpZlNymD2YaBQGrUCI
39/Z77Rxa8TO+8I7Tz76HjNEtF7BaeopIbEy0la85MfaVENGoRzFH6qS7VRFrmfK
br8x51lw/vt4bQrnIghZdMUodNCKK2m55V6JiR7vs41BPybx5sh80GIh1JYFyGKS
aM9YC2cxdwpQsVY+JXo8y4aRF2yWYdMIDTIp29crfEk=
`protect END_PROTECTED
