`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v6hTzORFhAkHU6a+p0ou4ViMYaC6m1tKkTNoZWo4LfiiWLv/yj4Fc1VGiBHkKiQ/
I6MO4p2DSQhNNpe0fwUQRp5q2L3S8Q/5qjXp1BEOecygypctaKAcqdRm8zikBXUV
JW6g5MCoWqXnAMVqziyIlzZvf9E8icaDWaUB5l3CJf3l2+txun4iFToXnJOjjB0r
3R8A78qP3PhRWFIZiIrGZ8/AC8dAamcvEjU7OOzrr2FbmNEne4zR1Xc/vGtVfP6A
W4+zuHpLcRWnCd8oj+8mPxAoAguhoBFO27c70AZgZYcJ4QDuOmgeOAY+iHaLtgAy
ZI0h2E6JYreoTIO24JDP+/GP9y9akhslUc5k4HdnTn6/KjqbpfCJewhfI7SOUYbE
kSLE06iiuAZT6nJiGn5KfNoE8GoRvnr38dRY6Y5dCKlCX2K39pu88IeGcGo6pMq3
wtSe/qYuivZIvaNRE3p+95256ZxuFp8WSYUwxHCYZwnkhzhGvwqDlQ5hoebZceYh
OSeF5euf5953uRgx9MGuKZNvvxAuOw/VqQ6M1HcyEsELsaO/1GZBBq7y/J0nQmp4
CJoyNBC22Cfj0rdMYJy2IecuM3KmyeJHsIbmcR6NvpSX9kqzfDBe85Op3z6BIDuM
4+VnwN5YuFwfJbBWIvelzOc5Da+PyXMqbq3AfZYd0SlOyc92xAqOlGt8UPbfNUHG
MU+K1sFKjLgwNklLPNK/AY3vUzgakb2T3yn5jsUBSqGMrSqtX4U79DDt3WXxokuj
3RFnWw1y3OXiUhQ20WIlc0fj2arV+WZUF3+qcqxkepgCUNuuiHXMdCKJ/9ZiXNTA
xjgvZQV5tjXNXpymCXYYg6sbQvHaHrBvDaqXul5uxhVkrT8Rx71f++LlPsxk691D
UeZDWUOEEs0OT5XDLKwsIrrHX+CiLDs6Oca1rWHBQCFo/YggWSscKg3wm1+uGf6b
Mk+yEH1X/KQCxSzCX/qhFFlGVdQVvI6PpNyXCw7uy/UCBjpbyXuPwcLz1EB6vev1
hmo8WrHLj0dmXtHaH1bisqxddRS6rn4fYPq1u4XQZwzboNiBMhN8tw4NvftFiMfP
KwGSjFTuQIGRhgBiISRs6H3Tyoj7Nwev2hwAdq2IQZI0bL+Zn4zb478TjSXsi7xP
D+CY/QnB1mB/OI43Koh1xjfMi2NyXX7tTa5uh9E3oPAY98jHKOHnnU023vjlrUNj
6wrfc++XQNmz5J7qbj/UIhhOw7YAcQrCasMzVODUYQaLGAVW7thM5S20ZJPSuLGM
th5ES5A5lIqFs5LyQJwJBihmD4I0h1YfRW7RQ/rJVJdX9D46DBMe9CCeZqnA2z1q
JkB7E4mOtTg+WyRl+6eZtIz8oXfNyL2sTamTxft1/QW6hBckAAK4oeetUN8p406R
J3h3VlnXfszH0SBkSViwMTFiZE3jDkZDoOfSBa5Kk5Zu07cwfRC+07o4K1vKg9OG
I+EFL0ixToCDbJYjzrRZ7ibYFaYBrqlEkdXVEM71b1acSy+G3HudSHT5tEWG4oyp
b1giGQyBevkXwwvkRRcvVTgIaTh8hf7ZIUtKeEqcsfXXvhd799N5N73InqY6K3wv
oRYnTQOZiDDimlIcmCfoSZY1oihyLLp5Y/gbXc6zPWv6z7r3eHlSGjGA1PXr3d/8
d/Z+KjrX5AAQmXhOFIpsmBiDvLdx1yD4Yx/2Z1PU+gPX5or/2AxmtmYWNIm/lBIP
bP3XolWsCBbO5INvWM3A9GvQ4C8+zq/buP4zL8dwGvYof5QkdNFKW4NHjwEYJPHj
+0jKokXVNsChE8TcNwCJgbKrecXgOYn88lfbabQEFaKMYJDqUqQe/AqLEjN0onfI
3Bmw8xU4URYy3k/IBjiOCDkLWUKQVFbWjBJWQ4bXC7jUn+6BAjV0nj1ALB2m9RjM
8yAHBITxJFP+4tpDnEYJzzAIHKI3N4Gr6kj4OVoaBIFFz1U4Zo4FGMi7jZGBtfh0
ACaHzgJ+WtCElCMNPQ6IhGojKZ7DZH55qkbTgDW1CViUEQbcz/VPKTSD1t8/tgA5
tNbcG1FoiO0iZWHX+mUF+Lt/w29P1ZOB+roJJq4+ouzOyajWLz+XMBo+7/hfc6c4
3pUSsIwNRZS1qphYvC5COWTrMo1G8LCOZTCqBmci5xVe9jr6+ggbyoBZgpdOF+Ca
qcTetc/xXFMU12rgNzMm/EdJ5ZdQzpLwNzMpbzDFbQaJ0qhBqVA5393m6rGQXpFj
6THgh6+l6rvX9GBIRx7leVF3JmLLdWrGNyGh+stN8tKwc0H/Sx24hu01pzUAqeeI
z5K0nBzH/nmZjeKEdVuRnARbYGTIs2npsIqF0PCn4b4drFv7OxS33IlDZQ0WEPIt
YmYlNPJMx40yi9xuXOKIO1f86WJtdWdkCiPX9j0D0kX61r8co7N3qMus9YmZbvTw
RFUvGfy+gRWnqAEVHHlIYn/MnPk+bB0ABu8N8oU9jUlwvFw9Ahoo4TDhIrtTmejR
BPjZTDwz1MX/APe2cKQaAWMZPTIbq2XLoPJQbRAxo/sBcMwO0CyIvY9fH5gStZja
Sr6O7VwgKwUwDQA3pu5TDnxCD/MstnJa/Xy1XWaO6KOAmLBRJ12BuOsfTEh5z6Gi
4uGVrdWFPZPVUHdltIyRrxW4L80VfLNigpnmeRqrJ3hf/o855ewnb6OY6n5D63RA
0MXkW6zGoqC6TKkxTPZ1X2ggXNMj9lxehwjQAAh+HrDDz00X2pQzsZc5pxjrSSzQ
5oTscLbGdoMpw4vGfvLAFPBtdtpQ7MOnL0DKTLHre8ubrMVreDCTOailtAq4Ey2m
JJD24/hzJcvNHfNAr0Zhqb9BOxr1uio7vFdOml9hpXioxUfjb6I5LkLgXhOFUT1e
agVmzs3wNBbh0pv8Y1qMwdDqwEzSR20iYa2G6+UC/t83s1YmGXPOdDMkHoJVQDXD
Y7pyfbzHol7g9bpcXnRhudt20GqAE4VuRxByNNjj6jq85mc5t8Ve3keQQOXOpW/x
rPaQ6CB/zLz8L/XT55Dv923I68Q1y63b/znTkGyifdftVwn85xD/FKs/ZBxDP96H
B7jsRMf/DIDtSA47X7gMRAD+aBg6P6FKFi2cRDeK9Noafa0gXPI0YNrb7ElyHAy4
qCEiGW8n2dsFmipm3rv9Gi44itPpFN1eNU4CYqcwx+vpq+eEM6dSFiSTdCqx/KYL
AztF1YyKNmvozI9rsG0bOUXuuW98OKQqgZGDZEqNY8piP7fC7Qu/gnVD8rAQrUY9
TSyK8MLfb31y9fpsUvlzlU36nE0KjOzjfL8B2ij4JQt/7ukgFT43CzRClTwxG+TW
oyVD84WsEBBD1i6+euTnsmtgjwT0BkqDrVzYpvQbHlcfXlL1KOO0BdpT+vCOxZRh
7eOaDwf8KLpiS7c7TpKZnQEBaox8FxQZ2rqrf/nmxLRBjLAwKpw0ePnakEaflFWv
mAF2YXtiyHpT48g1TyHtEYgkhp/up4Ph+SYdVt/eJ/mFyDxLf8Q1sH20mGJmtIlz
OziTgQ+WFef0KT9BzuTm1RUzuohu32uym5UR9YogqlGkep769ZfR7H15j9Zvl/SL
6c+KP8KEDsA+Qmp114/wZRpMzvPDi1oT325IaxEb4vJkHtZ1BC9LFcv80yDRZvfd
kG3byjk2/BMNC3+l3zxXg1HNYPzx5QMjGyYyvW3xdoydpvzHAPRE5+g+Yc7mYoHl
T2T8eGOkve/vKTdUVeia/b5EPS+koy+r7KhSHyVd1Guot6cf/7FrNnUiY6ec46BA
FAMS5ASLLQZv0dsG+QsblV3HDandIDcXJGY4AvCVrLlv57TjdTJSdemCnz5hrjAg
SciKf+yse5VYQ6wWstHRBbl2HmxMHMKAyloVJNFZx2LFScRzc8zmusZkIZs/97by
pYINa8zs68dD8BbovJ+cJ3wdRH0vQpslJzVbMsYxcTPImBuqT0fIFxgAIN+C7CYy
NM0roLI0yL6uj1tdRQG8lAKih4URTR+VndniCPaoAJ0OZlUbVj+GViPr3Axt44JX
tYlsCXRlVkrIiNCBYkmozV8B3pvlDAdhBx+VJYspY5Ak2wceHbSu4u9BBIxl4eMu
hkj7CdzM1pc/sCTgcbRDroSxGb2S3wSGTpvdTTPWKJF14qOXmNI5zzfuzflQyiPl
j763r0je/Ew+qKqa6siFc2tBQYjI8FScHY3GsAYEJndd6NuTMAubL+vRdjRdgdq3
UjQ9KxanlOhkZ/HOOm3X0nmkR32VwVAagmrQ7QuNGx9pctybPMNpJfeWFx0XqKkr
pHif72Y2YWeS+n1nzYu5pm1ehEOgADtVXxIZinG17w+UPpLg9T4ztSzwvfbeZBSi
N0IBBbXtsccQkmbN8/mYaHQsCwXpVgc6APXkWufE3MxfKk04FIVg72nuBoVj9nIt
JCa8gOyDGGczonwMJzhvaAEzEcDXrEIDPXGRcL16NtQYmfUm+wokgG4EO4gRND9h
8EHdF4RydIKehaIY73kKxtCAMl3SzHAsNLBByJKBwrV/TscmYpe5T3Q18IfrfwIN
o28sSzctW1owTC6/esy1HP8u6NRSXnpQGKHcgdmQZt3Xrh3NEBNikEqi6AN6IpOd
yPlhBbo3jh3b85+wm0LyMcjkkYp/S0V4iMh9B3iiuv2POC6GNKQJ94y3700XZ3JU
1bwG/ha7DjfOnnWBRwjkOXgWk/E8vFG1mzrdcu3PcY1vpr19qibR4Qs+w3WhfnoZ
CLgSA0zsgJFoFMIYKaFTSoYPBRV0cFfxOJ8OkqPD43pQn2x8b5BhMdLG2zBSfPnm
YYcbpNxm3A01VRoPIh+ATv8KPhcaaPpzWxdJoM/lgk3ZORihqs88Fm8UGp7/MnSD
nL1HR/vfRULrje5hQNL2UH1Ro7I58vx/fFv2C9yE8mEDkADe7h/Ba6r+WWzmBx+A
xMqCsiybhFkMd+aMA6kgmJ5bSwpcqL/tKj0cbCW71YOld8iyS3G6VVKaF9KFfFHD
BKX/LRzye4qJFC53MXu1CrLdkZ2o394WIjfqNx2aiEpPLxefQ57Er7pGdEqTpFBU
QTN/gZZQLowBYqg3PYP3AA==
`protect END_PROTECTED
