`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MhIRd0TiocsiT+zZpliJpbK5kG02Q1xmVcdw48qGJRa/0ZCPLUR4TCSu7CQyC6wY
CfGiJrjjSHTsY5SQNnm7/OpDgt/MIF4N/veWaxfgoLG72F6by6vTDsmGAOl0E8uP
B1zTDQlkztX+Fic0QZM6o1rzw7fy1jlEGrsKQeuewYj3z5fAZ7wk6AS9l69vow2a
u2wgMcVWQNmP9bgCpacMO4LPmL81LvyIdZTEZs2Z3KQU7MkXHsfM8FTk2CSL2Pxc
17/BjfwlN71lOV5lHXIFPrncpVwL7CjHk+ml6DneAKxqWky84FGTbyTSaDV9M0p8
4uXKo6kCCZeiBzTrIzuoRW4q1OohwkOkREZ+64eGY4X8n8RdeGcuxzmVWNNg7nZ4
+1noku3dSpmjrV84AvCbBVnx6i7tT6eD+4Gk+pBLC/4cDo9IExjNO/Tre0rNXupE
KqFbZbBkDVYzWWfp396uhGZ8B/LNfhwNwGg1wL/t00praOBsr0qB3xNtuLDs+dwb
TLOWWTgBDI6X0MmcHAsgCg0yDrRqD8CyD7fiWmlwke5UvsnWgUdsgex+HoShWM8S
6Kni4qUetAUKLurTDnLR8MUTOcSBzwdHNIE1Hw1YqMDpGB75OWiNXXoccdosM/5l
mypSlqwzC85XStkfxrfjJj9zexbnJvEG6OrEffvTz+EpxfsGFpbuPKLb+Yn8P/uV
z6uFqlQxc80/x6BNZ8gtgjGdOZf8SAXQQdJp0GKoypEhTX4FI5837gqoPSuwJRTt
/WthE+upid+KFLX6fSYb2vIYskB7iIzHMSOGS/LclEFhVuuKFV8JY8bYghlTxR/5
7tfoz/ya67eywpvXclpfrotBkQAqA1vx5zIYdZ+B+jR8OgWPmD2tBK4BcmmYIIJG
MLap2jRucNiy9c2oaVK5G/7oG+nooqPtJe5yLkBbeYQqKrR8zecOLjJcGfWJm3HT
RpyR7n0DX72s8prQrz67KGcw/AbDyn6lzkUSwWyZmRxKc8y2xsfJzmftxEre12IP
iELQB0Sdfz+rysl89RgPXb/Ndf75hoiGK5cz1ItWmg/f80l2id2wKEUpMSlDw/Vm
FYfJWaaKTJZlLXVSbMlXR/UHDASos8pNTojZWeADm3hL5JABVvzjvJvjoJKweIxr
Aq643m1BP7k3SHpgBtjvvw8yiQnlfVzqXOUD/dIyCR2EAe+x7OWNfR0fCTnUd5Bs
/dqyA8kWjGUZecl5Y4CdZXOvaVTzTXyvJLIbboxr9f5zsDd2qIXW5OrfTO8MyhMb
3mf+ShZAw1BPnD2kSAGHrTiuR9/387JSZMINRT358L7CLi2QrKM0mdwdJ7HCs91A
6mKyAcQSFTVv1Qc8AjF/DGlJBKAfmVtq0LmJuwQzkE6ftpwdiOM4iiF4qQWjrZrU
BhR6M0bqpDQHm8yaED5tpxnarNoa4ioR00Dq1d8J+KjkKnQNUrWRMmkAIGx5Ov8C
Zw8xqXx6gVNvxo8Y6uM904j0FO/8JCDaaIosfwxA0+7T3yGn1QnanLpzhjtJe44l
0BQxyskFtoZpsphxUKooCnorbajbNs1bTlWl7H5q3rGp45rJhESY/1RkE1iflmaO
9/6GK07cFlJtBgDBWRBFi4dyg58DXumJhNMlun0ZTQGeBQT7mZCddexgnFfvOc38
09JUPlWhqP9D64sG6wjhvcE/pLshUTjmJnwJN/ErETKhZCXDGRhMUUAOV0BnEvEa
VC/v/PZtyqhZjOIg36bjb80Lb9ToxaE8dOKt8XFKYJXoQ9IQsJij95FXbQzdF8l9
9rBQVsdqkd38Sq+lN/ixj1QDRheKfoyBrs1tPF9JuSy7Tm+FKI+l8x36b0VJSV5W
PDp8WNdu3/MAr0Aq5BtvtvttKzp1RroL1ZVOu6U9eP93rswVRD1eJQ+bANt/Lj7b
vVld4Vg5qIqCeL1hZQVW6gfdYsCfh0Wio19t44vnQnwc9fW1n4+Tabe/xG1N41dP
0VTBZUJ95Pk+9mynRIraBVsJpbMrL4ebahxA5+8LxPsXmAMBH1V6ebw+fklUfTeZ
2FnPjOTHcs48SBO906GhcY3/3Vj5CZpb+MPYD/gzIuI/25TtPstf/i9Mx1oQPfRc
rJueWzaz0EhNBay9kTC9RAEcEdlXiioSquuNucICGEkM3g8+PbsT/AGpSgvgwtWG
uI6jRjdwPkKSJReKzRBnxfIvLrFkVxm3+yzI0D0P82b8ps1sLCp4R7xNbb71eXqQ
nNrbrTR0FLLENnEP6rPP2gKrK3XArO0EjSjFd3sizhv3ESCXS+viABGD9a+AZwJT
QJHNz/UtnbLuz8m3k9m7s0mMvJTNtA5ZQ19jWpKUkBLUT9KtdDv6kImhPNmSL8TS
OxXied6w0rGl2rSbIWyTBN5a6aQdNOEdx+dQitM1iIQLoyihOSycwA5n6pn8K/Be
ciRScRKJB7osRBP3dfYaAJCoshNvKuOH9OV/VYRQEjQzffB9d3nRkC0mULGG6zeT
3FriO9OxIykMsDGB6ipzgb3duHXGpUArqnWzo2ySbTJeonOgntBMHvEwRMEoUm1C
RYsN4R3BEdAbSn3oP9EdWWp9SNFl3eZYW2XXJgcD72r01OStuAUNZhehPuzoiHQf
eFJDwOMIXQqqzp2UBWqcethLOxz8w533g/arIaVn1aLxYjf+8g9mA0wfMwUaF4LN
J+WwuqfcWfPMU+ZVWlkT0iGg1XU5H8DYQIPfOhvXs6OUxW0l7/3MeEq0CmI0fWse
tjD5WYebG1SuzE3DLI2vuZ0u4O+9GFq3xOFtT8YkBLb8ObkGxemVMJjj7twqdFS5
uGZyCH2XyB1cfQj6hTjWRwe2nFk1hP4EyXRCSe/IOuGOHEAcis2bHbrzIecVgEnG
Aong1Msdlj8N9BBKcqN1DiawCxTr9ZEAO3lgCDz7spcCQBDf6LI6qk8IQsqboVBn
LgP/oKxhRK00QAVS0iekGu5D/QK6XhxtUIpEDAA4DkfLd/cm2LvtVOEeGdpBDotW
Ip8G9/QDQk/PjwDiNFzXKBAfX+MDgwiKunyYrj5lnstM2ZyuYRSSNuF/4+BPAbWk
akJFHgG60T7sEtAL4zHN/NpYyEcrvJdCdbkEfK5N8DwQiWY+86+ov4b928Y7iBe5
Ixj0MNkqdJUimyl4g0aN0At7O6UciwcfyaQWg3HaJtZ780BxkEKRa6yY3j8WDWxl
+qcITZXrPZ6Qjk3DJBSSsLzXH6gjWD3YbllgcCk35ctcmEXLwK/E5kglv3Gb4mfW
9yjijl/sBSakAVP+lGJaEfU33qDB1kcsEdFeFLOHxXS04hzd+pK4RnlKEn/tMymd
xHxyT1IPIOOSKZ5KSSwsUJH6L1I25ajV7TT/jNKJiadzD1nKqjUbcKy8Ks0+Zjjz
AxMVPuzUnXbfy13VUlLmL5lH9SXhF+r9UQO0/Pte+UOC3O7P0r6Y899lXl/NrhVa
pSdI9zBNJxUq5VLz+kULcx5ve4PSyeSJ90KK7XS6AdeFOltxVbwLPMQDBCoRUl5P
mulCYtaLGpbVK+ZFnFUkdRBzcJTexop/AVictvjnO9HWzlVhQD/63w1LpKB12S8m
unDcEIp9sbsBfv/Ci27KreHlcgI1kj9MvrCdZfgjFN3aTe1bQRex2UFfkSeRPhXU
PTeFrS59MrqLSXr5JWrwrVAwZiND3eRwPa7zw1q9bSqYI80wqMFFPeyO7UONRrF0
S5RxcpeeagPk6N3lOaggVn07nzLHI7mSxm8ZQpBMgGmy6FIULFqXAqw5Wt3ZS9Pl
lTTiSDxE25GBnooiiMGRrt/KSp8p6CYFSlD2FFN4rY1MOb+BjbMeKp0kXm1C99x8
JVLgEGk2V5mLQNNd5rFeoowCid3UahMsp8ZV6S5Ypssznr6iHSNj+mrWIYFIv8nc
zzfATk176eRb1VCdlCM2q5GDRXsNVFn4vkqoH73jIQSi3sGU467HjL0JHMrRgxtm
mU1X0JDDPHFfLTjGplo6R5isHcnkpVpfC0PZP+VMMmP44YNunRpVeahVBcVwM0s2
ICaLu/b9GNKZJhTRtq1hwAPKoelMxbqQqTiuX2nfOjhW2WV0AJZKsjkUWb6Uo4w/
f7m4kq9OSKoLpTDbG4irBrwVfPTGKaSp3jc3e2Es3/fuXdz9N4a8lzh7XEbTXria
QdIrrh6SSMuHWRy//hX1RGD7B6BjdA6gAyJS9BrTUtYd7lnVsjfFclgA4PgYJVfl
Rl9ejgNzDoV7Tooql2nVrxDQA5F7dAHR3cqYGFHMKOyupQK55FnPmirXxXrsCqli
f06MjCESZxeGigsFztS1TyvURM7AYCjCZ0K3PrQnt3tBzSo0qAmbS22dGjigu9/o
17NpsOBECvj3C+QVzJi+zmMw3yfg9huh+/wLVVofJzn9i2f9FebamQNDGVcXFXeK
5g3XDi7ZftP0E3XvDKl6qkkE6zLJF09C77VwSST+psh1YayP/vMln17iNSpZxdnI
g3fGalBlJkMbklXxIBM9w55Kedrm/46tXRpojxX4ZNlYuc+SucFQOwywuE4Q9Uhy
DnRevmggPjrx3qXv0kVadE8Vix4IouA6y6/OWKGHVgbr6S7gTtUui5u/eNjkepWx
EhJnr2/c+ToVSAot54hKtqclodpiwJ/M+13WYxPY1a/X/CuXCiP9oKqIB7pVgDOd
2Pz3SqVXKDMFdvVUrERt/eDJ9mjsrURVUp0z0jTku1/LRzIpDlx6WV6nlJ1oeibp
8XGdZ3oa8tSbFKQMKQtcWYwUp1lN14QfJzT5l6aB9jyxqmsfcLm6nysNeEosovoI
LEWeSLgsTcENXFd0Vr4X7u7NtPzCtaOJhTLDI4U0YQSd4yaL1UrUuXTlHBD6OsQX
0bSArEM2NEjXzoZl5k4Ql0dakknLRHxXQnJlzAj2ECfZpSq2ZRLnVCKqqpOP7WAl
IphSiQ/KSYWB8tP9mpUjQf0odNPkzIhjkAfwW2zBBaSDwLkbPNpYT8f5+xFuBVPV
0k5UT7Xx4DRSkY/VdWHiNd0BmLGENhhSeLWO1U8gRraUqrSlokSmCuT+BDjbn/G8
nFPUIwNnRe5i5eMG1cBSJTWECja6tdkxEeIljEmBB8HEnw4WT/aByaQlTOjPiYHm
W2DLFwnORLmpjbfOC2usISDJJms5qDGAD7YdGeO+ovsXaoBtrM0SQ1tlpSGHP28Z
hIdyO7v4xGZYnCM23kGTVi2LqUiV0vnHo/SP1fE67mYiFM6bmUWtl0KlM07sBRed
Xj7BWOLH8sH9+XrRjJvaeAolNt0G8LY05AR6WXmWu3LZN6hZPLhX8GsgsvZrwRul
vJcstI0uxGacY9e8bwNUAH1JQjuOtVxivsIQlAwowXIZpWqvukCG6yEpQXqCrK9J
ucvd8mP561r2s64SfbqjOitaCWIpRieaTfJDj0SNoot8/3/2LDVkuyRtKyErcjll
vfGpa4VhEsfpAxf4jsMuhZwCEtNE8+ifX2oDALTOKrkFeakd9oT2GC+dMPY7/HMq
Kuc02YyLxCiuI2eqZSGCi0PabFmAKgJEeY3vB4E7Pj9BWLSJP2ZVVHZ80xLkSD7Q
7rTxCuV2kxmxTMfAPxDycreP9qiDvRDVlR2KUP53lw4ra0wXM9hWlNucrrGArhQN
q5zgZ2XEVWhHZYFWiKCIaKzywWttJh5L0MH1GYM0QOTngJm41T0HRy2l2rzbiN8Y
njS/XebI502Osy3261IloiFGb6xSnfdwfsW0E42JzDrlicb8ZxPKKlXE5FCHdPtI
N1Tqov2HaL+HM/YfOmn/ADXFnBWHTF7e6vdyaMX0D5BTXD2FSSvYOApFLRbqA3sz
J0KWt2MPHqb8NIZsOiGZYE2iS43w8rjL39hLz0dPN9rSvHRYZ2SXTs6TxFO0K91Q
RrCHwrlhI1od0DSu4BBdD64ia0cVLY3UkgzrUZRbFWBCAam6P9BD4Qh8MgjgoT06
nK4wRMd7K2cEjD4qShCpfhib68FHjfxvz5mjDvhlpUXKQjULlUpg5lKn6qdmfYCd
Ayt6l0irUAWDbCk3uBeA+zWBo281NKhgSQBf9MJQ4DV3Z/PZdcCrSZJ06QU6Mzby
05lQqqT7lsaxrjujz33dJ7Qskbt+Ciik2it8D2np5wa/RB9tqVDAX91fezZJd9Qy
QX5qCDOv0qORULsk5SM1XGXQ99LmsVCdWmOLt3/kVnS5UMz2HTS06eTb42sVlATI
GpTs2ELQTCFlPTCzf49CBwJqTeBdhJYhUzlDKSZ1y3xCwWn03hToyxnnG2Iy6V8E
dBlzYhyS3v1ANC/4xnLg226Giwrd9HeAby2Kg2qXVqLRjmjeud0mqnvJwvHZ9SP7
ystk4/MEOKkxTFm4Gl02mVUGi+OXd9Uzm3vmjDrxs/Q+Avkfdnnh6t9TRq+L0X5P
j9SNDBGyNtEpSKXJmT1IKuK54vfQWpOEmnSyZyRFOVOzNeRvA9SkFGg8LmVrKMaX
cpzt1JJ4VFkFmJ3tV9bayCJ0HxW8UjSc96Z0mFM3VZq1m7r1UZbbpb8VUdmNAMsQ
byJjIxIXcgOeAnEeA/fF40jSb1Vf6de4ivwMk/H6+YM4KxjFFzIC3NMrEdYKbuEF
l0jtsY4LXB95vm2DUSVNQvIjVU0T+fx3cC0iiyr2VmFJ+JHG1RgIAEzPyTEcSmWd
Cfk2hIQEPlddKN1m8QNH1ZgwNjGk9k7s/tN+ZXbnSZs0vKK3ukfERddgLcqsMClG
y54sqrFCsVNKrlFXGM5YzPBTgWFvncH1UkzNdOsQy14yMjmc87mp8SC0grQT34DP
iqqw8kHjEkqvOf4JMHOSME++eufYyrgoZ7rWO7P2emKKzQBtU12iw5anZg9J/8rl
0NDdyO1DgG0iSgMvjyD9IgEjw4TdzFTHCFc5m2ffVPvVBbFqwMLLqGKZu267L31Y
7IdhzRpmWs5P2FmoQ+9+ZR5xZc5ABPpkW3wuI57t0jWHaU4Xu+aNTBM0pxfviZRR
ytegOeHzHjjYiAg7Z72zOrF4E4zvSdvulQvRRZxR36dZZY26gHCU+7BxINLctRZk
XtS1ykVV/QcmsNAkw4s1LOEou07TgG0bIop/6ABLRdcstSJZU6l4+pq1J0hmNGFt
PgSn5IWXyRSvHI3Fee0mYN4QZ0AMcEvk8UgjOKV8gY65y22MCwDnAABDsaRwMhZw
BA8IoC5BhhHq6JiBrjpkm1pOfRbv7THUvo/BBhAQQexx7IpR5OTVHB6NH58qzrk+
8zy070xo0FoVGHoaKdLZIZ7UAmYcrELP+JLOmHcrE6d9L3YvfWf+TA3/msTBY75D
VKFr0hNKcEnL5kjdvhc0itB+S8GmfqbEQXroT2tKashc2LphpPyXKGinajTz6+J8
vK3PXUGLGjIi5P2SgbJw64ng5AJU9UxqOJGg5xyYBrYHpsfjNXvs6nrSWk2Xl/hl
dPf5YvXwnizXjI0JlTNsCq0E3IxDn6zTr4vkpDzFomeLvecC/sDJQEGPrSiCVkz9
y+nqhydCPnYhoO9pseS7yihm86ML3ridi3kO8/pOGScR7Gxqjn+MrB6kAG2lHGyG
mbKRgRb6kisnVAmiPY0+LE2saIb0hP3Akbz48cb8iFRvUh/z5wo2+JAmIenmuOfN
SKoyyWZw39MSn2X3PkF0viIlfIOOF1hCrSGHpi16gdxUlSoxDKinPENvZvxbTO37
qucpk4gkJiTBXTa3lXBnDsCjr/Wdoj6ooGNoELHU0gS4mA/CabhUDTzaemZKam1G
vyBDwPkZkrF1z2kWAgFp4OhfFiPz1RPWmipOnJhIO08hJMeIUGeRUUE5/E0k7CpW
RuneFOLWJJLbU5frAkTiK8LM5/cBlvrKIsSf2ceR0jCmUPwep0Yj7sqpSI7DtJ8X
chHS3bPyrlmf37nPuyF4ZVK9XXjl1O9uHSPpYm4YIsGQ/Uzi/OyQzZBoBjpdH/QB
ALlGo4zyrJxdkg9qX3gMPhyFP7xmFTVsU6hyZ5dM0nC/SQVw5Gyb6W2tJvMXClwR
CopamNTXZYEvO2/SFsBidTVAawkBvAzRpZPlP+KFvC9SYy6mq2rITY8uBk6B+nx7
VMHTBGeFGXxDD4/zxnAvc7HNYBNFAayKxTXu+on6twvCTHUYWo8rR1k9+z9IPmLI
DhHIvb3kKeGz7xI/MNsT8sD2eQZ+A59Uen0/GvVmbmW4RX4+qlYWuohrCTWAnauL
Wck3U5PLMXr5Du0OLEVu10qYcrOYUOD4Sp6qbvcWn7unJgcv7rEgJNEmFCVwF5YW
Bm1nFg1ozfgB19CzVhp+fLYi30qAuO9TQfIFBeIa2u3783v/EGClnf+uwaD5reut
5K9AEwgqy+p++4+IgLLMJ/VrvawznwfVWglKjvli37U9HrQx44VKs3l1eA5C8gn0
New9CBGC1wUnh1MqYHe+ch2du3zFTiwZFv8f7SZLt63TiKtn3svMw5t7pAEvzHgv
4JCSPUyw8q9D5feAGHmBpgaj+zwk2J7h9nJhTWvDUG5m/nRONzpjB3in+NiIWvEE
2GlmJV3yk21Qeajd0QyBFdG7f4+AlQ6B94fD8OutEiSChP4ekJKti1GvIEzkIPCZ
kAWpYw8nawaSLSyoOyvSv2BxWo1QiyzN8ekt4IEppn8df6uAXM+iO1Wto2Dv3w8K
9IxyQ5IHDR/r+yQNvFfSbt4qfqD1zF4/N3+k3X7QEp+c4A6SmpBjTMUc3IT1AxBy
8MkSHCZsoWD42Rk9gYLrajX0MeFovjZ6OV5mWVUzKDR+gK78MO8Tm7vBQWWco8wg
rYzVuT0lGH9IzGY6TxLbKn+ReNU2QJ+lEvIq3y2r+r62WaxlWe6/EGzWfQkt3+48
M7SWDJxFuQF/8Dhdw8obQZyNoriJf+wmtmGpM/2gD8/udjPiBhoSClB2MoaUMQau
qHb/L0peaylw0/N/YcqL0x17qWrf34lDRobHxIrJR0+XRQYSjlEOqF1tLcYrMvrf
TEQZN0UtGKZuytIZe46NeERlF0/ZNX8ZUtEe/NpdzPqTRjbd9O5yYdzlO1IS4u9F
WfD3RTEox5QzaKaunKAihdTW1Ef1lXtHpehL/JeIOaTzfKXq452M07eKRS4HfRNb
qUZNHIev2wcWjBvmDyzxBxGPCz9cFoDCdX+d7wSU5CSJnSTc76V4MujLeA2Ul+tV
kpkFmOzwHI7xeJ6ww2SlXxFzv3lvuSFAcWZJ8HPU/eQfbe+FDvn/MEQX9qn280kV
+xN9IZ8IzmQgJw+gBFcQd2bNavg4NE4GO4yqdPK0S/ZPD9zk8iQYXxzshTWnofkf
p/IkrDuenSyX2Vm9YXYM2qJD0u8q+Lr8ySO7G4YHZ3ShrgtFM58dbWE+Wm5H33UB
8YMcg7fIe5AR/saKqqa3PYC7wjt6r0diD6aYVKgkgNqHkKo1I05wnv4yB3yioFrc
QhI5fYm3BKfjKwfX7wmxmoueHAl7kH30l8zc5B8yhEoU3EvtCWVOUbrZPDcsCxI/
mcsIvXV0KVaD3utnSn98lrqGad51RXR/Iuv6gFW+duHwPacwogdhcOBUofgleohJ
xAG/r4vt6F6O5GR7esdhu4HmpWFZL0zAsU3jefu5A5Gy5QiiHdxiVyGi6RUXzDoO
3ftMB7ADVBSsVXHlicC0xIdhU3zweRnzb/Oy7mfv+1wYUgQMplyrBDg/nDR44RWK
nK1LL+Kwwzk5jnMgK1QGSX1egBYeXrYLMcfF4enD6NRAlnC/bAAhgF1FGwSzNduO
ysnz6uhmioQy+qxCew6BsmygzMBDXS6X5LCWCjgjSyPD47UrO6dwK+b9Y2VYeXa2
p8/zox2XqEVgrxld+4Z2Y4D9cNe0v4KjZXGdvId25NVx8uax3ZxOUCduPbg2AeZM
FggJDuWhUA+E6pD8CHwuTr0poaRqSxKYCpGrXisvzPU9MCU1ep9/FKkHD2H286Fq
gKCs4qKVaSX3edPpys9thJSha5d76Q5tiYxDOIB9uDue1zDNd+rXu8Aj9IwyZaD0
v+p/y4hqB7wA3qdO3eS4s79r/ln4RY6PqOBbrKaKOkRf5XmVVZywl/+fkY9hqKmk
5v4LzglElS8Oaf4tgspZCJ6+NpPJzCzSej+u0ZbcSv8HqEGnaL79TDOzkAJEzYHz
CF0AFOVqyrHP3BIosedFm7wlFHHemWOIa+nS2FPX+Z0+H2MnJ8XzbNJ+T+eQ+sFr
6q63qoJ3il/mawdDcB9Shfd5rkHV+ZBHF46ONbe5kQ6fu37GXSeZBdYGTh74mGIK
u6Iu3HyS53+L6gEptCmYtBAwjSE9+L0jXQ3IiFRNNOBHFE1yEaEIpB5KkNnhTaK+
3fIxV/dQyToN9tWN0rBX6e6HMyqnh9CAnr1uKrmULVJrpvSOxCsYbqOD9HDXEgUv
9nAfdGl/PGeVAkPGrtmsYN5Ptw7d15zUoT7yreGxBaptBnSLW4gvNDmPuKXfWh7p
12DYG8p/CNnhFPdLcGKAVKCvNFpWWZwJQ52m7NwcUe565vo+hXIaOu5pbaLWzSNI
dU1GtC93n8wbb8wvilbfLe0aqvsJFe1X4zI79qGhcqb5v5xmWIIr0MSIbrtcaOzM
JRF4nEpWcXH0U0e38xA2YD5AxdPlyBDYqwDTbo4VyjObqN6F+tdaaSaLbFL3gq77
Sxw41iJBk+F3mjEeO8U6f7o3jlqxroyHMWPm7O1t/rJ986S7xef0yvc8U2hDf6Sm
CEg57ZPXXdeoT5bwjji9BNrINy2fBUg/cn6zrS65oNVXVpUq6kP7dFDRMUkgqCq9
vEKQZLgH7QOGiHXNqWUKDWtNMB5XDSnIoWwghIbDga0dyjD8Oh3RH5lsGFrpQJO8
k9cHAyG/qr0SmJJpSTJhf33FKKe6rnTrr2Hf76o0hYo3soo5REKuu5Xs5mzyaQBv
344m1Vjx/pfB+kIGCXhG/1WTi71pjNbwaP1z0mYtdfDmhjOAzUuD65qEBw8zpjc5
N94QtvbQXeFhFS/eZ/xmFjjlOkKWxarjW/tA7KNRnsH1v7DYwtSNnOCBDlGDN9pu
aYVPYKKMhOk+9n9t/22MdxQZP5FqNHjuTlQrdGosHYcZwdtTZCbH9xPKekRJB1sI
bhGEyRBbD1UVX7jV1o8e9TE/8Rlzm7ilhnuhzZ7JrmNZ72BEEivEwWrIwY7N81VO
FxT7cSgykXx8ZH7WIcDOPgJpqfZtHIpOHmBhjjP43vlBKacn6kFCH98hWLCBsHn9
NctBu4Yr2TpgQtvN2ETa+5eTnWg7xBfVqHGOdip2kl0AuNvcf3av8+rei9Cn5A1C
/CrJ8I3j2LccFm1D/BSwa7Vqvxh7gqPtuBGXEe2ZwCGMBIWj+jeAeY/sxX4sreBM
YYygShFVOsGOgj5Fve9Dd3e/PmMBsiVm8zR4wRGOtdXw1mV0y322Pr4XVQ3tmOou
/Efp0uciFLE0ZTmVEl534mUhqo1hQn+wNw4PCNhGgra3l5WqvyyvQIb2U+6QvwAD
lKAEXVrDYviURZStkJ7Gw08wL3a9Hz2itsG+sgstLmXX+foPKHPE6hEfWV2tXJIf
pOSctTkxa6E/rMwwmPoSA0BOg/+DC+XLoXGkVtDksxiyrTF3gycpZJdwPFdkUnfe
wNfGTN18XabvIS0AmawES4oG76xyxWNrobP8GpFky34H/fSxYVGj2njKIGCJOl0C
BvspI7c7MJZcguQ+gnJQVmgLG0dF8OifqDEf4z4TfKZwhClJiY7QNlH19bMU7h2h
HSMTtynufOGC8BQfoBhHWybtg4MjY+LZ7Kh6B+piuXLnk1xMDg0pvLn4TtRtK5MS
t+fCyKc9GkPabT9+G5UImq86IPed7iUbAOEg9m/zTPK3F2q/NlTqmf+QbvQKHsS7
L5p3mgUq3O57OPRO7YymuY0mO1KzHhOjG0e3xSiuGHOgAI2nhps0+sUlTzMVKFtn
Rzu1zl2D+tNjbrScKffRvukZfiGdGv4LnsU19E84KirGgVxlTcqe8GXMrvkRIWQY
5kmcr2ICHqU/VmhTyFvmsBJQzPmHmakGBKCOR6EuJR/2UEZptqJC+mK8m8fZRicz
4pl/esUjrutFFVf4NxbTi7qirp9mSEr3OB3hahCzRiK6tBlGH+A7YlDkHISNWpp8
A/qzCaJTvlwtRQJl8sKbQejZI4yODD0z5PcSVWZqTK8U6IRbExFDNopAcPXrv9Rm
qyhj8vj7x7WkFvrdeAXzlukJPSrwSAU/dm4dAtVDlu6RTx5zNY71qYX3vQdUQIvr
Z1UqsuWiaQOl1Ai6UcLrFjYo+Az11Z0ieOm2QoScqevQIdDhhRyNF4Jl737JbQO/
rR1xsWssonvoDcmDfnos7AGWRcIkL7G31mMXyq26q8SSZ0GIknVz9zfcgVII8K/j
W69pnf+5jtDYTVMqtkd6bFfXkINwnKtX6NiugTjBRvxaJu6yZtExLxP/R2h4Tbey
v74a1ULBis4h9TeFoWHbFRnsdWsku0z13IYGOpV/8+rOHrto/JJmbBCgIzpaLesc
qyxMwuai2EgeB6JzPECtNXCS7QXhoEp5YcIxTRw9AKVCXLeEyKMCHfmaKH9QvgjQ
KT7Lf+IXdL8HMB5wmFm/BFMSzyFASoS8+yBtZ5PnsEkD5O1s+FLQ6C5786ZmtC0+
e0oh4QD09fi9Fh4Pnml1N1VtEC9HOYuCCWCwJZD0kxMVDKhdZPd196GIuiL0EGbs
YWe288fk7ch03R+rUrT4V6CTmSsvMFcdClJaG5MGl8g3wUl4jHPf1R6/+jZMQEFJ
MxaAQdEabVik3QOADHYKJ1k8HzVq5tciTY7i2NtTMZG1I04d5APGSwxIqfMu8kRt
8P4BnFD76pBH5ddN7mtMlJZ2J66AnSm09vf8L4QPDWINq+Nszuwo8LaFRPmliE7V
VfQddtp6ZorlAlxQt7ZT6BSivEFMmv6H/AAs/tx651s/uK+YbEsgch6G4Ok048ZN
Ei8Jd/+CEa6xI+PrjCGGgLB0Ht4JKk3GZTM02DScrjSPshHdJoxPe2WUQv2GfVHw
9USk/XDtFhR6/Ehtw73RpjvHD4QdfVa6cPmV5TlEus6xCvaVrM7k3bLo1mfAB/PG
Y/1UqoAPNiCrUfUuj6+kFcU+m3Ew7L85mEBSyAMMaI8m2dE3JHbBwls+pWrNYALj
oSYTmS/EaPQuxq6XvSV+lLPxKMmDuR0t6r7y7ZbCYhGUOBcYlTIrsAg1XnI8g0c0
UwHfh9oCBRz5FwVpVCU3kY0zELYYBHen2WgsKaJ0YjVQA1qdv77HwvNDxRy8nxie
u/Xkwx0mQwJB21H0bgKjNTXvdWwzyhV/28OstdLe3SCqmQAn7SShLD6vMtPm9uGg
XABd+CF3gaI9E+6qkzbZUejEP33ZyMUSA5ybwsWFgDf7eoSIjHijjf4fH3WvBGu3
ZgQmu6ba9N3P3946R8q0leb21pWmRaQrG0mTDQJvrQIwYIIzd16/BapAYMUNhGtw
Mo6VeOgRzUIdw7ccihw3dabBZrgN6Nr4fpsOZgxiIri/11li7ISSVaD7vLDPAfHx
KsiA/mQIpbAsYdTEL00/KU4P1OgVqehti8WsL9DLyjA4N/hgHD4ILCwU3m6jw3vN
LP+TZGiUw+5Ab/6sf7kd0Hb2en8CbWZZi/XTL9QRi712/+g/bBU5WJNhScDP7WvE
tj/n8WsYFzzS0CosV4Jivp0TMgdNKZk9Slt36l7Vuh6SgvphWdLdFpKSieftuakZ
eQlXsxglO5/qshmqxpddtCr6h6ojCeuPTgFOrSTlsc6vYTDKaBY9OsXbaiUHmSmD
QX2YAl4tkUwvMrwxrmG6UERN85iGVfPsmr9sbbhSxMrtwHN4ouQ9Z/RUYrpDns7Z
eOqHTsIPfRT8v27+qzlCq/a1VgqMWOurlQ5OfhE8MzDn++B1ItJEanwVBW4KY/t+
YFFGylBXRE1YxD1wp8HSzxr4ldk/cxxi/lehYvEWzbNTAFsrmRI5MEk29RSwiJ6X
8wvkhwhCv8jQWITVSYiAUksgHBQXC0UpZoUprJ79/5KYXO4LJ4CKJ5P77l82zLZi
D6fq9c6QXz3x85XI9dIExm1kYM04/sdaLw80m/vBkyMRO6uQdi3QkqDvE5EfzPLR
bhUoR4tb3kAS8VsvI5p9tbrAafey65tBRbeHvmT5OtorGFymYtsNzFWWQM+vQ8uP
iYIlF7mB9so7c/jOi0nxGoEPRFVx7YPX+vGM9v2MB7MNY/QDfiLg/B44fC63VxCf
6TG2s3zGb9AqkeuKcn4xDivY1FG3w9HLoxcsIruK5kLDb7JU2TSd/L1Ktok1SjCo
ZZ+Hzv6kDdZWljJiL2CYgnN26eC6tWbOcZnd14GfZbAo3+jrdey7W/RAG+ZNmkPo
BqS35XcrYdFbTHGMYMeOse+kkxjhJleuC/HS2DcIXdujlqN2UGlWkokDY5wssYJ4
GwUr7jLxhB3ag2+hlZ/NYXyGqihaxvCl6goT4+kALeWSwz+w+T8zJ4QmL86ovxic
7Vq27V04WJhTBbYvWmFeN/ysp31dQ4YcBzGgaHPF+wkdzWMudc66JZIU+UOK7A0Y
5h2O8E4kuewlTudfx2OE0B6O+DWeifyzkNUIpHy0jXiMolHab8sIF/IN0QEyPZoD
k3JtpGGlyjIML7rYfS1dAk+MH263W1rW0o1cr90/H2a9lefcKbawmqPCywiV5W/v
uwvzLMaild98tXC+R3xG74rGkj0Ua/0vBLvrCR6JG/UZ/Ah1oCyxoIgSkKN7JMrW
pr3grALtHFLp0dcYYVewK9d7J5tSXNWmQbhWR2Y8N/xTynjzCezqxiqsvJsVKJki
9Q7Q3PMFxy/Ibubw8exQxm2UpTq8Bps2zDH3jAJy48Hk0MMfo0hyuAYM8yf3/ndc
2KgDhJXiTa4HLT/B9PmlV3kMKsU7rMyA86jVE0CiVVUGou/aveSNWkqDa6ji8cRT
k9THczLlJ3Z3RNi16xOzVpHkU2l9ba+wiRimQmGradOCdLZ4Zplv1kOAVJyTd0dg
0CHOEKi4+BVaFrNz0zMUqyb1R8ZDGmEeN7jNbNRyXtc5ol5FZQt4fRUjJdd2o/AQ
/ScHiX75lV1IQtxROxPXBCWTHOZNx7gmt97H29/uFEgKib6+5gwBpUkEOzquSJP4
GGALST4kJVLywYH2lJgo7X55qSy2rx+rs6HGX5x+r4g7yGLlyyKkqmsb5V6+rsoY
0LvIsh7a1HqPegQ17cH+1IWywzIQVpyc90FFXv3LgVLiNKcQa/ek5UHd4TpcIM2q
hoTGOAvMX1URNcasN6kIeWLFBsGU0Cyswn5IxQOZ5KH/3FrdlGfDKIwDMkjB6shF
EEZRmT3ReWxffwxKXvmBQXEOxTkN//yTZ4QAJj1ws5bj5L1R/oH2x+26+pZUjYY8
Wwxpq92W0YOkqXtvHqkQgcaMbIl2VVzxB6b6c/mmBzLCJ7hqXM+Plo8Pt+xBUWm2
RiXVEW9ZLwN7HIxT+LYhmHD8XI7BXZJElxxaNqo9P6fpTSFPyuHDkoOsS6zdMJW7
SrV4IXkldJuodkJa5Zry5Li2cViG2+iQMM0aRF4dvDo9pQ3gYRGq8ul6SfWM/SEf
8dzmNbI+2w/QHIPj1n55uc0klG6wKArG8gyBwdlyJED42sE4+HhHmk7vtGqZE84f
6GXREeEFkvYy8rr2UIyNlKSONWh+J9v6t4+AtPS+rk1F8RnyfW3GwRAH/uohM20x
uhSs5zI0UdwZQY9FLQQnVvvwnXXxbtOJ11qj3zdWVyccITU+eAyLP/7P94crf1db
KFIic43vs0Ud9d8iDFMUdpXmazTJ7mzg7x7X61nbBrRUWxO3P9Z7FGMbmXSK27KK
MB+CayzruTmzF2FrJ+9DWtz4RAjudC6sThG9vGMmFBoyj1aKykRS9XFsLDeWIVxZ
zZ6MVEt8ftxmYiyqORyoYP2dwMIfo6K/Ke7iOSSwte6OK5LgtGoc9386W1DnBfUW
emw2OWhE2laXaD88n0ZhD6EVhh+ElkbI1zhhXgW+EapRAsAv9NJCpQTmQuMJVbvN
sfVZjbYIqCcPLncwaGIVKe8tW8zOhC4z52phgM8dP4H5y2+HQWbx5LVNaNGEprVz
VDPAKicze/N82K8n59e1Mg9V8L4XBUypGvuKK83yFVCDg8FZaQopHRnK16Hiaqx4
dLRgsw13IhWdhrMK6qp8NiY9ySH+cvIiE9Lkm0UGrNBe407stOkPuqfwaMHdEjSD
O/0RBCBpZM9jCcuExRIU70ufmbJQ2R8hYhl3eHULaCxT0213AlMTrVrwOP8O6Dqp
VhWuJEscOmmMwz+Ecw8b+Kwi9MU9vZ4bWKUTxAs3701WVRjxTbbOBCS6VFbO/2OW
7CrAgRt5dOc2h2xXNWUWsIbSL8zeO1MJfmlWR1W2hG+XCr85qTVy5rqhq/ZFTavi
hcCP1vxIKuxmmMxKXK6XIdHM6ly0RPp3Cs/RrjvZIbb0wgoSd0599vNpOCP+4BAc
XmvVh/Peaesu1GpZHaOeG9Kx8mKf/fFW+OzAf6U0GlgrExbECQ2VuYjI+YZiznxs
cCLqfBxIoGOCDd1h25LKhFa5isoAnNiU3BP9a/OjRDYRxHMXd7EPOUUK63Oe1bm5
yDuTb1mUJ4tNAo7JkFimuYXh8Ydeax8V7G+1FEeSm8Za1W42KotO8HRAYC32B4Kc
fjylY/JP3zRqCEtO95YH0FinftuNkEJ778dbkxhskkz7qusvz+A5KlrpLeczC16b
rnNYngEx8a8bhIo5cM7znXC3ncHVWbD8ToC7GRVz8EvEtSHyVJrkvU/BQrBK+Ho8
oqYh6o6JmMZHnKTBwNjLQTN1ze3RpqEBypafYccb+R3RSYi/s4uGvzmAvfMBVQok
uJ8OzPM3u7rcqZy9VWuP05p19FpxJy7Qy7qQpo0kJgPLW0IUUVb67vqI1akh/OmE
i4ckTcBZeuoWC2Gw+9uEsJpf+kMnGLbAoLYt8e41+xZJHousBli55wjv60Sh1iKu
lx+A3qSx/5LKaeezCASkv2Go5KjX1mrupLMAB0L7RPguR81oUjA3bQN8jYbMG4MC
Jj4VsBQCZi3l4HX7eE8jc+ZjaeV8NDI1gGjK4xsvrb8IZpGZeKAz76FLj643aIaL
HLlRar5cd1flPo5nmvDwmQT0saeskQit1bgbSYglwPF27+hNPnj6OfxxfU0ch76Y
FsKtdwJGUepYYzuUe/oxEXV2ajHa1nZ7L9CgceOKPFcmWOWoOIE4O+um+g3bBZhq
geqzqrNvACOgTcaFj2KTm3kEh8OATQnyBQbDwT+9VKFUv3B1pZi80fjb4KIdyila
7uDeRkJoWuibKDMbrmNkIVclNEVsqZduIqJg8+iBQQw4XG4qtC88w0z+uiGme2tz
XPvLT+QcewSfgA+YsXEeEh+UCRkAMMPlAmv5DnnUmTcMm1P/NBDCtyr7jglqmOcK
wvBYJ49qA7Jbc7qj64THkAAjHr5hVggJ569CtbRoshSqppEc3c7+CbuJ/vFkYvct
FkfPXIgzhfevak8qSt815vE5Nh3bEk3HQmdv8HPH9aa8BxgrBfcwNRH3z+OrFrSE
tzI6X9SLcgzuK+ppoLaacc3+dQFFfDaeRdp6YRm/BBH/+v8EkSaLXNsNQgbvasm8
DRUP+vRGDCLVWeIG5P8KIlpIExPMcgrZ2pgoAwa3uqHULijzdrtiM+wffC+NOPYR
zwvzH2yZhbZJ+Y2+deDE3A1hNKARt+jbJKZbkKvpfN2wI9SP0Qtu9kffsZbOIV+c
aw60JdwbbjWicdwdKa93iSCXe2AH4OT4GLYzwRgscfZiHzNVt7KvMQnVnUuAgqOv
FKUyL1BLhpZzpEIwIafZAgkaYmejycbrwaQjOA2qg4dwCFT5WpWyCuvRrxTdNBKj
QrccEmdINtIHvqT2D4YWL4z1NMKRFwTZPCPmzjZpPrToZ5AU7IimELpAFkLzRxli
MI9FQgNC7iCFSiitAuZ67d5m3pcMhJcHHXANT6WvPtagfo8O/mOzCk/o5Opow8zG
gNmZhVlpAdNVy7F6FE6/PnABZmm+v7mve+qqc1D8z6huDvaaJprdQzsHj8LrLRr8
xRrwwT1d/tl6JVdlQPTxzO34OuQo95/rtTM61FrUlaNnttlJB92bSEvrm+ePesvA
FQhWUR4b1JrdZJTA9muFQfCLlLimxW6pZwShL5QQGHOLAtynsz/vhUbjre6WAwWA
lduI/NS3pMmESMYBjy5mf4B6Cj28cRj2M74ybE7mtsL1M6JbbtBCruxrKJl2rWj5
Sv9bbsXuHTG0uuiOHfBFbTFE72NKO7jKzd9mBcJ6q2hxUrtWhn/0smHVXHXFYM/7
UX42FhDBkb7WmtMlfNSaQD5sk0FOVJYlqlaqThmqv++dV1E5aliADkdctXX2w04u
oceE0jM+PVVOfy0JMjwEA6YdcGu2PVrvCiQtkX5xzGVT1aboEB0dkaD56/7AqRsa
/Uy/1WFmzeXldyCQOoKyIoFvnADUgJLmkn0qPBfct3qLyhKf9sGOdU3sOigtdrWV
pxn7NL3qAnVEGcTA9u7Jbl9WcvWBa4QOs0VGxRJNOZPdFw0gs66kAFnvaWpXPOaY
aYzsqIgm0TrYiHOsPto+S4bPX2TUEgt1nrDQOqPVGxs/lQ6SsUxv6gdrJ4WhXnue
Gc8Q+JLRRuKEDar9/ZNas764EhYDBOcv2ySyC94pA7PKTAJ+Dt1ci/zmXPj6WX+X
GpxQ1cPRIA0OBhAxvnrM7Dgz+IiLj03IM1ABScZPXgsB/IRjPS139XzMI7dczngE
9w6MSoJK1REZOQ83QayPxOX/2wHM4z+ifa53aw7QYa1ppJCEQizO9gStmkfpkD13
UeT4NaVuht+fKAyPA1EtsloXLJqoorTPdeWvJdXfUdTTX+blYx61R9cBWPjI6f95
2IKV3rgxlY4dw6oLcO1DPrVPWqP5Osg1rfbhX9vyvZ5U7h/QQc3uOY3U1X4sAMdU
flTnhXdPxUqVHtoaJT8ip6g89+3uMORPR49KoVa30Qp1wsktb3/S/E9OBLukqjPp
N1XM2BpRMApD/kKs4nV0RDgF2QSqledwq2nz37hCINxc4Lt4joWwjs+aEQ2j8YiW
GxveSoYXibpkG8XvBqwi0GYnbFjR6rptlS1o2koxUQdFIuhXO/gzSC4NUdGX28QG
tBbvjmUpzaAyqmWSMG9uiMdGBUDiqsE8xU1bULs27vDJ5VItAyb0ZKCNKxTp5oU7
jBHIh2IjANva1YglK+/Sv40Ra7jVL2vDLuqBkx74Ye4QfCtZfDu8h1/+u2ZY9MX9
9AxQCWN0JJsNPRGDtLB/tuwfP9kqENmyBT4l6gXf8PDO7Md9hqgVmHYXsZujKVFL
sfi39J8l8+KywYQklPzvoMXaVpNmPuj4n/Bb1zSH/znozYt1UZy332KjDt2tExeq
TucKjvnKxs2h+MGY+W1qOKcVzO2AzPlUxulfALfES6mU4q83nuitgBMXt998y0u+
CX15sj0xMRP/+qq8oGPH8gJkjizsrCbhzzkkXi1vX8qjjhFEEtNBDEtqCdCt7s1o
+KOaLyNzvm27LR93H+8hIgI3ZZ94JQnUIANO+ByyB/7XITNYr5cICDf4D9RzPKp/
ukME0RLQFG5KtuTgTB8MAJSwkFdqt51f5WL7TbeDCoYeWX5wHBkWCawEuVrX5m5B
1pJuMLvZ5QTuJPAF3ntuKW8K/QS++DZuov1qyEtMN/aDRAdODYbb6lSvlm2T8Tq0
1WnubLHR62x0T2BJQ0LblFjdqJKDqOhmMUbQg0mIS/c0eGdGiWvCPN/1Goq8q0Vg
sEQ95jK+dLf5HIfLtzzwm0El5IGSJHhJO9DmePpER4VoRu57tH4ybtawLF7Nndbs
`protect END_PROTECTED
