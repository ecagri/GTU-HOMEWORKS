`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1tZAlEUJcibwneDifEXO+VUBHlKrtw2epMPfy5usDEDAZkwVVGTL4PwfkKjSm1Eh
H5pFqLhP7m4gLn+jxBVv/KjhftbhN0WAWJlBBNpA/zUqPL7rDat77twRPfzicnfN
cIC1cTiFRieKJh99k4xL9I6YTf0ODmxsPPvldIUWA7nfppBbBag1LVvy/HqY6Hvd
i1kGhiIsg2Y7s3rVzLq8056zRwJ4mRRezXparchJSlyespTpyRxMzqEnL0obuazx
Ky9JFkriPZtKEG05qYb0QfRpPgOlByzk5oYpbYrgKY0HGNsms+dz7gFy7fHSG9UA
SY0QmOi9T3lnLzWl89YXSig/f2dNs+opCco1EINGeoa7Sj+U+59c1z5sKvuazI7z
NN3bNFjPjth56D872svJrVQyJmtP1iJRwJw/Mf5XqjHeaH+wOLUM+KHXKe1A5HP2
z9K4fpEh92F24rCkAz70ia4rNk6fIipbvtuww+3G86vjxUN/uYBX7l+MxoNC6EgR
viupyR8wCc0urtrXYqnpzAmrztSuym2lEWPSFlbMhMnvVas/8sUxB1gweY4F695w
Zg8ZPaQpIjgutnVbsAxs9+KfpshmZFX8nF8uKdDvqD4aTpxfKP8Ehnit0uDvvftQ
MhJ+++T6c04W5sTtg9MzwcGmWbge3BlYgKSFatNuM65j2gjbwmSWfB8zdermxRM/
LccZmr3CZDwJ6ZH87alLekVhZ0y/mW34Bee6tNMKyrY=
`protect END_PROTECTED
