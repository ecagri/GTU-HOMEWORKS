`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bCmni/BbXsulCCuJFJZBtRhUIYKg8vNyED10LvxkMQf5OmhpV4wxDnJ6QzZY8grY
ilcp4jhh48C7K4Lns4XrnSpg9j2OHC1VXGO1ebMkLkl1vGRpbgui1qRNswIFXHwa
Hds5iOh/JZXR82LrtbZ/dt30JwwCNISlawTmRYm+QvtfS/vhG2Z4uiH5WZ7WURYX
iZ3Q5c6d7eeGaCXEhxyD7ez8bCmgf9Ka1xHfVnGEzJKOkYw4IzPhBJw9dYjrRoL3
iXXcaDAb8V9FErR8lrl5EA4HSIFRs9pSL244gpRHTmm+lonjTGFaSaGIllAl2Iv/
YCt2tB+bqTIiXVaMjd8UB37lTyeMLhS0mCYbxqFBP9L2dF/NY9/itNvChwqDnGWT
flC5e4fc+ZzLCTCJ9mN+JzqBCCsmH5gH30Sr9hTyzkRqk3RSwdG6CLa6sj8+ejZJ
rwOJWzrrr7ODSOvmX4c2Y+r8Ke9jpG6jDiqkaa4vWQeJ3X1c9Clog5xOX0CGU6Rb
HQpGeYUcXUXStmbafF7gc6zTURGwm/2yvsSTTvXPtfR+t7PerffMkrXPFVC6V2ZU
OgRmNViDJy2iPt66nL/iAg==
`protect END_PROTECTED
