`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vgUYrPw1vsP07IJniHEkVcNVjypNwmMRAgFC21MlPEArc/uqdYSt5pRjQjLqDrO6
xwzo7cDDYrLX4ifYp/oHrg7TPfiTwuQAHa4KTUKdawZTJncxEDp1QvU7TgDSpdep
smdZeectblzOfZ7g76zFmBMsLJuq2psBeSGr+Il+TgM9EMgLrNHTRaXwhKI1BRJG
JoOfYxt858838nrHT0xj2dhn1iMJ0SYnCU/FSpQGWb5L9hjzQYPfJyBouVlE7B1A
x1Q7L8ROPHXtnA+StAcT5unD49d2z8xLyG647GVtES795I7suyUU4dg+pTbMx+ts
ojLJmJmh9+z/YZydDbmLij1qB8nzwVe0pGUP8QLu1IIMzcYUgc5kP2u1QoflFu+8
WZNRoba7NrQshWJovC7PMgs3/i3/EJmjwccZvGJU4iDGaQEzvdeQhpJkkMyX1ODU
bu/xoJk35lZC/b64Yyf78gm/xIHs8p9vEtbD3JegI6QKMX77XGIUVgEMJxDM3zgr
XQebgTV/Uka6/mRkEfe4sABAlq8Nq64sXverU1bqk92+14zqttmBFSBm4E9tYFXD
Qkcw4lLdq1vjYBKglGmfgC2I7b5e2mKjfugq8/HWFd3Ze0z7RDvwcXfFC5m1E70v
7Bb+AS/gU0oWXfampLsuwqP+MTSPuwk6PFLSVcoX0yg8Ei+AIzZ1CDf8euz/OuXB
3vbAou4/KnByUoPTVFpb805rt7JgCEH/+rgK3Y4lqYwlQthTif4vVJ1XGcDQg8YI
V+VDgYK8M1QH4s3vuQMn9gML7MrJbTWNuusv6uGJMeBRFQw9ooLrSkp0JYL3Ncbu
0N+CzqSAn89D3XFZKLMvC6P95TaNYV9PDJKM03/tHY1fFwwYwrRqu6dShIJ0KCgF
8H87ZPfoptoFU5T7Gpl8z4nWKHtQFs5HHjA9G0gjEROJ0vtmfgwvO2DfP6uaj69M
nYJy6nSiOU7H+mUQA+iosQFBIyhki8WULi8OIuE2MlNdPT46HrLZkVHjAxZiyqN5
4Hv7+fA94weWcLeD0HpPmFVzffUC9MeadodBefyx3lkIc7G1jZc1nnBaavqBxlGV
9va7FAv1hxtGTFztF2tABjjH960DphDmt4ICRI1ytmXcsQ3tvIf0D9xmLWKvX1Af
+Q9+SX1DM/7GVSoqsosP+sBhLWShd6a2KXaYTkSQyR9SMyeljjJbsuWZDlPCx95a
2FMoPZbILIW/qfE2jppHUuMHWCXKXwcEP3EFiRBvwW9jRmsCGg5X8/4kcN7vFKYT
z+Y4XqdT5Tjg6z12oryZukhTsyKvdSCczSbSTVAJpE4U+KWRtsPh2z2zfIqj/GOF
`protect END_PROTECTED
