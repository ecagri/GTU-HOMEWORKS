`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BZggIjTu9oDJcD7Zq6py+gRXiRMqxyiVPYzWyEv8BdfWZ3gzhLX3xUFvUWvLRy+L
X2BKOc88OllEE31ndxnGUh590vWQ3AZISbOacC46yoLdzCkpoq7ahMSHctV3c4+N
GOjnk4SL0C1sKdjKkVlcp33oMiIuD51zeNdzPRYQC+5ZG9d+CHaecsNRN8c1ytor
9JRZ2/rxaG/j6+BCXf2nc96MOApZxrRJdroSOByG1wofOGY999zgsDWTgmBDShJX
MtU2Mn8aP5gi8PqTJw3/7FtdoFkmZ/FCpWARbr1t4zV5n4r+8NmYcNjAfnKTja6j
FqEWGxc1a8ktZDmPY4y3GbZituoCxKC8+JZ68LS6DKsT1513B/vLJLzH+yjWOq4U
SDQ1yg3kjTm+95X5oG2c0g==
`protect END_PROTECTED
