`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AG4XXckIGmbrcTxTuL+FfGL5WjEExGiq5v1EL4W5rf9OnLlekumP2hdvHm9UA88L
EWbcGBuW5v4wIgPahwkVRgKj4cziP28u8rcWm3G9K5CAP4zleWhl/YdCdGVhxaXH
44bjMnVdExYQuYAL+NvuC1MATW0OCtWG6FBrj0mn4qgDkQe5T5o5+IufHu/JNt3M
+AzA7C74LQz0ci9T74LPjUcQaiYqsbV/xIpk8PvS99j0phqrpo2VkiFFdS1xBrT2
DXRa0Du/7Jnxu7E7aN15u+X/VlpR90IaMtuZGvWXkMxYG5wKKIxZXDSHgKa1BT09
Au1Auq1hmGtCXQqswrZrG6vrIxRdo0LK0Z87ClxKxPQ6sOCe8SrGHr/bNaKC03R/
egQ+2a8WRWia5RLI9cRsQ7ZGBqPD/Dfv6nyKHPo7+LIAO4hR6lyZ849fu+49y3Kb
iKvSktRooRg+/wextzyX+PpKpQV6Y7f4+di6z5lkxMtAXCjLWvEB2fOe1Cazef49
TZ5JKkrhx8JjyrPJLTWjbRaQNdepxOYBX/QmH1p+zJDLQFCikzJLwv4Sg92g2aHB
eZO9q+YnqJONgS1RAa3e3SqUJg3kpMKbMkxefLk1SoApVJd6kFumGHDBpMCwUEgg
pezfAFmVX9haA6hgjf0hVl+Td369xUzKm3IfdUeuV6mRUXQMKr0ROQQfyAl7w40R
5pP0Zr+So1ceRLzhp6Duzigvvi/P98Ah6jW9qCVVezXRTmJxSGTFNRBEa80ADr3E
idsmggHZqpHkiC9HMHL3/OyhgL0iG3w7iqADRVSuQzQoKxcuWn53sFopbBxoMZXb
LUAgCcX+gy7gegV4HeT8dPqbBGFF3lvsbNJNmQSRbpVFJPlFujksCG/RC+MXgDVJ
tu2K+DINysE9bTaXh8DR/8sadW1YoeBOymZyUp/MPMNdrA1Aht171AdXPaulBjW8
mHehKT+yBSvcHeN7kBjEpWUQokZIQmSMjR3TdPuyxjcmkW+sZUSm7YOsAueNYZpg
vVz6FDdnEqfdxxKyjlljoO2RPYdNiSJfS3wUrsOhRfYXqS0YC5n57cXEfy/fHXyu
po9TEm6NfXpxF0MVEsImTjR8eKysAS+iUpm3ha99gPHWTMG2dtFePCqxxjXM9Cxp
xVfhSIP7qq722tdy76INT2vE2bxh6jtt0aQVFu4ehqMUbOafEWoc1vPIETocEOqc
DJwzH6t7OGBxcpTV5UQ2voSp8OyCg8/apT7eDmlZLVlZhMFxIcyJCD7sjbZ28VLS
V7ox7W2uz+mu9KyzNy89LvNxSF5fNMGNapMIB1nCL0mPCU5K6Hn3KDigE/M3lAdO
6WJLTHjaE26ywI0f1V2DvktczfnPVvh9KiwUZireMUBpPumva4qLqJuxTbVggawI
Xj4DwX6vb6W4E20MN1ZcSmTg2e76zTkI3ODCp3vurYMof8yj4iAEmuYFdm4knGoM
CQHpjG37P74w/HxKhn8v4/GGBGegjJtoCTmCdO6Ecps8r0zRiO4GUGpnnnrawBO8
jLaVNvv+XbQy2/nIUNTjB2VypyOV3ly9lk6TD/AmA/GN5NNq125XX1wTotl8h1p8
fJiz+9X8Y6oQxC0KOP7Db8L5OV25FBFegs85ozyssaLlToHvUNdy9ZEBdEa2LTqZ
xFvmN4cHlbIRv2LFS/UqfWb3d7opCpQ3l5asa5TXLRyY8xOn7gxH049RjkkPJecb
5inZQeiWSHsRM1CuXCl3gI1nawAl4ZKq87PTd5qxEEFPsWhpHYtncryFvWsGMFzW
LZcej5guxHUMmiI9Fm959bmZ9GaHggHoIOy8oIqK0t46lwrh/60sKHKHNiITjyUT
YtIcaoxkybJToke5l5jSMV/XXSawZSuPCc2BAPIHDRnF0BOMsZ/6SYXc6XBrjWsT
6HycyaufZpXWZ1RKTE13X4jB4fdb1bmRYxtJzAatpi+zgWappTMxEj5NRJatTC2N
ZPLXLfiXKIQiOlgECGPmhkmYvzq6DWSUFSANgthjPILqq+PveaMWpyQ3d++3SmDb
r+hb8Mwy14xrfBGvzGInv6zKLnlcXixE7ud0rvAy2AlcCtYBa0oUZWjUou9kjUmS
g4jeor1caDfuN7onelHkObpDFkUyOpxZ88m81RFb/GwNapWnmejTgx7IX6PSVo8W
RSWnWsNNX5HigwvxdmNC+mbY5N8sgD5x0/ANIW4msq7s0O20AAAnjmGEVjh4DFJk
bsX+KFnvkES7pWcmMaCyLP6dGcYmSDOzs8EN9gfKhnYbol19QzBLamN/JbSMQZ3e
t8ubKhATfYfeejFL8cJhEqk1NUCSJj3822/NoajKv0eS/TrMRwfciamWyOcQc50Z
UHkZe1BJoSu1vvAfHp5FhsbH8/WmCNgE3AB2d2SAdd0rfFh/3hKYUGQPIzhoWKzY
x93+goQHrtkp/4a2pVr3Am95VPPnoXg2G/AYdS3ryb3hbAlsVX8DYSiJYkCdMFy+
uMfyPnhvSO9exN+YbnA5hzJmTVQICcVM3DsLQc1VA6Yqd99VEq84KJNb1TqhI789
cZDliDBcT75+qTnhOFnhDKhsE8gVHGQX3NatDUbcHfLDIJK3L1ozIav9EMrSMdPx
cwMRWRivxFsUWwl779F8cmDhzFEAxI/Yu+9Y3oyFimT+SJlA/eKZQFYtQFBSFU3N
XhiwnDbOE4QxgvvV69LPMybPhzQ6pphNt+dmtdU1PWd8ljGNucbaT/HbRos3XrA1
VEk7HiKZ6f8Vg8ktkSdcOsrXyfca2SzPnGlw2W8/vbfBcGnxrpwKBG1arvxDkyXU
mOvXngzg6WkMgMWojCHqNWLFQKMqtolkhJWGCGj+3VfVoFg7fvGxzyYpFnnKbP3J
oOLB0E6kOyrEevhpjeIc6dQIcrd2whc3m8nQP7+SDHZ1YR37BGwQFUMMe+WnRDyP
IxOEmrQlbHf8vR+atUOuoYPc9vQ+q1TvrzLXg5mgKWb2mdQFivkjTkLXIy/TtApB
MOycWdmr5h199YC4y1nggXfQnwDZWIOnuUssSZkB+Ffb3BF5P1LbaInW+HupM2db
1oxOrsE5e4Qb68rZ68TJ56GZNqyF7ZUgasQ5KzkTX3mDXEEP9av/qLmxEywkfPpB
z6ApmAc8ejSBWtI65IuSPtC1ZisGde0hXdqdxZKn21OxVBIRPfqOmKjsrxAWUXjV
xDJ0MZ2It1lt9PAyWJUNM0U2oseN95TKAJz8I+U4gkMCFCeld1sTgXvr3gtqfoDy
+rYHFswDuMpb7cXNFxH4N3fKUDl63SYRZN8f2USmdiIWtrrAiWVVZmbcPg8PMKNT
nalh789Z7WJbRAQWH9Nh/p6Qa+zNGdUw84eTORvfrjC3FaWpTliBZnNMmkhaSFJ2
El5hxdA1gCkVESAujAFei2QuE13XHxY6YuC3B1ZA16/t4jDBOcpEfvwrMlin8Xt2
RpoZjrvnIRz9zOEv76pho4K1UGocmHvluLNZFBZzBEnPZjyT6aL724urbo005PtQ
qCn4rfu1LtXW3CN+OwJf+PiTgoGlQ8/e9UnyEp7DZb+qEv/iMxzFAJCrCqplfc6N
lnd2lD/F0391AlSGJN8XtHSuMIZzlTpdTQpd9yh5F3YIiPz2EJ+eZgDU9twLumgC
2omuokwPMM965o/0zNyhlXBBxZDjirZxDDh+SdD0qYnM9J9SZ24/hup9PG7a3tAd
2vVn/uHbZf8UWaLrFLzcEe2rkaOgFzJIkIVApjsXv26V+chQGhkzux2rbISbMptG
0SOaMDx02YwpSDm9jRKCVqckO08LEHp0BQW6FtudmMiU9QSlNu3ciiZF6FlRdpQF
h1WkDUZPG84PWE6XQOig1i1ilw9iyfatg5r+oDINS9qB/82YC/QwWGMVsPLn7h4y
fqmW/+6Friq8X52XVTY/hIASR2d4Zo2YGZkJZ/RNqAS97QSZdd5hNH4JcxbXuWqS
B2dpycXOOcAn3nOpFrcFamHGAMRO2FnyztrkactADdBIxM1xRD92OSNBfLGhNimG
wmMM2xTCgTqbSdcgsENHspZWFp+2dOuMu4SilKh5H0pJia9ENQTWIxSob5vUMwUp
4n6T2XHzk/PyylEmzv/DBvUii7/xEfzNhYME01L+k9QIsO+wchOGEhBY47kZVsTZ
O8A5jbK1FP5Sj3exM/F2FOOOepRXiDp6rA91tNokrR+mX8wdDJM0l4ud/oMiSojx
jWHW9LlzkASXm35a6QdcsfsM7Bd4EHn1j54XxMa9kusHxG2mbailiHTfD2dLDOx7
+rf0GJtSrUjBUaQVYfVonC3BpVmMjukvwCKxuE62xBGjTJCNSrH4OUUWgATUZHJr
FNda65eyTQV8AWuhANMfXo01RN0v/SBnwnqWOiAtS2zYzyIQM02QX3ndnCMgl+pt
rJxruOsnLb+Vadg/sXkK8Vj40fRPY0TMG48DlWpU/oQjYPjRFIW0ETzpduaaRF1t
ELhJNfDfar7Pl0mg00f0F/TassseF69VNETVvhsKv9bjxX/mdfyjOZ7XddUSGv2G
lcOdRDQZZLpc/9xisNszNKrje8EpqGomYtxzYFfGw1yBiyPrg256sDoSWTaPvIjx
PTTd376Sl4uq6/9NYdZSNP0EZaDRPd8IyJyhHrKCXuLfw+Gi9L47Tgm9qA2PT3+o
2rEYeG4lBcrreRpYJTkyw92/3TjoLs65jtBEXQgt680IUqU2g4rOnam0xwkJid4d
wJivU2wSNLmsVQqJX6oPi8EjiVo8Tx2Cq65Aqz/u92WY4Na7mYTB7e3yjVn0c1L+
fTxZi9vAB34h1n2HgtA2JKm0fh+YB5NRdsH+BCdh7dPcy1+zTBGfOLmoO+HE336X
4BFyIEO08v7hwnl/lmlALdgmK3RoeZpei7Lxpm5hA0Fr7JuE7lDUFDnS/+zU5ASA
8Yr326Cr9Z6PoIGx/PdBLZHQDceQ9Vv5Oy0XBy77qFQfNgrH5iTvquhsGnd7ftdW
kzgy/ZtGu6+/+NMt2RGK5qt3nuGElbAvQYRPMHFQ0wGTs5LllVjde7njucSiRb1T
V1Q99jdRZUsogcoRpeNH++B2ZzJFJVzGeNhMOe6Mr+SNZ0UKRXVNRioQeQHn62+9
wMQC4qS9KBbe9IMNDnDD99kJpvnEhzTb6yGUnWA4+zKfdjwR0AASY214mh95QXWp
rv1G39mdQOCoOi6T8tmJ88LinWGRAM/MsSb6UMtacRG398a0NEzVletJkkQkrnON
Km2zL3VPANAcpzmONS4bRgg8iQjJ9Fsstcj2JVRFXCR1v2RdO5/dJ4xkeIRNGsvp
VzB22mtVdF9H5yuwaMpHRCL64emF0dWvIB5j0tTpMewmlKcFn3rarbAwhEgB9C0c
blNOSfEFDklTAHg7LlIMDvrvhbDt1V9LnumYQFmmEs8syem58WoutxrdtgUYj49b
oqYjfS3qYGfYuNTEhnhI1QHApDtg6z8h7ifoDptPbEqM+LLtT2EHOClaL0Vy6LOa
OXYd1dNe54SIUcrLmXrnEGbMPtLNZKZcrlfnLZbgtNH1kF9DujSvMlCZJpeanIrF
U8cv7VyEHSftMi9irHGPir9GH438i8l+yCnzB2y+8MEjQEdMeN3yauSRtdbqx3Xz
cogi0/eCsIMBf73Xo7qdFw3VlvC+ZrsKimBhYGQG3TT/HjAqpGho41SX4RmaXaW9
JqE17K3CJ2rSnL5utxIvkew0eiSFYL6WfVk+9sZ4h/Co8U6QFeaFJWNBZ44QRR1r
HUHpzx59a7BELT4GX110DVfJR9R0IUOjklfe7+sKTKs0ZQ/NzBwR5TCedNckjboZ
qiDeNBJbdbA+WQ5eP70+++nDMAFiFPlLvHUjxQZnwc4uw/sJhfUZmPhlclTbTf6P
4CiwX0jPKZF5QBvw1gPLdi/aYz2rhQC6NlWXuvVUgm5a4b+NcQ7YbfZcyqj6KE1J
JJqVTdhdCQwq8iTixCGAok25wa4MVkeSHDXM2Fyc6D24u59JAeCYpQR7UNGbxLs+
rHnTkLO3VWT5fJvXrRylt43Fxbi1mtiGur0rVziqoszaxrmhEOCTXwGuqsqLskxf
+cBzs/NholaWvSna3XyykXRMSPOgh9sfUnHGbUzAUiIeC6h50X9x6f0FEqJjM94W
C+JkAzT2xqGIjJj5gDmIYS+YrroRQa+TKiCLYkgumHnqFtc/Zp6Yd1+hmB2eA1JA
UVYSagOtIFaBt9+EA/JUgqfUMAORzMtJ7VkpeMTCEMa5x2Dg+k9v8DOJ/rR1iCbH
/OcGix4bisOMk5B3/Mo94f9l/aM/xUKB8IyWCMMolyQH7Yj+YWZOy6ENiJs35Ogo
CReiFT/p9ItQAPplxLJq8gCTJc2gA2BxHNUlfOnL/LoMADZSnBzj7GKN516namrK
x+c+HOrTBrGkCoBLz5t3OLU2kH6j+ov7uBMfZEtt0wWWn0E+zb5iXKiAUvDyqDaT
S1Sfhiaesj9jJnmKpGH3vMuqn03LQAU5iJsB1g/Ck8U9mJLSnIsbkD4Y/szchN3O
4mRbTWb73vPtRu2Z6UjaC50aO20SlbhgWrlVcplHqle2bwywhd7SMDAdI3tMRQmo
RSLsNHvXSb9SHbkSKJolmCDHRhFh1jHLF45b3Vumgcd4CZIiwpoohtJR0s3uQ6+2
yc2f5EIyXVh+viqjYQrVPHEKZy6UZ9ibi1qguG97f+oSGP0IEkI75tsWzafStL4N
5Xb9ytcK836r8Wm5QBx8LeYROn93WaG/PgS/Qk03A+P8DFORbLv2PgrP1zjNFfR8
dlHmLrdPJIzDHFsH78Jt0derwyZtgGU1jqef1r06gUbKQNmJ6MHCX4fUa0QHyI3j
EpwCmapp2Q+yKB7vaWl5JwyMDJ4/z85paCZo8xLux3VG2CYhZ6N614lSqawUp1N2
uXOOfaOOceVPvR70yDRYM+RQf53DoWt9Y1u8Fz8abKszogUFEAO2NJcyVkAzbz2V
sdmEfHudN+ICXRcILD4pib2KV2rhM7shJPub0XTCi6F73HIf8BPqrokubBbmhs1L
T52jVZUf0dDJbnf1pce7Bc2TttAVq2ctX/eE1f/74mN4sqGgykEcYshFEfS2QThm
h6L6Yxcu6fYs9zx3kT8pUVOhXvgBbIpbJwkUBor9g+0UID5npYOcrErkT42SSGuX
Hrqcc/sxlt9tUGR15+G9n+SXEtIllQ4yplTPA24J4QEZEG5gLVdF3FyiJj2OJzhL
txcwPijBZPSKx2YX5AfUa7Opdn+4cgAHaAO3cP605gEcNluP4eEFLZD5yTC8mCCx
zOwGt3aVEYKRMrm6qNeo45M5Djt/xt2j8AsUwIljvJmCVjfdo1E0vcnzA6wc3x2/
3HSPp8QSEXH837maHQUwnqYXh5+QB0o33PQuENQ2o4Jdu6+NgDBwxqiE5P1+b6mW
oEtFNuVXnyYOI+UpgWlBHgeppxjZBEqTmFxs3q8QGLFg9EsxHgCvS3TgBC1MSWKJ
7MYCFP4uX/ec/wtOggd0N4Ml2HnpgONOQyC1KGCSVbx68yjtsFJet9jTX25ZcCFR
JCva6KE+4Zf2PKQMZZypnQf4gwZ8o7orbvcWhcDhuZjG1W3yTcXbmwIzv68I1R7X
IMF8ZD3ucn1Eys2JDDmHfbnEFhPTQIUihISxS+dC9kd/263sizzPrIU0DT/mmKsK
2qxc6bZuB63pB5aSGWjWGZU740/SI7ev3cdV4LWHlFKk1dzU3qBTtLpJ9Q+Hj5XB
EVwrv4u8OKSVErqQv2L6YCRWvs7n8DguhrYQ2fyO1N3c62mpj3n4l6vqVGQBQ+OX
vgpaMW3XTOX5VUuFsACvz1UHA5V+IwrQI3fgNyRaL0+jabd0DVTE6nqkZ90Z2ZBF
SNSkb7metw6JqVfP0Zu8r38SBoyImr5401i8ohEazp58ogSmeui8gh/2Wp0S2YGN
/u0c9uDNlHnFeYQkPjq/dMEVTlgI7EeBQgIdmd7Wnpej7BB7WTaaM+Sw/rYJYHy6
tVd3t8AOZzVbuTcz3Kvi6yX3kfmmyKc9mxoMBU3Ktuem4DdE+lj7AXtBuKFf+6jP
pGfnGsX9XLlnPGvjkZg0ijttmzo+3nKkX6v1Wv4/t7Lmpc+MfQ8F3bBGt1+cMcri
vOr+Ogs62zmnuIkxVfQKE9WlFnh60ihKMy9PrD4Lo9DhgHRjwIKpBQ3sXdUPaHUN
hSn9msLqqyWxAwUjh7FBEGOyqRY8lzlWl4rXPMLqljboSnl+oYuD83Q74BtGtyof
GgD2DZJkxZiHZwA+K6zNUhj6nseKmaSYZohfSlBNMy4uk4pnjxLuhoqRlEyvkqYp
M1qAOkRhMn8TG2k8FVmq0+DQTfIMSKFxmMvqcHg+N9AgF10egYozg9hS4j6j1yqU
eLzWaRjaDNA8GCOc5IQSVyiEkeXrCdMpw07gXFuUYQ3ArkuUpxge7ZObGnmtR/cF
1u3LdVHYesc4IxhNoGL/3NVx61dg/SjVdzjtrrcWrVy+I9fbwHqlGmsn1tsRsv7a
oZs5C8Y/wtrdllOx1NyDJZyCPZ/DOFxQhR3ktz39tkm2xVJyMJDX12imEqwhAKNp
m8JVlJjdfzD9/C5eDdTE1pxzVT1pO8b8n8J0tHbvV3AiN0EWOX+NiMJiHinf1TN3
pxxVRo3r2JyVMbBOvg2etawe93PApFPHotSxPxKHOPQlj6Xjktt93HV2gjiFpZ9J
MkQJf/RuZ8p7kpmD8KfkWFCwtbVUKSSVP9w5u+5i7wdtTGaZ41VyHHPbL0mAq+KM
fJ3FWx2nDfS+mkcL4EUThpaaOZ0qRBPLLr/tLjACRfv6pYi61R3KzK+qkqBa+9dg
5XqBR8KkGWd2BDywCHBaUaaI0s3D8wzfuDNuoMzDMrJ05/cTzlALoeog02gRBvLa
jtt4Oy6Ys8MF3qG1efwXAzV8GxP9FdOmCj0OFK4jOl6QcoUGiai9riyMfmGAZ/tW
6ndHJexpxW6DfSQhlTCYuUpjgjMM1uexISYd74kaSjdedmpZkY6nTjCg9vKx3UrU
8AvGecNw1ZiPRo/CXs5J0tqWIbQhJMxMzE4Y7mDia0SVsle+hTqLpXnGL92I7Z6C
lN8kCk3BjUl1UQsKiSP+SKfvvbCMvan4m2uklAFAcIUF8f/uUXshY8BEu4kQTkqj
52M6Ir4rxeMP1P5DseosdZcYD2GkY/Ls7i0jojM7cYOaQ0RgX+zhUsrxQGVex0H2
fhESS0LuYSawvCNu3X6zbCYeozvSxHV0jDESRf+SgcPRzLXJY1oF4Og+to8xEtIf
pRcRTVdmF43CA+Mzak2J7FhwAIlrn3kSQVor/YRsFL/YM0DwnC+Q/3G2iRT8ftL0
L3eVhAbogRGca5YpKTR5Fek5H2TlCVSyf9jnuwmiJsNXlrJ8Hg5fvbSzn5fwlkPI
mX46i7qOgLUuNsLWxMT/jVloDo39M3cxQyEFzf+9hMbqD10I1s3DC8mp2Eqi/81b
Ej/TfgCwV2HELeewgmouS0exYGGkNUDtHzdTv6WnmMHrGUS03sS2SI92E/Hr5d+g
Sw8sVLL5qxPykNfVWAOYXXgrxsTKpayE6LuB/O5u0WIRPIRURAskzATYvJDExb0R
/zPHD68++lzEqPKSTPyULfVI/Mpf9FrCdvBe1sECxqR5rpfPogxJqNRF9/ZQYJbK
AB43xMcYPoUxOmntoQKv8+0MJFpVwqsbwyby+s0xo+bt1NtD0Vhsufyn6gvRBtRQ
hmF/G8r8dRwyx5M3ddKkxKbONkSXfm1G+9qiB9ZifrEKp53XiJEo72Zzik5zhLrP
dZDvjcpp7pdEvVp+xw9aDz4thNkcDwhzL3efc33m+4/NhhhhLghSc86SwSkxxrPj
zGzUFUP5YatsojexjeY8yagX0M7jmmYbq1m+/gn44akwr2urlQXEHAhQxVyZZBcd
/vUfGFwZHnKNuGWwZLhrbL1CbASvcLElTKnD4VnLPswDWiDjS21ql4relWXrfIWw
WXmAUXFya8PARgb53QbYDllwgPVG5/Fu3Gl3odrqb564Ly+Uyf+2/H6dduKcUiBZ
bIYvruqDtuye75vIuytO6OuuHfsaoXkyYysRt/G9KLxDh7+qa34ZI66TlYJBtHNu
HlTJANF0dj/7ZuOhwe8xf9Phi27rP4L19rB5G0uGozgBv7xycHWsZgzq2z2JuDPy
0uIUTMBd2NEVsKopO1ZTz/VPuA9omEzBRofT1i08HMUIgaomym4Rzv2FmHPBCneb
oKgWjbLJLwsGH5hb9Mvn0W50Qe/hT2Y2eNbIh0uBJ8pvi3ggrIlHh6bqRddavrfr
l5+zPCzj0rh+C3/3S76iQDQ70Dwlt4M7vQa2uGGKBvqVybLrpncdizBffPV/PhdM
hhxGcIu4BWScnAdlBZgpvDewMBIIQKF6FRp4Lbq20ORlOKKx15i2L99HORwzg9Ps
gyI2Or6fn5WUivp2rqbE2hv/r9HFz3bxebcEiHPJFYgnc7S/4wWgGgFYsOKGAHpj
in+i9tsTEDaaQwvftOMTXyLqYhKAzf9u7GHhTJKYqAWnLFXqsRH963JTCLancqeb
M6kOewelysDBx5i62Zuh3NiubQ20pTka5PLLTRrJr7JQswLLllWGRRZ7T9xTbyaa
wELkVoKe5cM8DdoDFaHbfwxI6646i9alqEZnzvqRXPWoDWwCjAwbm8il8aVD/Q4R
fFTes9YCPAIWX9fQrEfGRsBMFBSNyziPZl8TIOQ87AN0Kdm1QnBIUZqK1SNIMMhC
9N9cvCqQz+tzB8CiAvvAoTIONwjKRJIoz1K1Fz77TITHo52nIJWjOowH6Msa9uqi
gSaXD8FuI/d4ZOYBUh8cAJLPrAN8ALvUED5I/ZkzBsGaPQJFjS/3/1nKFyBS8At8
HxqoErOYFTMG/NamCYELHF347bveTUyhvDE/i6QGTxXRUoOa5nCaN4AxV7vqtlAx
4O9zIbkjP9cYAYfKT1uZQEhA+gE4sqIvK9bE68p7LXM7BBu/ATmGwD5oOc2LAfy3
DHQIGtLbgAegGGI2FAFsG/393ARkBqQL/x91s/l70+8ApA7ptN/QfZX3OdcBbJle
fVCizfW1zWDvHyNlx0Wc9SsALlCSSeSXeGcPyM0vF22pU5MDb5mVGpsyUEfPjhv0
8n/TP885wvvBq529gW2nWx6N9yvdP8UP+Myd7/lCQUfA6WP9cHQgMbOj7AxYyTiJ
NDCH2FV6eRCxR+OIehFrNdCVQdRbBhQPtt18E0+G7sBHluKI11UEonLO3nX4oK5Q
SbG0wNqv9Lo8VMPe42zk+EHUwYH7jpDlH8wU8ZgygGtIRrTFcUfU/KKGzDnNBBCE
HGeemVabPaI0omHw/e5FPFZgnCa3+wM8YqgVwaO3OwrBv6p5pxfFc+RJ+smSIwDx
+igwUh5XSVvrl4Nl8YEYc94PI9hiu+S+kG1RLiVb4bcK2rxJIJL16WhrzMAESjKD
rkz8UnA2Y/9gFnuHf00SQZBaUvoTIoDxvA21VF+30IouVNJ9FyZkoWr1J+en+XY+
jhhyHsFzBoEwzd0LHnV4fIMrQjWHIMbIibTd5KSpzg79jTSYVlvZ88nluEbdJ15Y
x5bvp2wYjAA7Tbtv0xoRLYH7aAwS8mgSULi1JV7LP9N865i9PrGaS1+54cD5NLY2
G4kfePiNfo5QXu/d1UVdXRLtbLmRinHmXahjPHggV/bN82mJV/Lzbe0j/E0XIb2U
x2g6ngW+2PCmDQ6Lo5SFYo7enG1gD1/xggnJ6QiVZjfuNEOVeP+0WY71u7teVa/5
L1g0sQ1ciYWNobHE4dm+K6LDUYCgsBezW9WNP6cVTUfQo41Bb0OSFX0fqyUfPMfD
JDU7WFiXAdvXzBckHiBukZOUJ5K0iatAZwhCIZAOOi444sLg5FWQyOXJ3Gs4o3NG
1tu2V/YEwvhTDYVVP8rHAarKPwF/+/G9k4QXE+f0W+O22Vxe9wNY6KbIuhEU0r6Q
YCpH5XvU9nliugw1DfKTnwnB1ZFXp7TC9cSfBfqnGOn/a1P0BAc9QRT4yB3c/yd+
tH9+rCz0YtzZTPsix5yFhV5GzrHGI+OwoA9S4tCQzcvM2kf5djVKfv0AmWDycQDH
LU4MbFpB05ludfZ5PX/tZDM2x0BgMiUjIVqnpLWnXJyKDrcOxCSp/t4kuyIOx0cd
h4JWvHvPJQpfND962ysKR5G453CHTj1IVjqDKNqHaRf9RUDZlumsi9OdbesKDZv+
39sHs5Pf6/6i2WRIuQ34xIYicxF/tJVlISXNgjF5T0o5RVNaQtmK5VImCHXPf1zt
b52RZW0XYdCa1TOT/L+DnFux09GAo4orqLtUoQqJHw+V0B+/ppinKQG6ggyQC313
GN5QNmjaGCMlBGXIG88G/s4e9sBxqmoRPOid4dqs3UGSbvujvXXMX6PJ7DLXRJmO
gTPO41o8IQXn56MglzzgWXPq1dek2+ExIkjbuYd9Bjh77448lE6XavKK+fO6KVSD
`protect END_PROTECTED
