`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YAqZtlnWDWyvvCp1earMAGbiFRT87t0CDX3EpyD9Hi94SeYdqpCbIW3e7DFotocx
wY369LkOGn6T5Omxa1boGGWS8KJPtj41/6SpJwVknkMhYOfsPWSJb9j9FAVltxwq
gxKk4XZmolTxv/r+rCN1hfBF/S8a+0Wk17LbbqXcg5af3NtpBLHO9IIRXwhOr03d
7u9e7WmVxCf7nZ5bKVl/+838ak2PSQg82ONgI3BKu7rw3ULuRYN5GeuHk1reMGuT
ZhCmPLa6VDogPhaQF6EScQQ3qq72M0W2bN90fdHahOQgAKfSSQaAQ/Y2X6POjpoH
8oz0CaaUxdUT1jMge+LL+ztx3tirX3je4keRLQxo3wBc82Kpq0rsH0OuqRvA6fhB
on4o0Z0U7w5PJYhFh7dmOIswhsX+S+ZYl6kyyHo6siqixvL7KgS+ekeuKFpaw/oQ
c9HCK78BfPNJn0pVoovDxeaw9JP4TMqv/m7bNp8MtnRrdADERVPgRq3TDOW/fueT
+JqVdeu2TG7omMFRkQl8atmnG60zEBGbfEYvdwUOJKgW9gK8nWybljSdmdElkoc6
1AxLB+yRULMMe8ItPL7RcOk0OCsj1AkXsOp/H3fBpYsXmFRjuhpuLmr5DGew6JrN
6LTgX2dT4ud/txgqwJnKB37j72/Ldu8Yn+McZIqDeU6h3mwcsLTKQDuXWmgt6YO8
huW2pbpxwGa/ZlWrKtYQd4kzGJv7u+GfcKvWENSmYeO1qZvyhX6bGI2W8z85GFm8
Ygz0BeZNu2XM0eAUmG/QcfCuRXTnCfObHQnUgrONJkT0cQSDznnjdwLCnya6NcNS
nTV0j4/szeTqfWuv8jDA+gFM1PulHAgkiqEQ1yDdavspcSUeG6hQp0q1WiPLTiRk
P8Or4x1qyacA8aRIRRtT2kK90EIGy+kOUHYwhldYcBE3jTnjfgUWnWna4YUAvPQi
M9gDmteJFdlnAIU3iI3+V8YquzPLF48Y9Z9WIcoaUdwYCOcwFipJsocHr+ZidJ7h
+6g3kV3LLR8MFambkc/JZXtDXkW7vO9xipxDS8nKOI3n8GJA7rWPCz6OwtEwoFMp
0583+bSEIe4EiSPxOhejtMLF1ei8zxJc07Kn30eDymgTuudzqMroHjowOsEBdPFr
ZJN3kTrr/isVCWfOLJDtdD35PBb6cdxhaNAAu7y1aJH4zrmBalAHZZK4EYLY+qD6
m+85GRU7F3hd0sX2CtnznLKuMyPu8Ca161PYt74pxpDXWmaRfpKB4zKIBs9O48LH
EFMK5f1Vfaq0PB/HVZrRRqQS/3oE0ntdkOeiJn4xk7V1OLGcQaXf1Yu513zPPqG8
jEj6KlsaTN2mLaVU7KJ2ww8+D5ugcFwNi+/h1GvYNwLZaa6m+WH3V/TIuYU0aO7/
Voj58x9PPsUQGJyk7WeiNAcASoqYMpTwpaGw8yOQYt8RuPJBPAz3VvnVXZbwTbLi
VWZbqnzZCnfZtwkvNI9VEgSbhTvQGmHHqEsTVzNe6ybNR9iOWTr5R3CWpFvi/XpQ
tU4pm/bOH1bmyn33wHy0rTyZiFQyChu6Iwhw56NZRVUGF05n/eIut58obST1FblN
RjAIT1g4ZcaKp4/hbrkrzDxr9QlqGFWZpXwIkq1P/3wVpvgMCLpAGB21hzF67s0B
DcEVFIVLAIHTWudkKBQCQ9A0FiTDG2GfboodLOG6329g+zS7cpjKZFYU4MsEo9lx
NjBXJXqlj04u/5QTiteih4TB9ryNFkDTS0bKaXfCpHwxgq6IUAr0SSzbMji42kA3
ghwFX4lb9qp9QIfNhFC5cf3zzL6Bdbl7rgAYQAGQdwdzadzTdm1seQLYbBMmi5LQ
5/sYusf9Ype2/5Dcx17NCHM9n5fMgd4iGGTaJ+dSKSgdTiR6LnrFIAP6YwxWA8YT
fWhBbdJh4EV4s4ColY5FETefAyzCgfpzDmRxMTkhv68ZXlW+LqbHP52+sAJm4uPF
1pdDEc7QQy8e2ufSStiSys3UmqcaKus3rmZWTY/bBCGiKdSpaQKjBdJ7VlVPoCpu
it9uVlH3QPeOpY5wSZPiL/yEYIb99e8oAdiFlW9IXLRbiENIEmivNTf+X6AkHsV1
ogkCj33kmJO4ayTqVan7W+fvg7nLEJxW2vwMG7Ch20d0nDDqSeRUjthBrs0kANqw
l1OllcpvreX8VFnStcsCvgqCZW0rRf7On2ch9ddDnBM/bGHcMdcegQPCPUeiaYlc
sbM3wS4kQg4zTjIKZmhnvqdQnehUhLlMNJROSr+H6TuXnr9KX5ZPMbqvMO+ARc6h
ORO5nC8I+8J8tHnciLsgzpvI2Va2Pxg7LWySHzXwZtpVGXhPJReMpda/8WDff7j1
gwfcgXwbwx1ycJGYipZeKX3RXGOhn1OeWQUujdcjFpbMJMehOIrK6i2Q2/+pLLIy
mwn0OinZtnuq45tpBVsHUw==
`protect END_PROTECTED
