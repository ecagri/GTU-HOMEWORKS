`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/bjXfQzd6fNwIsfPYmEo8XaH/airBs0TdOXl7WO2k6AGUFKGQ3+phgRBqCo0OeZg
5tpkNC636lp5XFwzRTT4+f8ugU9dBuarj7HbVvmLjGJUlSsOqBX0o4X6gk6RCPYy
bF/pxKFKmbXMOwy2xhYIBzszNGLjCnCRVMFQVdR0Kz3SKoZMBUf4snA/2ce6z/mc
TApJ4j1O1YFzT4yRPQ4VuIO3iGZHGVQH4pglzOje5eiwMYFvkO46ryKdVfmVbFTE
VPHIVBsmkkt29vN2BBAh71dSx165GxGT8WD1h3r6Zcwc8SfMJtHJmADhkt7rm7in
Fbg9L5dMu0AoG3mrlkVYEJ2bbpcWdfmieu9PV4a67AAWxoqJdDJkx52MNOlbn8OY
3ThO7pyzCAwJewUeWhefIsztFjAoV5JjtpOM0aoEnHiEbBh33r23TDqcYLBSQUSW
DJ6T4CVmm9UvDIdCDcUdBnkgBLMUA/QMMEOF3ggGYPYTl+RRWMM+jBxxHvaaHods
Wb+u5nHN6w+lI22Fr9gYg87KP7LCq9Ftz44T5My/UdA=
`protect END_PROTECTED
