`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qT9MWP9TJT3B4xawvc09oBXRECrveiXE+p9HUy+piKuDTjbjmtBbh2ukPcE5z0Ip
u9mzk+bFRSn40oToMy2xRCTftnN9KERm3EABpW0tS0WGOmk6z8Pk/jkMvqO69DMA
3CyTzXtOKQTi4bWeQiX5TALwKiXUXdiJXRBi+j6xUWs5AOxX3qmCiEWfSRnLlYpA
RKzbHfleA2mrVZg3TMkFAq/gLrGXlcB5fK+YHzkDoioiKAkdDMhpDc12zUMLeN+t
1RyfuMfM0J3Kq8F+6LqQjdskeZtbh+ToGBzuBmPzB+2u0ikqaOI0RkSZdCwMKW8h
dYISIl+xsrUK1S5MbuifZMKt3kKIj48D997O+t8vezS7g+1rLB3AYCFDKg1q78Vx
RtRa/aT9uDiXTIohhdUN64XwXTkBKZUggCBi1BayxAfD+0EJWgcUbMRtWXeQOvvf
l8tkgfkcWb8FaZwqxbhIdIKtFUcoY3E1mTIduPmPvVbZupUp/j51TcFJq29lLKXm
lHvRXKfEnv2LZKS+pORu3mhwJOyVbDij2508VooH2PAyKZOaqcH+YdzNiXuEDhNN
dQ+Qq3KQIoSk8gXE9EPR+lmKSMUpOL3NN0GXYxycmOc9Tbxs/ypUXe9tbGmTnkgN
jNfxpcoq92gwWJC4uPR0ma6BN1c1n2fuh0KpEqgaVP69anY3Kv6RQ6VxS1IzRVj7
Gi8CUbboh/Paz89ZSCBHcFHkLr3K1Rxpo9rdZsAFDDpCu5F26kh189iwuNkGTDvD
t7/hdPlrULPY2c2U+B4/e4aUoGoT9bwzT8zA5cYshauEWr16VleSb0Vzao5UnaZd
V/vtCQE36akkOW71cDjji+wTR5IDHR0TDCQSENHNkV4lTdSiYdkm0jLrJw89rFab
9DVilWBuZl17Sh0sV7dfE/bmLYoLIccH6xrUP2bY34nA2+uylnDmewI/JNJRD8p6
`protect END_PROTECTED
