`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yP0Ic+hSOwPY3QY7j7hCbUfT3tOGU0zNomUZoCIfeHCDSZu40kbRDuk96YgxQGPk
FF3zJdDGZGZrsw+fVsWnqHmPV7j4U4DlOh7vjHL9QIl/GVkRiLCxIhIgeUr6scYX
nhA76Dj+qYaVq+Ey1EGKeNAWhduqqT2lVNIvUjtiNFnhpcLtMzlVwI2qZmfH0w0e
gIVjQlYNfOLyyOupwjjK3jiVcRYQH+oJhuggQcjTEnCwezlSMoqugIk6a/w+lIx7
zMJeuujTe3coC6UXXkL6hwpqXjeMWI+fvwIh/stQVormJZLNGPW7hmQC7pjdFwTT
91JkfJZDcW8vmd0VdF1BEyc7ZouXb7DjEaLgPf8xdU23eqImRWcAqu8IfhtJj4qF
kJOUqJz/G5aCEPu9w3edp9KIYBXiCWxI+Z5jNmWmY/UbpcaqkWpzYKLG/f0bFRep
3JLSxuOHFYrYdTJmV+j1vJft+CRrAizY/F382DrloJsez/kY7bjPoC6vv+h9+O5U
rmYzqblRkJG7h54xwECI2Bq7eoEz+wu3FQkOhX1ruI3PiRDJprx12txwwBAigwbu
ToM8asF6rlf8thlY7HF4UIH1oPIoVpOX+ftXRFO+ycbTFgD2nSVixMhx79S9wgIA
v56ky5etyar/OlFIYGY/yUP68tM52EpU431GPcX2WzSjfKZ2lQCPTXFqOcEVUdn1
yQgGhkZyvRJsO8P/4VMoCRiN9gb6vARK36P/ZmAZ++8b2agaMr/grrE63o9cgU6L
wp1K7coHg8NqX+eWKW5fxUt1lc9fPTqKoZOnPaIgyexIGG0HmLReojwARiwgLxz6
c5508sh1K6Lo6H19vwdqpZTzyEwHI5ySpcfDOO909+MioP6bbwESlQVLiyKCAvuB
1kfGW4XdLOzMfZdXLHoqhf5xAICNLXHt3T2O0ADmdOZLVJOr9ZreEr8dS+d29GNt
GRs2iygPTETgIJe12dLYfWBduAD9wD8ecmUwqoUjBRl5QWcVoDDDH0jtU8cvDOfY
ZWbSoGal07lCRZrtmZloHNgNrD2pwUyTFDMJGifiOXl4j6wjbIL86wHif5nnXI11
+BTaN2C+d45LwM7lqXOxm7nuTEqWkWy0GnXTx53MYIQdrQfo+kaq6/J5F1agjgdt
TDjmeQYWBZU5etkZfmmL437QSaNaPZTnd+E6cZwb50L4WvgzBPmFv7IozjLn2B0t
CRIXNVbqMoUZrVjv8tOCgTnlEmfKmbLG+ZaCS3JoSiFl4VK/bqpqiZnAPlNFU4Sp
RWI6zAdUjrfO43tDOgU5yawyr2pqKAhQe/U5tlyOqKmy1ZpOgSYkfhn15GhUND9t
eT8/6QBpd+QkzjYOo0R9lKhUatJ7Sxcal/A+ABuwT4KHyaAhQooZH4Wmwc1pPwPA
qzCkTvLPWaUlQr+OhaUKlxa2j1qsOwauiBmfrE24VFxJ4yRXg46E3ZwCbZ6o8TtM
+oMGppI+bwNCODJ5tkoSYM7Wq5t+epgoMPXsvvpOx+IEJo202yqyiVazyyTnYd8V
dzlfcatJttdlMsB3p4zj2m2RsxbDYI5oLFhPrm4/qwQqzjzDjS0VM0wqFqbC7Qui
vmIPzCJER+ChZLR2h6oBgQpr8XfFGSts9BLevnmdrqtyesZKnJGu1EJFhXflAOOU
MpSKLX06VK5xmbIN1REbdxXzzhHLdZJWqkBc06y3OXp+u9iB0vSk5FYIxfCnk0Ib
12kxz8/Nhb7XFfaC6i60IjedENhrcaZSaxf23RdW6adCQ4LmAZpwz85shvl5yH2h
LiqB3vOFgNi/I/1utyxWvwb7W6+Gnyq9gR69uK6K1TDs7/Hic1GIKuAjWa3yuGCk
JfssLIgdyYRWakvZHb1PUQ+Tzjn4cDJh1/I6iTKlGQ9hbqlcMTEjcrpZbvr8CD/l
rdeMq6O7xHSE7sm/ecb2G4X/3sPiM+t2X7YKFm23C1dAgKRUxNYxPt5lYbHPfUDB
pzcIQP63GTEQzF2U7i9P88TWpdo3dz15ITuhi36UoS5+szOXHr7hZK/MMMQPwonw
cNQ9NpWT19qcihrtwqTG1g==
`protect END_PROTECTED
