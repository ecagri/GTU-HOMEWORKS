`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LXvGS1edbbg0q8//3TXazELSn+hMtCLO0Cb8nCYL1pet0ts9cjGvOLtxhKpyIyah
9crfyMKDQTfIu/XEarLbesZzNfwJyyXpBBWslTeUhya/DeZdsD14wsEn2qZtUzq8
LKolPFVTz4YcMpMmQd1TkP+XB691+k4uXm4cKM6o/JaROaWW8Itqkw5VMVhHo45Q
TdEkUrvBRTHH1CY5DVhEYM2kyGV+MYciQCVjESq5lNvdR7kPL5YTAa+6RSecCDhu
IfLOgsxsJSlzo1V4naw7PJr+6R+6WSkg6STCUNZ1hl8KnNU+1s5tR8wj49l6iz96
4LYi43/ifrpknru3bPyjSUHnuZKzYlH6hO0rjUQWQ9vm5tUzdxmWzlY6WcQoJ5oL
E1FdrGhMcyWg9PDFmWN6n4OZ8Gc6lGgBwpIYZoVq6U3K80PQ/pH3VAeKCHWdzopC
/o2AUdJABW1zzCZZ3fZLgYR3jnMUyPlZ8mfONp2ykzFXMpncrd4Qml1kEt5QqbMw
qjAeQ/X01fHGv+fXGRcdhP72tnXsAlebMinbNz1WP4ulrlZbVoK3q7QAk5wMpzf6
EfpT1Sugk6vBwajSJS4G5dDH4JotbV5TYHUdkTRSQnpEIMivRDwgQq9P5IJemUOG
MjF5XFBEN1dNpAJyahrr1jA4p4xZqKiVIjIEv3PlUKYYhrwhDA3KzlWeRX+oFXB6
Y20b/Cv6Q45Jqwb/Dq2N4MX9rmG5Dm0qVnh2dsJ8s6lifxsqaIWTkUUx295WFpXn
fSOqPe2GwDWjOmeArthj1vd1hdKx8EfrHzGvNW4O1lWq14lysso+wvY899j0kLr6
H5rztZvgxH1js4GmkCKKMQGAJ48i4niaJf1AXf+xxCajJxYrpT15Km7hl7NJhWJx
PUgkiK6ZYh3nGjfdBaavSoBKObzQvuIg10Dyd86w4guUR5zjW+Lef83zdO+ic1tT
BK8hF36y29xxBD9xHdzmeXXBBZoLxGgWxMXDKrIMDV0gTa2x7ZHJI1izavJTnT2S
nvf7KMmueKdpKjXThd00QCj/ZBydjOiNvzkw0Ar7z8QoY3tGYiVxrsIMZqlbNcuM
qFx2oKhwgTxoUZ/5fz4YnQ==
`protect END_PROTECTED
