`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xo0SmuGrM6c8fi2tF931PRyQwbXfYsC+arrLOPea8X4oKQWkpi5gjjf+Fu+YFW5p
/r2wwdO7QtRWv2EHd8s3DOdw6B2rnM+Pyy480IttuGbjFsp/0P7Uo53V6jQ/hvMB
vOjXqk2IjDuza1hrCwrZtWD3f7IQnafGOCS8K1C6UmoQAGjQzAoCQM0j0gzqAL5c
gl5ReHc1ElDd9rt9oNnjgB0Qhze5/pd8FaZtTUXuZW3mAdrRpoXZzf1JSmDduZjb
rI8tzOj+gmpqKLGT0uSVqnZQ4gk9ecRgQkkN2FhRGVzSsCMogsVvEmqOsfwxBgdj
0e8DIndlwGG8ptmlLUquMGUL+9UZaK8jSBbAiXcwv8RONadItaoyaYrkZ6POJR4E
rGW0+fATlrXugZnm25b+I2bvmBmrv1/crWJjtwokOPKOnBeVNXx/IsoJZD6Nl9Xt
Hs8eG5kMGFz/kDIb+bO28gc4OgoGJZzUFpXvs7on3VuyThdfVx6LoSeZ/ET/UOlE
yHReoY0tvxYnDpWzFl0m0AHob3NJGqgC3cjUEe3cerQR2PS11BwRtIQlCOTwEHV8
dO7lbpraE3Uv1TdAn78gwk73YfDjgcA7uOtplMn/bHBUilgrELxJ2/1+XwJn6TzS
adhNuHZuagN4oF5Vr9Ij2cpc9CChBvGhWyXqpiN4p3lGhJgB1hwT7AUcfmOQ8R6J
Ju8DqWYeqbEJIwTdLAOSlSEa4NxydLWsd22Vk4Hm2a7VLV1LmvQZCidR6vu6z/fz
ePN0xKnm9K53tGFmWc8ITqOABZmBJPvbaTG3v8RFfYgPAT0mbWMufhUavHnetsjS
`protect END_PROTECTED
