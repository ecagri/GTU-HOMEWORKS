`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CDMeoKk/Tv+k+XSlOlLJE8JKo0ziWEa1ZKqg+y1c8livhzIIcoMwRpuRUxEgoeYC
0KN7IVu1VqjbewkRneJn1PV5MciOPYbXuPyMnEF6i+oKIzAe2YTNJSM+y8jGXCfv
9icXOcDxFym9T/YIacK7ZPPedTIPgyIt/vvQra4Ofeb694O7QPX1062+goHSMOHI
r+wwcf00F51qmA23MYtxzPvFTABlQYVIbs2PDZHd/eq82dYbG79ZVhqWckTItWBa
P55XAQm66UaVa+Ol/PKZhUPEOl9KdGoQB4T0GAYvFXIiZsMnbsFVnfQ+pEqndcHS
utfZYRIJoGWyUEbXw374na2JiseuYWuJQlVIC/m9FtrRafeEM9TYvEPE6FR+psRf
`protect END_PROTECTED
