`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vF9OoWlm4dnbu7V85wbL508mJdQg6cOzciGJSMSJp6II6ZwkgGq2WqJFc0SAsFH6
kvu8hlB5b3BFkz+jExqtKbiY4L0ZeJDymnYDavcnRh5UbulMt0YnLHy/UYQl/3EO
FG0jZUi8YpNXdggQJJzYAY6s+dzMvvEm7VaZyYzKISz/qo9oQDJ9wKfij4wK4ILV
83QrEgaPAGKwfIv4vIdUEWMQD/M/LI9zXwFWNrttvHTmPfqRKzYt329q3TsZJ7B9
sPiknm8kXhC95GQ3Qb+CTg/5OqRYmrWvDihkIwASOkdVijh+Sga294GqBR85XOiD
8iJ7gCjxM9m7fT1q1DuaXhw/ISe91Sqdfal8A29PmQf3GzgOM7ltiXWxuBvvz4yj
rU7jbXribQpeR21coT6ZRwkactOVMFFeT1+maExU0poC371i68mO7h9AgT8cwqB7
EJacecAemyMIvKhbL46kheAIbH0uVCpgerjSctDSqAotPhUOV/XC6jkp95yQM5wN
m6nzrxMFn3h6WseLrJtJz68lAOQ3K8hVgJ3t+myOsec2S0n9x3fun7TS12pd2MUx
ZcbROj1cCfFk+GOr1N9Qv8VomFgwO1lPG9mRcHP441EzuyL0j7E8IeFL3+vWladx
iPbzArWSo0p3lQ9amDaFZlkXx3ABrHRUXyf04hARA37a2MFNpp48He9OJ1ToB6Wm
XpmoESKjwS+n9VVyUO3GohDRZN0PmDUylYPxEtG13C0sPC6WzuAxFCXMefmLPF5d
GGPCqDUTG2Nz8TUaQcNgYpsvGHDO4c30d/P5ThI2PDL1S6bSXkJQgrfdNhsogUZQ
rNQac6tpV2lGFZKEKEsd5hvePnHElBA9r86+55S7DHgEI8z5z1MA6o2++7fka184
ZP+o0o78YslBhIwlgD44IV4jURFbC7q3YBj1V8esooird1Uh5OqSokDYdZPV4nSB
7cyPz4KubfFMq4+kDQak6HICor3OZNYjh+nuNsTVkNb78YUH2ChI8NYuqFdxdieM
phbBwWeHj04vHVgdB85oI/8FzQQR6VIvUgcKP+8JpCehY8GoSjgKS1zsg/6tGPAk
6ddsZKadtPTTQhkjNSZOey0oZ9NRl8kD/pB2ZnLwPwJYKg/4o34zPsBHJw+3lxgt
B1cx1Kwgi2Svmwg2qLeH295HjZTTNlDdZ9v0JWxjNHf9GP2vmBxGxh2lAonbNmGo
4mVF5Gb8tTei4Dhur+7jPo05/BJTgzjXFBWrCNM479xofoSueo9i4Dhfu0ibfSzN
QnDkATbBouNqP7LWa03SwTe6Ls8+L1NEY4MlDM3W3Bpq1aWxuRTXhJrM8LjwGH0J
wsQ4L+hWqFJMScwVQ8OTmEL9dEeMxHkBYexbI+3tsPE0ifbX0kmk8MOQeDyzhVJi
YmdAiP6RdIQr5WwhwSb9ioZhGdOg7YVz4XsJTKwfcmIOWt0mMUDuHA5O5PI/ZzEv
DSrQr6knQpilAIGyZxSm9zkqnOPPF1Hzta7wELxIDFAFhnqpqpzuiWvipinJX9q4
PKcDGHlC6cb4yjtaEP+l4VSINEr0GNVnEG5vitjMei3hL85HJl9SAOAJWoAo5Hsd
BTztZVb4sKvR7PWKyyaaxMPX2S0sX53WlF7P65g/k0ENTFif2zkujwx8xQEZFRga
RtUuDscDjOMbyhdidyZJ3QHjXekBUCQsTrkEQtK/PRclqfycVZTdRxNXV4A3dZeb
ybe+UdcnqEd8kOi5GpHxP080YRVmRxvV3TGEfRi6whL9ks1gva3gzJYSu419h1fX
Tij2FskVkiCsLA50bFqPVZRxyMSj1QSu1/214gtrgIhkpZ8UBqRkq3XnBf1Wk4KJ
/v/lLyfXPiZdn6YAXchP5kUDZ6WXR88oKQfzEeGb4i1RENgMA8mvvxJ6GgHrMl7G
QC4/8VJPyj8JVkQPtxF9V35MZma361aj2k901/dnx18mfajHVLnjdn4qm8NamE8e
nKuPPoPr/PBbA4hx8LK8WzWeZe7gLxnaEsEQNc0KY8MwOCAMPnMUiAGKQEEiwvHM
qiS6uiSWUB0U3keXXPHnGHGyY5Uqd2F/hv7Gn5YfG23FswL4MiRlG4eA9YAO4B+0
0tCnYVIvIGB2XbsKnTtmSF8YzhxrHshHuV5mRMexDkl2HZL1A4XqRuA+k21/bw8/
ZJi7TRwyxgqjgayuJfwsmBiqRrb5WMO3tkubz+lsV4e56GnY74k0K+YH9iTGJudl
DtTnvCuNyjBZ0Q8rJsvr4QFJDMwTMJMM/U6i5VyfysW6W9Xp0MB3ZXUaLHPBy2Ip
x9xA6oqaAHrHhGrnW0NQWGsqjiGD1MSfNSeqdL1/uq5Hw9bwKsLDqrEdY6Y8fq9n
vgnFIUWv9IzquyUf2bQ+lyJ+ulDScY2hDUBAZUmD/68AOfaI+mVJPmYRcHP6dWtT
vsb29A1rY0LGlAKpKPMiO2Ox5MwdEpSgQ0dO2sG38+C9UVkhihWg3gMztHb5gdxd
N18QJUKcckbc5H7nC9ndWY0rS8QzBIGSGp2UYdJX+bMfCxdvy29vMkrVptMBK6SW
rmGl/37D+i3scXBsG1NRuuRu0cJP8q8pMFGAOCCujLSCR154V8Glc4n8N2wYoZaa
0um6S5pwM9Zv18xIcXD8oXNNgD27nCxasEp4vNfZJeW32lv5RnnBFxL+r7ISoAdq
YMX1llCm5ES6j4ODXs3rrDO4w0O+r8CF5TlmrqRgwYX33qDxhfFXqKmZsVdVj91p
Z4Gocn0/Npe/sIyA7odtiVoh3RXJzl3jhm0PM33wBXIWk/XDXbfKzjBNGJIWH1wP
KSeFqi5Xsi+g72cwip0+4YC7AYsHKveDCXDaDUMfLuq0McEXX5a3/Et4SkZiwMKH
7P110e1xLjFICwq1nPPNeqNbD3+G+WN2K7y++I1GpHHPhH9SfCI3ZHDPaUqncWOO
YL40FNzlACU8yKyVtTvDYwdO0O51X/2xtTahuZycTEKTTPpDly5AeogngSL97IBd
n8fqdDb1bmw+MjIsTo15Z7Mp2pZH9x/3Scnr32aH7Vdeee91X7gxAYakLt9kDocD
GvGx5TnYY1rXoviNuZT2TGpdBKyevAUAO3487Xg7i2rAaEfgYYXOmB19bwNLAvA8
2uf7iaecnhekRzUxNIbEj4vLz19PDJetpAh4Hf40SlABKNioBc3d+nma/KqOeZgw
s2K0xc5bP/zZOEQn+bG/jUiSEINnTi16KJ9sdDmkbmhf9Ho5XSon7GoenMFFDUqM
lr7DDW2G6dEAoxMataWsUTaB8XB2Zlvk3r1PoYuT+17d35DcFgCiEZxdllt3rlOo
HKkmLaypIyOT11TskKcY0hQfHMD+ig1buaqcyyIqOYwXkgxhTn1BQ3reAbAJW7EQ
TyWo2dBn+iimGTCxVjc5KqL+qoEzb4yqFi2xitcSE6Z2REhs2qdue62Rm5K8gfYl
6DNub6bhknHpiutLpNdBgQuqdeAxPR3vf0TH3jM+PXYX6t1uKPU8p1HMUJ1oHi68
jbRzvdBAKBHj7ZmZ19a/VspMdu4UjKLwogY5wAwhPsxPFXkn6bz6PE9La128M7zO
OM4kkW846Om2FYent4rtv5CPqCUNM2mszWI4rpjN4vydb+6wGJC4cZPQVqO5Rv5g
6cZWBJkzBIYRBH35xMi5XGaahG8KAbRZA1D9N2p3lFF0UOQ7IFlB+do0h0/G6uJ4
BtT9lBJO7Lw67ollWsd7BtnUFrLHI7cN4dnjPq+X7dKUWvqbw16UoAikPzJb59JJ
QsedeeZTgRin2nnvfIj5YwIzTJDkRqsfyfCmMLSeqnY3FU8meqYMZer2r9RxEidI
4iSyjdTYmmEHM0AVJKQVGSSacbTIL6kwe+g+wEs1OL1VJSHpGx+m/NgXNaBnge5Z
bKE/h0WS1f1hfrjcOCa2Wvkse6ot6ZJd0nqwg0i6WTQETpsJ+4KNZgdHRe+dgQ+o
+XWWE4OeIn3OAPiVMNnmEMdQunbJm7mQpqxyewfhouPwENnDceDz63hshCV6/wLL
u12eue/Abo8chmJMgz2pI6jiCkf1DZf5j8A5oqlIpbWNZfMAB02ZF+CshcJCjRe6
Rz0BMmvbDGX8SxBkRuT3qM5SDgxhdGpQZ7qNQM2mfr1p17pDy1Qjoh2mcxrtHufX
9WbEJ1zaFH/+chvu2VUfeiCD1ZgUWj/moeCFIjLL125gWbeRCM7Wsmd6sfVVoJT1
ZO2YC2oLGkLsM8ZAGblUZscsQ4MGcwVwDZrBrDsNBMjC4eFS3E//KK+VMUf/Yu6B
`protect END_PROTECTED
