`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XRRFNu0N62PmtteqDw5GcmsvEGZNgB7edrX/zmNIUYULnf5Une7mxvQ1aZ/aX2Xx
Kl4q/4dsmgWX/8pGvsukb1t11fhcUF6d1y4wdk/9HObXXuCTT6Z+n5VMtcgCzOHR
ZA9tGgCOk3yuGQNQxksrKJbR48yU3r74/5FCIiRU8AwvGTRwG8Wy6k/YKfKib4LZ
PI6pPIHCoG8in6ROOSCUGgs26Jak/UdpQ3QtRlnt7pDf2t+pEck5dl7hhqbnKGsT
yAZBRdg/bUs127X+KRcsd0bMgwnGdhhHd1nVRocYZSoWIpheD4SmHqqOgQx/sbVR
CYJROtAsUmegHYM1yCULlpP4IfcTnN3AlkfVAk9aDbOfLAGo8ZTmdjzmBQUvQ319
3vSvPf6PBsbR+Gzp2Htr5Rr3v2SCm5Rar3xM7kGXLs4uLpLWH7US2bDAn+yaIxtk
`protect END_PROTECTED
