`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PZTUSREJa37SJFe6WBV2ydeM0fn687oSZggxGUfF9vdEVjw5K6hdPF2Kt0wKh7iN
JOllItX/6krC15wClezqm1DDHIaUfJrk8SjkjVKBEJ3H12HWvUqFhjWsT9bA/HLo
pkubjhV2oefKzzbxUS47CSQlqhxFehoAqTLuitZpkhxVrrsDLjBxZX5DyMw2L1Um
Eewo9dNrmCBVpZcS+lTxJ5ph29GMOcJJoCOVppKvlEcpjy08TY2VfbLzzrojwhkj
ACMKU9sdgAwDDjUZtFHKYlERJpXPmJ4NwmoPusoXV1McAGqSUqDTf8uvRJtgeKOt
t6T+yWQ4/oZ5k686Go8Wa9L+sthVARFzpt9lABwv7h1maHQJzn6E6uiUCud6gpug
HcQmM4uUl1DUvlTz78Gyw0uDnTr/u8eGwHiIEhr9/cMti4A5lLeilFavNJ0b7Ykw
rG0W0TVqUJoRFjBP03yxtijsN5eOrrmVK78YirRN4xEmnVEDUJDTH+DPcQyC7iVV
CvehJb5Wqemd9DiezrCdNN8Bi7GcfuULT9f7Ekf8eBE4ArLVX+q7qVtr551agq4r
YlHBJjwX2vfITbJQc9s1qn7sfja/l86OvDYnB2fUhREIEIZj7O71WrvgHb53QZEe
RQ62batLnuGuV6I6l8Ct5JBL4udJFpCeR5oToccsrIxeeWcY5wnkRD5PgUdSGgUl
jvNMTC1DQvkKcmYpXy+UxWS8mjkgQoFM/zDSbJ7AmUQau7eDIzOgC4oRSYTbgxlM
/EkbKv31Mme+BokDCls45IiZdzdJlaHBdMtrPRgXVy6F7NnFWeju0gQ8vWtePxu5
`protect END_PROTECTED
