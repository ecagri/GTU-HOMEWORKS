`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v9o9yGcdu0tegIfDj0F4g/Zl5DrP0d/xtwgzXrhtG3ApTDOUgbPPbrYN/TqOFdrD
XOGG1n1MHi1Ld54znrzf1rjvja5gO+MS3n99mmB7F17/baOHRtAupOv0ao8pl0EQ
8nBGXwJvfZLl6hQYknZCLUskyDZl34ba3Coi0X/DpvBJii+01TTPx82U0Y4wmgf6
RACKfpFuXYF89mlXJ5bnIPamNDqfFqEqRVsO15ap8UFvbfhj/oeu1A0AQH2Vdt3b
L2sfmrhwlcZOSyWWUeRagyUkGnwlAbNbBs6WXG4yIfyFHsiN2XQ4j8zLDnM4bzq0
lDB0TAiRB8r6/T6RkNio6VkiNAsbxvHsbbEbBqn72mSIHrqaP9XUFhsI8Usd322p
o1XzA+WvwwCSceJym6x1JFYL1VYm5X/r2JDZsKDw3vY1SCPojubCAWA6QPaE71OS
DoGR9eKsdFoER/ADVyCJBuKi7PYC2KjCEP8u8k9+/N3+Y1HGBDZqbNfaWnR92Vo6
ZR7CDlOm5+3xLM9GVTJVYdJkiR2RLLh23wdH6AvCNW65YBNLuuHs7jhWdLtzXSZk
JOA6J/Bp0v98nlM0sOgj/QHXZpsvCrKr1WhyfMrpUbdEa7nwNjo0a2RjvmzwW0jj
WFH6KaTqC7J3JQGcDt4xDVu45b4Qfv/m4trZeuDrJlWrWEEbl2jPaphiQPoCKtHl
MNlVdrfos9YXTER71dL08MlccgMaaIU4kS4TUBjpU/FV59OMhfC+APwrQNDSAx4x
XjtM7dpcd6z1u2MOYIxs5TUpl1mnDTt2qquCvAqwNBhT53/yzPq2E8gOT8meXqrB
lgFB7vkqEbkFF5LokktO8zKXiDIaMypY0VrJnDNxOP0l5E6U4JkFSUI6HMZo51pR
XVeqBp0PBqehb21TBNYG59pR24ZVEeDo0TRPCvaDcff0MECQC8oKF8SUH4SUD4Cq
G74TfNcnKRxELpSqs69qYQYOSVb2DKlnnZWczBWUNB9jG2t3wm+CLPuH3+LXTYQD
STJWWBEVqzLCThP/ZlG/FjjPdv/s4Tb/SseOBk0FdA+golCF4Kx7KafYc9rKFaGk
m1NsjsKuh3xJ2cdjppLcNponkGgkl55XXP/XGSLwPCbL1UBliHx16EaWcu3vM2Yv
lZ1hguluzApfetZZgiHmr/Bwjx6CTryopu1YwYOzlAYyORG9BD4pxKN1a7/jmfJS
`protect END_PROTECTED
