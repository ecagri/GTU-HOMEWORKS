`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XjDsg6hKzRu5Dwk/NH+mKaJeYOrYHTlM9hc/vkQE6eOihs0FzKN8yWRybaUOepdV
MX+fUEPXlGVrlf7mcgFC56Lyau/DsDIU3+kfalwYz5QLfNVJY6Quu9QxwXsqyePp
xIszq8Z+tzeTyNTkW15OOe/GpPNHXWIcCn3op/uOTzoYYXr5yh5VtPkR6dYuZ3xJ
uZ2Fxas4fjTZy5n6EzkRs+5e6ztYjEedifxf1/T9Dcmx66f0DDNKeQP8n3xb41wI
4jG2YeSJTxJLze/fNcxZ33b62V/bps9QUMeaK4TqQAA5OuI/DT2BhbMW2LXSDIyg
qeF6nujPVu0BTTb/jYxQtHiaJnYHfukhIlvgr9qo39w/K/ENkEpovXUFuLXE01uE
RgEiopNgpDeXc6oO1DV5+DiUQPQeudpaIakYE0ib1mOEg+AkSDOZGcIzo2PsDy0U
dJeVSGQ8XR1NRWOD1Z+hAhMUdOgkySKbTCQXO7INXZGVzx6GeG6cvaq0sWvkZgZ3
FjbV1TpKIZazYHzYfmz0iz8Vi2R6mJxxO0ib703yP1kTOY3pbrDPNatv1yjNPS+4
VANcYZBbaMWpKxrwhWew9PobdnNz8fqie6QZH/hZvRmek112zw/i7l377lWXEaIt
Dq4qgDqJViB5rb75I+U3rhuWbg1y2gKDJLGiSAQqXPwMZHIcUD/FxnVH+1NHpqqK
h4qLggKDMVxsZUqNSDYCYxnhNJ9+Nt5luPoGISJvjLMpqngLS5yEk/+h8iczdanF
+lhYu/5K7jvHS8t1IHhmr0wPLknc7Y/HBY79dkg6ngRR4LDSJJpqU68pvrwcjzKz
zQzcuz4ZWqW6mD6pnLEbowd03UFSSgG7+dPtqIvJS5dvO7UBXICZnWnvbzhLlV/b
A5nohL6+09CSQq9ehn9HEOAOHsWnjKjITEJJdFJHojVkrq4anY2s2uRaxbA/FYZt
4QiZ+VewPRvIf99g51z8h4OT0xmcdSQLGWpGIHuukC7+jvEKwZvw0iRivsCBiiu2
NEUUJqh1oqNAwZ9RJpBQ+tliMMEvNqDnLQCuHGsqMtgbHvlQ7LZWtw6wE8D/lJ3f
c5cmLy/fvT/QXnubt4dlNoLFTZgi5hSNVOV9VnxHXRs=
`protect END_PROTECTED
