`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KoFbGDZe/apRDI2zRMSvamSQ/UuIPkDb4WHfsyGsqWuVsHa4oeKIConb1Ng1Z7rW
5KT4HtSUlFnIkjZoRRtb7G5KzoMlp10w05sw/kH6Iy16PzXDdih/3qVwnTS6ewOk
Xd5NnPIorSjgoxNhxYEQRJCJ5kz3b7JzOH/dRoWO+XErOf55saKx924E1nN8r6mv
LEmDP4mVCUqKiDWY2LLru7jZB4xfyS90+ekzxyImfcpFXkORKHOJjiyNZ2GOywEA
CiKgjTXlAvsGBs7mwPzUyIzUOWl7VolamlFwHvCrPw2u+xcHCJNNkNpN/X9tS+4V
C+7twJJ613gAclW2w9dFOJZf5FgyZg+DEH2UAUluAEa+6opYTzmcVyAka9GLIU0o
iOp/rr6ZYkXqJdzFj9kIbABNuWnaFab4vAMih15cVlckAdCqv1VDUXOF90S11DXG
FULor/KILGIdD6tDtJl4DaGx08dTGFDqFilq/gZCEQ4yinS/dB7so+FJaPxc88sr
tvS3u+hKSiD3sYYej1JyR90zL9yX39FVa2yqPhBjLcCLjgF3hUOSko8Lr5sb3s1T
16DZEb6WPAv8Druysrv9iu2u0eBj40WnYytFvxKPkEd/JmuTaOpd/p5k8MSJ5ss5
lupchO88FcyePB8024LDjZqmBFNE1dqpocDqI/o7vE3HMWWxZq5yxJ58/q0X/XAz
x700bAvIcEFF6NvA/YkMSTqJPCREtJOHFBaTiS0cHR9I3HtjM29znV64UwNzPvY4
zFjUKhsypc0IfYp+k6TZqxKRU19FSfTpfWP9MDWP8ciVBUNFNaGOrXxcOMNoev3e
mofCESyUA5Vc+EbIAXwOdOhHbqRzyRr8YguM0I5yXxN5FlBK9TzoWyT1/5Prlpdg
OSrBwoORpRcDtWrdJkXBdiK+OcMNRSWjkyhI11lbnJqAKirMJfPsTIZzsv0cAfa6
jqAlLnsn6DqD2jDpqdNZmhfxB1XZwuNms28Ou3LtDDpESOQyY2Uh0GRJYruGfsN3
WZO7D3N5+NF2XjiKu7GUaNI6usdX44q7Pm8D4dxHwcir+q4+Pop9mSdxCzETemTV
K2Czgu0kV68i+nBBtWXJn+SXejnjsdpqLRius9fgudxPEbp3Fz9FvgiaZLCHyFIx
KOcLc5JQl1q+rnjtvSIlH3rZsPglGSDt/walXkb8nFZSVF9fYwp1MdX5lldKg3dV
tQb8+zepZZNqFG/N4PPsEJwBq7Ndyh0ezgrrOYwSwWkKEU1pD4lSDlFLgZ+l2x4o
M0Z8XSxPnsBEUggOl5LgRbjcpOnLkOC97iAoQ43Y0lyHVpyUK/9qNYnEMzDKvg8c
EB+ow9N8lXno5MY8ommHqwyRAjBGKMo1zlN1vlAN6VZebaIhcn5AuGExDLHN8wXD
oGo9REBQqZk7z9EB2/HqSz0JNz9J7zgW/nMpekaiu/J/5Jg0P/dHIbtsOBPJ8xeU
Euiz/jkLaufvxIHaV22ONhs6R00vkV0fmi4umi1bstlENj7aY5+t/Z7xjM6aKmaw
XziwSJefPRg0mD7SZ2nX+KiiqAGpHwAZSepVPanot8fVyOFN2489WFTQ77+nX58K
C9tl1Xg0rsX0oBhd71utA3i56vWsJxh4X0oB0rH2ejBqYDlg77jI2FzGYvyRTrJ0
Mderc+qOjJItElgOTRnX9LwnwrVviRFH3PtQ7SziOc3MjL77WOREZVZBnDE5e9IP
+51usY5PBZ2+Z1IuBFoQQSSCxXCRIAN+h2USkpSBwE3oUB1cQ+F1mYuOartXeh5K
mjotzVQfm2TezS/GOhuM5zAYC9IE6qO3JOtC5D8zaiCq7C6cyjMTxcZeQD1t3Iwv
NrauXcjayE5zW7OdckoPULWnPCcnzQAc8PCMea5c57Kp5mL0+57lu3mC4vaBPZlE
y44vtiH8lcRo74t4O+eoPtK1HXaOTXZz8a7zSpk9VB6i7YkKIHa6EMKrB+7pz+2b
eSxhoXOZDc6wLp0j+yGjXN8SNya5AGWRkEz7BmAm8/wTF00M+dwKlGtSEtgcjObg
foaW946Vn4FI6X3SdEupeWvqhaQhl33SxIBGAJV5mDY6ycbVEcG5meVc2VW8oSjh
Q3sHydLmwlR4qTxgXIDMy2AoJjs31Ipt0mEPyt/gGZwFyhu4tSu8qkKveMSqY8EN
l9AKnRY7Azla5Q67V0+9jAtlAadermU1tV4qNyURPqtYw4dOtGiU55SqwAD23byl
1RgvxTQm/bnSjjxVk/jqcBjq6CANGGyw0RGBzwQUlyXlUjZQGucvmo19lKOQ/Q38
5bO78xeFOUuE82kxCYW5DNgnraVteDTHmiBw3wyzjMq7Wjx2/oWfzxya4L550zsc
32Mn9eR2mtCDSQkwY8FNo8+vuBoiXuXVzFz9SclHUFnU9SexbXQIVNM4sH3oMI1p
9BvDAPOZ70rnZDX1c8LGCN8TDPsks2PVE/mpsjmD/Sw0/55xvEKb5f4ilRbDrSj8
Sz7Kk3xoDBq1MJ0dkOg1C8MuhLyvdBxi4GOBSla2y57MjuwVYC1mbCAmjsMZyvai
scdTfIe1S4+TvewwRwuMKVJ8IpYOI+DlMvaucU7euJ5soS8sns4cvlG3FfqWQaVW
Kv7XLs8wbRrkNjPOPMw/RcXj9pI/O1T5ZzG/wNn4UHDGms6i7RKhdVcKHQ7nktuY
SRTVnwmWLRj/R0a9oMBiiDahHJ2d5SAtrWdg6OF7EmYIgxvT2roafopdx83Yprbe
tLBu/2pUeHS/fcVHas/YxOf2U1v4NBbx2L80RdV68xXXy0uj6/mo9KtMXX7+MbUR
CbqB4XVTSnO2xw73gygDVohE1NV5fqrvXA4eGueWicY0lDenH0tBP32FRd1mNmrD
aa89hEZ9LvVTgJzaLMJ8OE6KmXQhpPtRIc6cTLg39H2zpW8vI1RfyNYq0n0X7egA
BdPCDWSgK0/yh96F4b4RwO5k63T8RYyRHimzzSqjqw3JEZsyhcKlkS1PqXlp6L3f
Vn2GyARpNOsewGY9WlBc/ACL+mABu2tX9UOlOWjOX+4qxNEgcTYhZ5/hkNpnngCN
6EpPTtt+lFFZVYtfcuUgT84hWkU3sOaaRfOuj+CY0AbY4m5mD1T1eLI2ncbmbqbx
Fke0f4ODTLE5tFR/mz2mWCEyxmcjbnSNkNdrpuzenSnLUDKk2csGcN3Z5Uz8AhkF
eSg7WxEVxuso5BhjYIOFdXzFbTfYadqxbDHcPZ4JC2oRsIy3N/F96q2XSRSwDoGU
PEhcf5ZgkghdOmNSpRBlvrrQ5EbydFCa6obuIDift1kWOXGcLhBUQa16G8yBPI1C
7u89je0/bC345Vd20HcSsDTBRcZyxaht6L8JmKnrekasjIkVW2oJHuXayUXmoxaP
24jLXDQjjozhkk0obbHPRvRp8wBEyfeRuuk0HbQwfqhrabXtx0aygA/vs7MS8TPd
qSzFmZg/Odrkm8gDx0BvcrKNbC4hQcpGGY7jpeGYokLYfQAGL0X8MdMxPhffYwzv
nKc6xwenIklEXhzMa+OXBF0ht4Y9nXCyO6ldQlfpIRiq/b/LyNCi7dAQVujMymlY
jg+jP6QsfbY24r664Lb3JifVDbF9nxMSZHlwN0QUiaOFQDrY8hYdnWfNXH+uQaFD
B/Cv3P+p7b6KeSWEUGhwwz5XQw0wY8OuSJlkNhnoM3ywHLeKZa2zjWPu2C9Pc/UE
YlSZzZHezT0lDZRSk7uON4j++OtImInq9RXZC6So0lyyQmmIYW9LlJgMTInSaVLn
WH7kS2i4eiLivZ90W7iEGxJTCFgPbvuPbXjD/Qzawvg0wwckpqQ4JPIlhLpauHKg
VqVZr7wOtwYMP7Ko20z7IdxYaL6GcsjUdQ7Pu6P4R17WTLtV8fwxn6xAq0WlUSln
pBacHy56hku0gnJJbVdZWht4HLegiPbRZGLgp7SzcJEJnp4Her+tBTSQSuf0Rvlj
ZAlVldvCDAoDAb/GhxWOkPg8x8bTBmEnNeWcv2sz0HVCxMSFNW+4tXQZ5VNpfql+
Wn4hInH5NFSQif/jDYyhBoNwdImtosbS+tDmB3PkhbjWwhTCQ07gUWbfaCC2uTwK
H94kmUcBeIt6j/A4cYLx5n7ekw6taz7OzcDEloC27b7lF4JoMJXP6b7WL6j53azJ
gfhPTQHZb2LS0veoSF0p94tWDJ6PAmbN6xPldaAuDqdIdKmaQ62fcn4W9NASsXsk
6bpOQ9aJzFSKVc3KZmq0js+jyiZiO1YELxhr8wfwOOyol3NqJWXOZ/p7q8CcEU+B
AmDlK80umUWLvcgQahVpxBktLjf6QFK9VgweH0a1e2VfcGGhtTGKXkRDv3iyuzHN
zkaZLZda8V+mr9jizlcA0/dlG49BC9ivItQJIJ7H2+ofCEnYDHfrtVSa1NlPG1fQ
VNj1xY3zX7zHQPznqTp2A1YRDFJMO8G/CpMjy6vNpASkHJkjzhafsErgRAfbktW5
7ecr8N2Bn1vE5sSpZixJnDwtVQ+gGiPSu5m9N0+0MbIw/7bMLnI35mHuhFne/4gk
P83wsxVICxpR7fDr8UJ4EfzgoM/nCuKEm7ci1YcOfPGem+wIlmJI1m53fVxICtTd
Hx1JAMubEjf753yjxzGMQiuae30AsmQ4wKorahtRFuIVrmf9YqOcKaVQLjHAziHF
KEQDJ5KouawjVFpLtQtttOycm1E/ppFxt3of7CicoZKH+f7y1S1uE7dZWzq6Tdqm
OKq+sJ9OH5t2oxNvL3KYjc38+f8Nm7agMSisq5SGBTlvnN6yM1WSvAxPPiZDLMvn
MVmn5ff7B1/x4WsADkgPM7oDRLt5nJvwlnM3ITl8f7eiSA1vYSqcII2W33P6u3pa
lZ0zuZfWJS9fnOBd6rk7xUPF8ncEmJFrq7xTtYE5fw/UvtNxamerJexjizN8nzwu
E7x8xSN3VYu9J/3XBt2YMTTXPVlTfYaSYkCxfj2TgJ5f6Q1w1ZPXpYvCLkL4ZAxW
gSXzAPn97yOVVRXOX/1WjsajxonZQi5wMMtPdFOQZm5XUBzLS86UJYEGhHJID/M1
T4pVNR2pBMhmgAA8/lb4F6ho7WKp3zm8oQaXxGMnmQoISDJ6qKEtsrC+9q+roCg4
qboL62A/GDr0e0J98sCYzaMEWYyp4ke4KJKdKZk+jkatDL2cE15WIm4AICFC+V+C
x4XzBUtQX473qTAgOB5pAVpV7L3OEZWGILTqVDWnvpgepYIcn2N8acwRBg1t0diZ
ra6x7yO6pMt73mc//9dXDluE6eH1azka06tA7r5s9TdO69HxLmwvLjMiLgV3mPiv
H2ALwQNQ2tZBDuAUNEjohr6okRye/qEO9kjP1hg7o7Y0uHqOFrnOB3StvcyFyMJY
rbKvsSKa2d1QO18/ro77Tpl8ndAwAjru4/R1KiWb7YflHTq/4eY/n0mpX0sOQvYc
z9G9FY69smH1WNubSHedi1JyR2NqAt9yCC+WTTe5Ag7en+/Q7+MDZ26A44wSyGKt
8wruWuTQOL4TR3vQeD1++zIPPj2oeUC4ZsDfcwocan4zbcwrmIiCmNgIJcqorHhW
G4u5eTqzwxTySRfYhcx/+2HGP2NPg61QiVjND8PmVk+1An8u+jROKFN17VEdDsok
/Qliv3fB8u3JhWKYF6CLaYHxC4BYbLY84oUoabJ5+Q3lljxAWliB34IlWOMgTX0K
6pMTvhYl+jL7yR8p9uMyQXPgqzuNOnf2sFpFgu1SySQZLMS6bxOX1tHK4bNyo0HK
nIdHzhFEBaIu2r/2Vhuy5WG2b5D5zJ7n1SH8aZp+Af11YNpht3n67E1GbAqFnBOJ
C12Rt2ENjCiSmQC2YhACkZCyl5owVg7oLMFFrgqWwWdNmBp955AbGcfTxE+Q2V+K
Q05cj0MF9Rcuc8OpB1sDp4Jbu+uUYDXRyJwrcDKqweyz0EkkS2/uRfnWQNegFjDz
0hXcFpiLSP6+diljYnDrRApq26eLyIEayTHMKfO2TKppeIMZWCFYn732AeG6f3ad
q+XZPc0JitZN4y4M/3IzcclH36snlzMJ4del1dh9Vcy2Uw9qRb2NXtyD1FK8KdTN
fmeXU4LVR2jM96y/9M1vBpgK7x9G1hKstQ2VY0zIBxXCi/vVSpCyPdp2UTJSrfUA
fMWta+Y9u5OP2XKcATO0W5oDvmV6cIZzVkGyXxGo5L1RrGlz/fUQ2ORJctoq0MbT
FVsoaP9aT1qXKKGfXK78ZeFNPd1hPUV2aA7TeRlbJ0P5ApOAIXFCjveb9dtIwn2i
qp0+PIpbm04/IHNark3JVbjovkoAkD7k4oNJ2x6UA3tkWvaqMbfxhYvB2MFy+dK4
88tr7OHljnAua4+8YMwBrpViC/ddi2S6LmJAfQO4faC592sEfeXfmxcQC6gzHc7i
bx3L7RkgANw7hWEvQXSl0KTDJQs1883RGuGZSUIy45kVbg5eNBQEmrFyffX3ljkV
4PgRXqcViRTzUekAf6qbtHrEWyF/h0ot9a47ZbJ4fFv9+E0gXyBqAiltqWLJUZfV
tyvyFPK5t103rZ9UZdd7MmhEtXHuQgLPZ29vHeHTjza30Hbj5EMEBmfoUjultv3T
fCBjJ8rJGSyQONmFzlOzQKTOEd1j0fAT4ZJ5nG4tXSp+KVVkSYfVB93RMGhTrwYH
MFJqtyxrLyiC5cuii5aLTaNJJwzSI7/13TeiDiO7qV3GAa/Eymc3lVx1ltItVeuc
+oSbT8bD85vEBrcsKqFaLsO6JAbtfsouQnYg2W5rDfLhMyaDQFs7gWwlF5211fAR
ZvSk8moEtIdPNq1kPiiTcx0aIVxFLEu0OPR4mn51srBx8mweeEsXgTjwsED7Bu1k
GE487+w/1AtSWpZOpRfpN/BywK68X+HeAcdLCA4m1NQQORtPgt1inn6sl3w7xTXk
wpsZfDxO0ECDwPrX1j40w7yW+IWC5IUnR043cWjOmo06PngyyM7wWanYYkyUew1c
88eaH5OyFecSHrhMqNSjKbOjOunUzcklEYpWuUmmy+g1Od0rHnyNhMdDug9bGOBP
xTjDMeGIUiA/Xl3FCjdR66Sfj9nwBEURg+SwdJQZNSqsBaq5AaemX7uqu/rbJ83x
T22nPqzkDAp84P4nHVSbONcUyKjyhsGswjrTFLx0IFBhqgEyVK4MiaDr4kuiZAge
Pg8UwFE+8MzqtnTWtfiPOEfj3BXnWkMdz2fxI9aSIEO317C1JvaJM3rF3yC4UwhN
l9uD5fEnw6y77twtJ/kFQphMtmffrEaoqLU0G+56pCk/t4EltC+TtAHKjhlOaTyc
jN3e4UN2yf98LYws1X2oo9laefIC5Oi+8Jkaa9gL1R/BQqp2omCSpnAgwktbgErm
nPoZzleY5RwZnM4gvGq1JbK7Cs7y5uzdMSlN/QPrs7yq8l1BuQodUIdPwOdyj54J
SQfU6i9LZ6KRZWYY+1pdyVELkWai5Oh5lCHwXaBp7eSUu+M42ZZnhjE2UnatBvM5
LoD9dlbTE5Hli6FXiCsX4PFgxfJJqRKMBJzKGVnwmsMFe3OFnUwTyqNvLDQ3+Ylz
kXBBfivK9R3LLZo0xyRTTmdyFnQVcoOBti2S1pLi2C8IExTyrsoO5pwd8ZKCJzcp
FJcfRlzVndKy0uRqanD6Wx8vPlGk/Qe7KyQ3CgGIOo2NIqlXCIzdTSKZEENFAp/X
PcUCKyPezeLCvA0puzPjiBTwI3QsCYbQhy/PuJNyf8/NOpPr2QZ5R6J2F0WLlLpg
egPi+gGX/CFHU3Z4DvhzlWHwdJpeiBWQWPSkURHrWkr/pPR1i0MDFNZhP+FXJdCD
XtueOZ5Z+S0lQJVo/1UmOjbiScGOWeKtAhKfuEc6/uV0t5SxroOb8IhM92ZQAo6Y
sVUIq91EQl7FEUSU9GuuiOo1Q3EiQSkq4wJAaXVuGq3ILkQFP0Gri1/yXUE4pLXf
R9b+CyqJoxIVKuO7MWQ6P0oS7SpJmVCKD02P2u087iavgq2q9HOqMzQzCYLUsMGJ
F1VopSR3y7EJ5e/k+9iPkQqc+oZW79DAnJWUbxKba35brqzRemJLkQGo5E+IwGDT
dgIOojRFHMjyeEmcpV9kkS4CTxQsN4qWv7kxCMKYD3hgB5tC2LHOYAJjZaUdFp8o
orTcW1MPIr0cS5XqzhMQ7VhBSiyE+DGAGqbNnNBl3lbCqWe+saY4XpiUMcnMO/Za
3lBeGL+N7n0KeawFPyM0Wtqq+LkJ8iT/JwqcQ4k0QPrc1bRliCxavvMLO6b7YZ6f
ck13hAj9+XnQ0FwVPIJc/cBsepyeS6fVuIpMoJs/FfjRvLq9sC6Ce5WicrOV32bT
EnusuWoc2yeOp7De1vUdqwrGMzmpTCUS1q4yUjLKaSToGmme+6m32GxJatpAqFDZ
oxBVABWmnYdLqCjquf3GkM5N/yKwbOOihFDqxzx7jOOMIiWezvOjd4Z7YacaJTd6
+jXqHOoLqVUhdehPCRwVAjklPA1F7HKgx4ic6tBsnp8yAGJRBaa+5mKNEK9MU0+1
CQ8Dnz21jDmGYWQtPK0dIzSyCJtz0rl1JZnFQCYFQXwy+zWP9by0Sa6gaM+DsgjX
+Lb7NQuZ3Dldfyp0z5EH+jBqQNuaYe3QnwZpJuilxmpukJ6BYlFzGgJIShcxYqy5
sR+1IpBEQn0dG1gdSpdNXKl2VXQN10LW0yYzdBQkW6+n8pTvO68lT9N0CqG6caL2
SdNdHAxJAnkayNtiAFupc0/FLORBVfataa4h26Y4fcUxsCWGVn6yDtoDtwh/Ahuk
P/PCZSmFET79g8ZybxeMB/U13OtQbu315UeHrJCNhJLDVWr1Rmil8XcsXAHHjZ6y
VLb57eVKIMO8ZwsPLP0CjIBZ12KNb1O/CeOEcPBZ7jbqlnAOAsIUQBUFnVuvNdvD
SnnBH2Gklvri72fW1vTgorn0nsFMVt0B0Tk+F26VGuj6qiFffT9tB6blUeF5sh2D
AMY6nhSTy8YsKWzbTdvCzh24sk485VXelxGJPBkzQUYm1bKPPvlzxdzTRWnH3JyT
2rbRit/0gEhF0UFoK8mWPprx2/84cS4pElsA87pVPTHV2c0LCA39+vXqkC0/LASY
DjnEZ8bMuDH2VGG1YAYa5p9JVj5KHIz3DbIUg5WK3dbm89FlAa1brOVFh0QiomFT
0w2xjcQuMoeKpBVedjj/WfUymi3P9KOuA802zh8LZjX1UHm15RVFtk3AV0ygJ9Dn
/d5Le1thYm6oIr/Ybs7C33YzH/e8Ndht11b6YmOlJB4B2sDODDaLZGCY0bvGCWfQ
FxGmJ6LVdi5rZSl9kn/5JljFtbiEKrL+vwrae42hrfFXFSlcg3vAr+2iuTjz+f7u
/q84IsXuWhpUe0yE8vsjBoMADFCOlww+Ky9szDQQhu0nbsi61p6lwz1pyci/KVSA
M7N7cHA2cwGGL3PGpE6OXRenGX5eknduxBXuEjRwPS2ZzcVOScoxd/8VgVXbfd1a
FoChyqQx2CdugJcVsXJ4pv3wqX6wQ57fbIHlqDogqpuFhcWdpO6b74q36cqiRN58
uuTVXJScGsgyLzdZbN0wrExzz95H4FYBh0hYc84GHyHmxH8cxvhlJFptnuf7Qkg2
v9LK51dQnZZ+MZaCDNG9jLBodMTz1nOB+Hco/QBXH2lwrYVLVeRaN2OJRNShjqrX
DO0VnxGzNfN3TS/HzMxczJSYtOWc+fdbbKbyfRTWJEAyPJBru1bfT9dEx/0gHuVn
uGoBk9RKuRn6Bl4OduhzwoOqd9GVLh1HynttDM8cQbkv5B9oAgtkGPUaaOkVgWb/
tzFs2H2BryAXTvSK+wbsBWO197tkRxAcgl41I9kHie3Yyd4JECrCw33tWVQHuEwt
m6a0ibq4lBIhy1mV1DrWtc5c0U6zNr4I82g2rrA1buGgHHSUS978nXnOm+ZF6oQZ
0dT6BWDV3a9MNdS082LMUn/RsddYPoE/BAmpQFfXVtDhEfJtYCnEH45rIr/hs30l
Av3eNacTBtOP8LTNvHWY+yC3hi2phxt41BjDVdpt43Kj7vtkB8EIpWImQRCcrRCt
SVnGbvmAzb+QyiA4EFOJCEV/1DqdM++5+f+UpTQx2qT9btTgAEV3pKb5ZR6HWBvc
0v4z7JpNpSylRtn4UtvzlOEyAqg0xNILWv6kyQ1MKiXq5z1panO+DTXZL9yviBz/
aN33wwuF4B3rpnOKDMwFyx1Wa1pxbSyyZpltrphM3izPCASiibW/6SroNSGBW3D8
QZ7Oa12UbRcRDQfxdfbdziYEeB6dyarcrytg/+64fE5iYWimZUWHuZTQGWczNrxQ
3f1XHfH/zpmqf3b2i3hZfvvyplo8lsUmedZe100d+E9/TQyIcLCiCoFgjEY8LIg0
aFt/TMkpwKwk9KKa/9UKJSsc/pEzWbn8CVKby6LmuSldJm/WpqMBeScHGIT/CG/E
D+1xuIES06yn/iCUdpBFLisGg/sBEwUItcFMNF5LUZFuU8pWKozkM3Jh9cFzuH8n
/Dv4wOA9z9No+Ihu0Il8n1yCUFdhK+lZmZQL/YzkgeIyDBZ1it9V8r41mRw2Iy2u
OVRb/6yiXJ24ykCieCz8DdY0OhbsgfhKnJrGPTW8MJ3r3WxC8eo8+VgV8wRrnzdL
O7raOuiKT80/sQLCUuAc4YEYBfHZduqWI8ahxMKOYYmJvWlHCuymvMTq8ebaiEZL
7xHVOClv76gdEy9iKX77zMtMvavxoOoSDHViNEGrfiiU5lGL5dVcAd/vUPHG4tF2
iK67Z7rYcB/7jpcEZ9wTbx6dYdVHd3LHBWVjjbKkZgNbRAbD73lqX9IoSfdKGGUy
zubNeNxOPP6GyOOT9ZAt2XqAt581oqkDu1+D/Yjnc9XVdbHw6Yk5Az1CO1Qriao2
xi1ewk87hOTNBboec0ljjPdvV2asEuSktpIKe7fSxiVs1QWd+FmU4pfpFyw6zoK2
u3DcqenVtBydKQX1c+/UuEMxE3KaZP+T7VGp8YlMuUcIbp6VOLZrLjDmZt3kqIqX
uMmbmSh5sPHx18C31gUJE56NUup3lUHRgZ5Fj0C1DZD3zfWswcCVznmotyos+0dX
xT1aJqerL0yDgUL4ePfD+qTEg8QuLJt6GgGkOe7X+AzUkMz+4JcCMXNYuWU8rtBn
AcOcFeOHmRb7SrUP0XXYyKCfEmFC7IVZ3dpwYWYUnJAuUwoyuU807QBmlpA6Df4G
HZjS1iMdIxesx3ojlUqLzfxkRAGbyrPTbtd1YkzdRJ5o6eV37w0N3lQ49nXW/tNQ
FxtfisQ0STWgsughlaOgsr8kf8a1FDNtJgNqTpS/Dt9fT7C+TgWUdRnks1YVRfY4
cakvPr27G+tCFymSi52euoI8ELNxYJ7a5vGbDURBWWk5rvHWj0v/qyYVNZuughTk
gunkVeCBLqH22N4VMAFBW2/nkKPWIzPMJ8AxQOMDIlTvvk2OZbDKKMAN/XW9T9Xz
PzFJB4ekgfcXoF4mLwfZWUqWe4709SycH5rFCIM993cD7iLMIp8qvAVnG2zvpZSj
7YqGv+SMztPsm291U8Cm8lNKbsH0Jijcq8S10TpcfXcBAVlea3IiaHs1z+HftRla
ojwoBbnT/wzT7J3g3a0p0CzU8xqBBC8Sd1L/00fQf3yKJe9k3ORobwGQnOjwTIl0
lSsrx0P5IxZu1ITd9l+UtAtynAO2G0fKvPIY4xmTs0jTksfPXiNE3ea50qLkdtaY
4xOIVRK1qGORMtV4GmI5JF5njhiPZGw6eoSQg6WsvdWVMu2M8N1tlTs1AgsBGNsN
mbKkWyoM5HxG9y3mdQ0N1yxdRNvJtVX6WS7ZoNZyvwJ8GqUzwkx+/tDoZHOD3YOt
oa5yXLrQmuTvAjsBVrxW4ByPs5TPj+csckijvKn60wsNlhpj5zAETQ6RcDLPQSTn
EMZcvfM9Q7C4x+H/opWBe3jQKvfxFAHHkUUM/9015Mxx38y49n+LWUG6zAuEap/8
atDeyXhVWXtHwyNVgdBERkfY/JFKSnvTOUMdQiOhKQ+zuDeomBu0WA8VKmohzzG2
dVn8OrOh8903BtX4ZaYE6Ry4+qAePzjM7zQapYYSZPVpbka/tTuCpu1qQz73D8lj
bYZzf3CUwQwFA/ynBF5hYbEfWTZAW3VRDq5Q4rchLnt9xG3j8R6IQtY9Jwv+o/OY
TRF1mMUO/PRaEJtqrGVHIZt2ma4zh9Yw6CB6gsLBC58+GshtU9GwywM9/CF5afq0
SQvWuRlI6J0xKVPUq2OFPxfpVnN/e1v+B/ITanJ/1c6xZxfvxosy7wXRkRNRwBDj
Ys2OnmUdYXJMjiIGtDeEIzijH/qJePaSZE4oHTdouQaoLQx94Gr+2uGgt2bEbcoL
+NUgujhpn7PwRyCyWB7L1W/4r+b4V5587Q97m58Q9kn2GtJ3zLameLTtlPhDKgtR
Sa4bFkxWPds/IpXs0gOQ/RWX037wLhzXzFJxdng/Ze2TaPq8eZVYelMp1VYND5gf
DQ9nHpz39dO14zPcKL1zng==
`protect END_PROTECTED
