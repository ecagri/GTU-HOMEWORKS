`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FJd958cw11FwNd25kU6sjF3IAwK3RXy9saAqlrJSOsmEb4yvhbZvgL1w+q0E4db0
MKORtdJcnh7WWqfdLM2nV8bMIHIjjZEeoFUiBsp3Rbqh9h648CEy/GidiXF11CzD
cL9DQUkLlIhNaBLQ5t3d+QiHd5f3JPBvdvvIK6qGtWjJ1H1EfTKek9JMe0Ed6cBW
+BSgngUCx8BOoUjMnMnVFP7AvX6A1WxUt3RiqkNC9STaQ0b8L0938Zr3ZV3vMLfI
F0f8KVZGTCAb/9NOVIR649VvR9QUINOVxYBPX2cXQfgv4J6GVJAS5nL20i6Hr77Z
bRKWo3Sm7ZS8dDXxDexyEjtCwPs3frCXys3l2GnSPrEsHnCqNmT1swmLVXAGB5bS
dj9owQyKsBRnHf/pTkaDmfEJRlP/M4mp+Mo6hsnWU9kWFP6l/lnQtNLhVRG+ueji
0YQws2pdDIFd9MY5t3P4mEmjyy9JuI9SdcFu46CCZ8TPKRzQ3B0y0pSYiagwXgBt
fP42lZ7Alo4EenqC8mjNd1zsehyNE3DUZfe5m38SwNMyVPwAH1CG2sOt8KYM1ahR
nUu6GHoLBzAXAur1zjgvJ8qNfc32VnaKcddJRfWP+C/wJvpLh5jG9V1xbQYFlr9R
WZqZi6gIrd/+wkmrvH+XKDIunAFZvwwu7TV9KrIkolwYJyod16JMRjRzvWrF8ijK
E7w1uiiUB4taYJI6r9i8yvL38SZIfFVs19tK4/uDgg97rCUaHUpNbSRStoxU5FCk
erG8YnaRaDAeLrv6cZ4LlbgGgPrD4/pDsfNyFwU7DQcZfC7tEvc+miyGTWLSM+94
vbqHXdQ8gpuxS1frNP4ZwlxSBaum+TPDxcLNuR3E/DT5jHvE4GmfpJN51cuN/Aj5
JOqyMoUHcVZsbr7ncgWWScwG2G6HcNfR/J2i1tBC+CcjrKkFlY9ioM8SkWHDZVoS
KaZ0xYDMy02ZdI40AsfMvJZr0SIq/IjlkdoMvHUZi15jd+vH5xOVIW1oNVLMgUa3
JxPdq/L2eVytZxVQrXYw7lsnqlmMB7jZeUyC8mGGEXV8wU3yEwCaYSHHomr7i1yb
UI81WsvRof0TSD26IwFyFaIiKgDH3qsWAlHZXbgZcHif5KkbvsvaanKvpJhMZH4q
7sfY+zcplU25LKudKD4umcdcFTIKiesK6TPLxI92DLjsrJ3N6QkxZHG7tYaG/Fob
1KE8l5MmyDMXPmTxrD4Ap2obDF/fkRMaaRhXdh5HnZzOjLaNaHGzxvtn6U6Sk7WY
6Za8MvuHie4hmx4uHXxmyF+1Rz5KKQ/6oiOjl53w6/KnkxY4a9aEe9RYeabcArMU
YcX3j3MNYEUzNVzZhqBJaPC5/WKxUSDXanK/zEG1dKn3syJ72qOpINQgaE3BYgLv
dcQIZCJ1cUwxXlzjkEK5OvlN+kDBeUiU5j0+2dl/iCAfXDomWfiBDCDWGuvmyKCk
oycXmauw1CqjE6KUWad/6BM6KBmb+n+0DCoxPHOSzAxion5/DzvUFrMLY7yMOLiw
cHsLESc0x2x5Z39eqC1eaDmlDb52mHkZuqf0Q7WGKodw+A/k+yUXB/Kx8dszS+YE
p4NiLgMtS67il6ICnl6wmeFYIrG0lb51t+0cM1m9O71HKbyvQuptAiN2YH/rqh+0
e3Q2oBcVOdMKiFmYmOSNC8PyPPXwb22AphhdO14uT2cbzywapmoT/wVDeGmc89zY
goRdBio4CTw0aPtdhf7w8ciX3J+67wJQqPDd6ojeXNFv5qtJxMTDoT0JwyjVrr3Z
ZZjTT3Vuzp2nvRvd3BP09WDmOGt8LJVd2ijLASA13BMwRebg7Hlzs3R9d0IHxaTi
b+qx0dzNp8BRlD9yZAB7p5FRmRxnjSaGKWgxGPMyX0ZjRsvQZTYSZN85C1S9nIfy
Q01RWnKH2rIrTW0SdiXQmn6+SgPmAQERGnxd9HVr/GwvjxiIJgLGbfsCc2Ciz+Ht
WusD5Y0twQM/TCpFF4AiYNCdhg7G0E7MMvSSTxBaewo/6cdSdIgkULFsPf8HpsM9
NQqAv7og571BSDCaq2ysP+fjADK6FDxgVfz1+zK+/WFMc4DhBdU2mK5RjYCS9ptQ
xyc0rC7z0dGfmnPteIP+86XMmWz+vTpCKu5sK6HOhrRBxlTR4xj9DRuwhJ0lD3Sl
GK8Mvzl77/382Sjh8ZUQvot96s0e7ir3WIhdDUTufiWfmy0XbYbIEFy358bF1SBp
n/EtV5nI4IYX2qw6/2/JTmUR+87brAFoFW2ZApbkQemp5X+7zzpsYjs+wBk2Y3D6
26aSbLdGViCO6pG+0PVbzjYeqolj6ViOKUH+oshfVJx/dL2UoPHOGl+AieKeei1J
ZqfZZK11fFdQsyNItjb2S+hMoZRkUK02Dxrc/aMAhswfy8S05YBcXhr5stv/mujL
9pvSJVI5hRTEqrZI9FCB1e0wUlVpDmmalW0LtsvBL3LWqULNZrM3vxrm8Xv90xDV
4oZDkLBicgG/PW7zqT68bPK1bRXuFPTSFuWoQ7ItisWDJwLpCKwGk6ITp18PcY69
Rxx51E78oSpRvrlxKuSkfVqPrD3nG+/mxo7ug9ffD6siZqMrMKUFdg6WZRyGuvxN
zqvPvE0bvljF0lYG061EUb60u6F30u/Ui9yHhyIGGXbAS+cS+/ehy7bzFiAPnRmm
IA9pUQ8169fA4mdvuvFkOJgHYu62oU7x5oePe0095wyeoSQED77ZRoRKu6sJryL+
TUqE6aZk/lmvosCl/pHsMzDPemrITdtSNXsTc2j0Mw0FjdHGtZLUpyOV+Pnv/twf
71edcRz4OyN65CVRNZCU+5+lAptSlJHADbfzyTNikB0p81T9DTGUCjWO1Lfs/OVe
ZPUrW8hf5/RmRihUoYC1lg1rVMi2TT6ykVh6whn5F8wEH5Mf/7heJ6GLzEC/owAX
cXYgyf7PXHRvff4JQWN6DtsUYHLD+07R7AjgrC3QOMqRH/tTh6PIbbeggnFLdf5S
LW5amNJ51v6j/xXHS/A5SUN+vQ0SpN63NW9PFYn17789lT6lhRsmbfkhgHOZoDPh
e67L8+4ZwBuDdgftdn8kXmaG9DeL8Hy8Y3BnnlLbAZHU4GNrZAWiV+i0bg8jCLXX
GY/bvXZcd/ratomvBSNjP9MNV7WQS/0n7qrX4TfjasGTLdgERbixHvsR2YRBgU7T
XAatP0sxZvHJRheKiPzf0afkW5DmLWXwOUcPZzxj8iZ8CEKJ7e9BcXP9/QhqRpI1
c/Gvva/TqHmoYu1zER/9TmYqcwTQGUMvLEJm0BXGMIf4MAjUufQBy9CKGSK6FrWY
EeO/9ouK8c25UuCwICVyNCYT2si5FyRZJaeDreDSTmIIR2CvKfNSo254sxQh9nJH
VHreYwwW8PZyFfAqojh0JL7PDtbdPfz8qCQf4Nl/KMszfu/hGV/3h8TR/ClEm2VX
JhNX3KKMTkq5tmqCdWaqfqPiAzoIvSJprIrsAfMz7zXB5FzHcWewH2jdvdH6NDKP
nFC95IWLlLEVBTWa7HOnIkMpXQtvmgIzydLbrgRXHi/Bv4br8OCdzZ2TForyOteh
yZw6FeSdyQ/K0DO+q0+JxTh2EpgE/KCss0/nX/y2FUIsIR57ZGfUTJmaTbAH3H+x
TY1wrM6adtgC2d/iMX0ffbmVI3nH5U3wrdt40T0K59xJtm+1QUJj4lC9qySuJxD7
lTspG7LFSIRkOdYyZBOVBaG64pz42C0WyvcKbi9EjyZOVGg6ToWlLaUGnFKiwxtS
I25spYGF3JlgKcw3T8hJo94XZyJACLtm4QvaEss3lUGZqXMUYglb7X3t5xDrpsaU
N60HTHEdq/tmldDdmUOCZJ2TvO06hyhA8aGFlp06Q5OTcKRG6Tsg2RLa8eAFhl7I
e9gOurQO275pcv4MK6dNzrPOYvuthyFqzrdJ8sgixRJZRYmyMabjSEUTAgpHiE1e
yOxuH9DQepzDMtU4+Ky1DC+/pQvaRiUTqatSBTL2azHcpGpNJq2t81/PXjQepdGy
173NEsAnFsHYzT0mJu6LuOEXewSzDxBa9jgak5xFxM621ke2nD4Zfd7ez5NH8KCg
FOjtiO5D+1tihS8b35rNAWnlKS5JywBORcnCxCEIIYduueE7p9JjPNsf5kOVIznV
LxoNqStduL/rlajK8RJAJZGZ1l+wflr8/1WA61EHGx9LzCLqhziYGXYaca9M6maV
x7dkJohUbGwH5niCHWZqj01ShkTZA4Sa0PxNMno4huY/swZZFDSf/iHctd2g6kj7
HbBL4Iv9SSvGupwimqLaxydLETn0A+uqDQshcXdcuoP/jkUWX2+0MQqWohZwPcWD
VBJtIzV6/vra+GUWhkygaF2KKDhh4Ya4iaK69/bHaq916v1hxPae1nhYrkkfY/m7
nOmOOQynjYkXs+mcFq3UVnhfyHL1KYe2wf3uk90rYkEUbzNp7ywQC5vixK2fb1PV
55vMXZSOvORorPg9S48CQLISYOFPMk87c2B62eLc5Dsdi8yFa1jJnSnBRXeFEiHG
1Pym/fqyICyAADIDBw2vL2KGYrfSjQJnFQUL4HnKDHm8AAHl4cEsFibW23LZVBBU
DZEHs5XDdV3acJzP8SwZbBy6kRpcYzZW5pjU5Yn1RUE5sjMdTnrbDKtAOwFxzjMz
ySFqciiQ+Sz7jzxd11azKV5S2oyjG8UTbb3QyEpefsnAXWF+xTpL81gsfDb+4To1
K92zGXVNUbDkcQnWS/Of4pUD+K+MCesBQeSlEZtT1OJqn8AAGGCCJ56igGUH7oXG
L07NXMeF6GqrVrnwW7GL1+YWNBnGqq6GKyQi+QeB78ZTF5abDJb1JxNaZs2nLaZC
N/Z4dmT6gMLY5BNhb1IbAT5k0zv02iiuQgfXaRhzPGyvv8gjzZx5OhbHj7Psia1w
ASqkJgrj8/YppK1AHg3q27tdkzriXWdZQbJKg96j7w39I+8WgAXK/wMgxY5qaX9N
1LzI73023TWhsNRplL0ti6RrVos8Ll1qpGAVlu8U49QkduaRZUddy3iQmUgD1SxB
fkx7aTM0AbkzwlOGJovfpS1Ph0ICmEKewFNrdxmxWB+uV3PU2qiQOG7T8VLR/zBV
RaTFDAxc+dz2KKqwfD7ZMaGo9ZAvfL+ZBhgT2NcWAB62FgT5ndGIMoeBHyyTFOe/
FJBU6CuEPmBUxFYKQbMUvvTNGgV2+NH1O2ONqZDmgEhlFvgzL1Vd5iRV71Mz9Aoy
0Qkn4QKb058DSwdWlLQFHMhpdzjWMUs93lnaiiPad1iF65r3GAu1LuWQbDPfrBQz
N8dgZXfnK0NUp7pmvnjy9+zkcchEgzi7VDnts7ieVjku7je3D9GXEPLJO2VmvvgE
AJdiUS0Bbjfk20j/KpcrZf2TDlv1sdiGVGhck4RGxcEXiQEC7C4EEJBv5GboJX4l
6ut27pNHH4Q4ufMb6AR+LO1BasVSTPY8BpcN8RkpspTYo63oQMAbfKcUPAN8r19g
ezEECKhczqsgZDpCDR9g5mVxrUv8Fxqg81tE2lwlfG/pZv5me4LYaMBVxcFozvnW
AfiSLV3Uuh4zHgQ1XGLVH6dbj+NT5dDAT24nimmTPJWt9KxwD8DDDste0sDqED8i
HfoRofAe+cvLbWhM2SOmOwPXp78B6wCJwJMiRWHUV7t9L/qV984RUDMVeEyuWNAB
soyioqKt4e7aLZqDF8ym5T3kMXKWjUDUO71XuCk53QouySmXruNv7H329yVre6y5
OCQ/GVRZLODLWvoeLB/GDtjzeO9KcaHdtZl8JgR3NBMMe9OBh7+MWoRj47aKqX5D
CRIkzqkEYynrKGdHyLn6tE+Hn66prDPX1sfGfS6DVvpeaqKjdAHzSmjXF2Yge6mP
OqNkKL4BQtHyZRrAR8C0SIh4d018+GnDh/BJe6TKK5ecz1CzdhhLfLO2eI9Ar2mK
n/FL269BnuujdREtUoPo9zb511KZfMkEvqTih8pxhQD/s77cKLpjmjiw0AyletO2
vi7Cv32S8eI8QW15YieHPlMlXkSIElHG7YPalnUqebhAwxPH/H2y4S9vTqvIqdJG
Ia+JERBYvs5m4IYxfbZ0i0i985Nze5KepeV/DsQ7+nGS2FHP6FJyXJupK4Ifw8gJ
98hj4Kdn26SSPPtuAIaTFrsLzQ3/+rJJo2/Rd8EU0FXZmaPfHxpfF8Dc0XgZBuao
e0nnBZkuGeCB66RFPazF8OTeVZkFvoC7IcU4PFTD+ubu0spowimuWyXUbmBWSu6O
Mx11ZqTgCAVC9UBJMQRxX0GP4PD1XUpasm8d4PCihzRuAwLWB6cWZ6n0K1i2sYwc
/U4djFwFpNB3VCDath2DRMYtnbQQdDwihuB+HPNkkAsaHPZ/toZuxIPzyQf9sVDj
I56oAUzu9pnAszowXLkhMBrqgchor71AELblxGv0x0OOo1Dwdbiu/DPhB15y32k1
SAMaVlR9W/CujJiuM1oCte05FENjsgNCq1K/ghA/gqiKN3ku9YpbeyGFuJYxZy5F
7yh04ObLJg8Xv/aMkIza5sf/hZ/sVpjaKLhNQJI+dGxz4AtIgj5+480JffsdsDwb
AEkXmUPA0/T7zXZyY3FN3M5f8MU7dDTXPy4EbLd84G5XRLr0Ft5xVEzv2NnMQYkg
9XidyyJHo/zq7uEyUI6O//pVrt5CDpbckcqlyY3UbsMvchlhy+G5gB4FPqQAPKDf
DZSR3S+89esTjsq2BYpgsAaKVL6EZtt5MH5qhMBtXtUdX6KG49cjrlxflOzUuG19
mROGAgEL5TYys/o1rIpCBdlUMbfL2oBbGlPDMCDuN/8GF8gpPhBSvurfYrKgUVba
dO9MWg0HkOAY++OXuj/VW+wpwXih8LkEKZhej4YZYrwyNTkwALOfRZQwSddCq6f1
kFQt6o+97BTFl7YEGuHxry+35PMqeELoOqDcC/B43BZMvarx+XfyXuG2ge0T6ddG
tLmk38s1IploXRRqtudkCYrJ3yVgt5FHpjdtbBn7pwEve2cNK+hxHnmAdzRIXN1h
1p6Kd5jCnZjccPzZ5UZn78xdwbiAgM/sKd/lYHArWZ0waOUcQru6ZKMAHhzwcT4q
gBmCJ5RvcsYw91t+4uKPsXVxogQKspRNDRVrbJXi9y6XUM9HqRXKdd/bPhYiR4IU
ei485df5PgaihAlL7Q0Y8kMeFfqeMno0yW9vIskYMJaKXcj7HbflHh+h9+PG+g/6
U8iVqjGKYxUAKKIMx1ba6V5vZz8/tCAp3iBeV/xvKRnBwK73G6BNHSBFfFxw0CxZ
Rl76ApRr2WVz7ROw29oH9R5va6C2md0JUcfbUC/NS6B1wMjon21xcgDy0Crmy9G6
D69YlZsea1e/u4pGiGRPjvbv1E1gi0I12PgL+nfWzvU2JabRM662m4zr3MXJI4QS
KkCrq2tf1POkHKpiMd8EQ7DNW8MLsxmr/RJGfRPs37/50Py/k26jKlAuvOpdxNu5
O7ko8H+7BL3TRTFsOAJSsoXWYqPqDIyBrnjlyq4vsOAPucerNvW8EcgghXu4iw0d
s0NAxQuygcOBe9y5RCxvVmI2jEHdC75UJW0O+Vi2tlJjzDKKtEjm/eXo9SrcRvvP
/dL9mKHVvbD7f2RhXKTikvXEUfHZzuD0Gc2gC8nR4fSDgvEC79ZdR7oQQOjBNXNW
XwgVrmutgYoBicHjfi33V2smKOW4YgxWjH/+woh6IcBBSYDAv8pi0eyhRfGBUizX
p0brSDxjNEPKcTTeMCyrQkzfgBT83U1SrT/Lt0/DDczDFaRQw6hDY60He5LYc0y3
eKzpUCaDREtSDdgOEr97nHmjG6+vjer1sR7fuq+OsWF875g35uy2THcVskoVLFV6
UL2cEABgrFrFDjQ7Sd9vtokPlvIq75QzAvdG6XfKkSTodXbzBnbHeQc1haZNe5ta
mBimFrNVkw6oiGn+Iso9OAY/YXJBEFkGDE/cnyP/FbOn/eaRp5WxaZb91ENuNyia
TDhP8IvbTYPTmc1aN0YkpmWxusyMuME4F50lfQ/JR1IJOGcsUH4DvjLAnyjL6gI8
euG4N+CdkxS3GyESwrAyRFGA7bS0j5VeAfL+ufggogcfiDN5eQFZRacxWJ6u/01o
y5IsUfXYuN6hWACxIfFr/gcgYW9feCp6hA7hFP07WRJr/ZH2cpv2n3VWOISCNDJ8
75V/4NKCibG6Epdd5DS1+9676cZ8QUO+bCmYKLXM+MuC2YDq59oIAnPkA2sWOnkh
jpD4NyVY7au/VK85dkl9R4K5d2fsV1NvtcS2rmNLefMGAEIyUWxD3+rHUrT3JSie
YAahuVFXu5pz813iJFJYbSl+s59Hghwy90nWjEg7c0CU79leFeam4fz49WDpxbdh
pmmpSIV7QBw+tUXonhfkCBl6ELY8FF/ZkkcX5NlzhnFi3RdOTGrK7FM+CrwJ0geY
1KLUyOSltJYocoxuDzC/3ZcWcVVqk4toYFPOzYFi3Udlb6mpO/u8EVIrQBQTU+sZ
IZhAT1RIRCdpMFR4jiHXgslkNRJ71E7TVtugrcDL4t+XeNptEdh2eAWXRyU+EkmQ
Hn40NCh9zbiuvXYx8+xN88IMBn6DosxWf1UY/M5WKb6aLAttofOLry9Bzia+KeeB
k1hmFiuhMiwt87pDN06p3kCVmb0YWLz2gpxAxPrL2u2YCvsoeRkQUGw4S0NSC1BO
TqOFppdYE9b0vjBIXi9rENTyvNKDlSl99uK8eRVtc9TwtcXJ3spsb4fhnO/VaFrk
d3t3FE0QW1cxp0aJhznJmbA8S3CnQpz229NQ4xT/NLXv9RgZmRqEYw4BImJETto/
jnxHcej5ro8tHPeV4ne0M6FjByH8QVwTP6LHGZ92XU9oI7nyH8Buz2Nl0vQmMW/a
QAli3hERUWOOTUP3d/dx98GHgCjc12jSLt5SpXW8El3ehmABknnZjNZMf2YbcavA
Nr1Wz3obxDeFQexst4X7b8M2zStsRpFDS3NKwXlt+p2n6Wu2NPCzH6EY81Hw2A5X
+dpRAVSXcuAVbaGxogVYNfIrU+H1vwqqDx04yhJ8JOCYJH+Q+eyR0z4i8nRDqLYX
4f+YtpMtpm5vRcntOtCRH18drm+TWQr35xTEq/V4nQ7lkUZ2KVxlc9aSJXOPsA9O
YPOy0LI6ftjnuLmTgVa/W/LepuKs0rj/1XmKsAICAviAlDvvTd1xYWr32apKhdRF
J3j2qZaa8T8QiiBfOquzvK4n2S7dkMRSgu4bGPoqyMLBKwHJYVrC4JrL+ls0KlR8
WVm08OMP7mhC8ofGDHlksrSj4pqgfk9EmkDsn3uVao7Arqsfy4zpl1ER7HfctN3A
HMhv80Hmto0JlqYuZ1w5WTlgDaJd9A8b9CbKg213G3yRIKDJ6HscEecP9q8aprbc
eGLE1WThKmUqmqYHPDJVij8G7jsdJzCiqdW7l9Pl3GrrhK6WAaZ/wXMgfLjYFGK0
uRxUeUiUptefT1aWWV54+euY8Mngbx2DRtDE1szTLwBYTdY9uYZ9wGRxH975lpp/
sqZMCgFgDX5c40fF+tBfCMlNsjN84hdxS32daCy6qynjQTZpGvl0KYb3TVP/T66N
xHoabWWZL93VpCy9WIdQsqOWc7ZVXtz6nCOh7cgLXbDWoORUqABao4qs6Bkxfsxs
5dnr45g3VjJ88wTzqx/LusziC7a2HiK4mVmfJ5nFDKiyI0MNIo86wwrGdxoGWqHW
dnU2NSlm8YJ/WGR4iDy4f1MJRjdXa6OjIGk4CSStS6QCT2UJpHdOlotHHrNH2UEC
Y+HoY3YGv8AmicctERd0tG1UzM9cb7eIU9RS/OuAx1/DqeoP38jiiNfWM45R+uSC
yxX6tr42t24KFv/KVYXZle4hhUf75AgCUSdZQmbsRpQtahBui8qNAiYDSBfoOyTc
rMJY7l6bZSAynZIigbeLM21CT8qLQBV4MzfLLyCIXwmfHtn4lXHPEm1d0T0Z9pjv
Lfwku9GbFZ3R48EU6JpxfGKJcQ1TrD+A/Yv4QCT2ibQ29pMLbv1nkEWDaRe9Rl58
+mO94Fr1RAvbvGMQ3vnwPiaYsOYeh4AnkCH1ZIQChFo37W6MNdnJ5NKej4kPTsLA
Njdm8Fot9HHPN5YFTq6aZg38e+H0nm9vn7hEiq+Q+0yzA2o/+XeTbLrZxYF5tBvg
kBTrCyQYtSAOVak2FYXp8vCRK4KrY/Sa5TyPJAWMHo+erCWqAKOHxVthVwVXqkeY
mP5zPiK4Ir36QHg28bp6/QKxHM4Tuc5pkCOspahNTu0jbNmz48YvUz6mfYM+78m8
yJKLHtI8iwp5Jbc2SnlKZhPDImNoE7TbKPxUH/oZEyxOmjcnzLr7CkLxB1b7YILa
TmD1NVLL1AVLHsK1cY5AG2vxnTX4BKOMHgI2ZDstIUhjsodYHU3oyXWcKebFdfGs
ebIIHq+R2WwYzVmQWbnYnSdFK3SVub7pld6yDvYKCONzEK8RIXxMJELeev3UJ4u7
YVz+jcz88RJ6p5SdIQcUl4lOup+8NfQ+9obVwVEOIFkjBMMLCv6fe3aVFhwamlPm
HmaOBiYV6j33aG7jHkhcNm1SJjgW2WOJ3aGaPLnSkWp7MJND1MsQcUQOhU2TgyQf
DovTf+KDtZU/klMFTgHk/EFMGpwBSuSlCGQYgadNKmraImnoqwtwuP1sMqFOzxp6
mcvMAA+vlC/eCz0jqTweB3cCoNZgLLidf2FXvjTE+h354fXE1NEiLQ4UA4uh9ukt
8OUupznC6Sxk5uLrl8VKGT226vY6jPbBxKJ98pwGiUHr2YoCNezTCGQJAZ/TlIpT
UpBlbmrQzvvdICifSOQ15kzpfU5Pl/0lepNoRMHHB8QsDOU5TJTfxLgOWARjQ077
yf5c548u5g8yu3LU7J5/qsk6oRSmyKp1pearxN7zZkqp4JzbaVk8OkbemfUuv5cg
JF6bPNdG1hUHY8LVi27UVbazI3ESVK3d7CxeXbgvRsGTIwTiFlOW0YhlEvJxiumM
OPiG+GDkZJZtCxGRl+lMgYaELMRYWiE8ge/H+V+hntpZYjLETiG71ZHmoetWyEmY
DW68Xo1/3RwUsg6qWiDglqU4bYfb8pQ9EpxfpmUFW+Uh2cUjWYVra+JKefBqStPP
q9+giYaW37tfW0PDQnlnrXep+IkTNhRBr5Q7jwrlq52ShCseajpwBln5l/zhYWcf
ivs9fVnrpOIpJBhvjmcXUkg0IU96b4mm6tsiq55HDvAcQ2QSBmQFnNPf184xRln3
h7TD6zM1Xj+6ImYtCrYuEcehTrzIEzXyFxGlml6rTwpOjFOw/Zx7G0+PS0gPx8y2
cPVLoyohvFTMzNdl5VO7RHOgehtQ0RdRvLFzuApGfoLR2SjE9DE4RAY+/YK0hyqo
WtGKJlCQz5JEcVAgFgjb/+jiWSzwyhD1NagL43vCmWuDapznpZTxFwhRL5r2/7xx
qt8oTlBnFhzWGfupA/iU+8jPhzSItpa8nW5F+j5CGAP5kHo6PpxIHF9WsRsOGo7S
EP5LvIFHWG2uKjIa8ifO0iWUaOR60aU0gyOKgQpjFGb4VrnaAeY0a8CAm5+dQkTP
uUeQFoz0G9UaplAl+uSux3gP1tQ1Biwef6m3BX32OBZdsOFRSrlvIxIHv4COAxrM
tl5rcB7QhytiGBlW6tRr91mXAKxA6TxI+nL5S1fUsFK79oNxtia3PZlRNFQyt9T2
fgOEZZLdyZhTZ/62ZZ/Rl7CCES19YtO8UQlsR4yhb/LbwnOflste68ekpLa0vfNC
nwYJsdqZO3Db+Gk6t1BcyKU1rhFb1ivpGhPix4lk0AHO4krOwQd094lRLyVJTvVl
eAmvSilH+mhyesTRb4WZO/xpqsChMlSMp9WfSUUAjTh0RdxaXxxqkb9JK9taOVqm
Vc3R/jDBWRJayDvDdUN3AiTw9Z2sCroKF6egLiMxIj2Fd89oo/hPm7va4riSyzxn
KQ4jTrLNwjlXzMbMJAjYasdOKAQQPEgQVXclsxbo+LUbnxoCBg5jCWd/8o4u+ERh
aQ+euvWmPSq+QsvJ3FyTtVzM1tDJr+16SOtPuVx36TdA1QMT+gtFg3FnPu8ctBP5
POd92JeRNDgbXkyha3R0sPNWb8MUXlfPa1a5/bxXstf22qcgt8Um5MDfek46GJ2V
DnZmgJBLXoGQU6AXBYgPem2ISUrQMKoFUnvOY/KhcQmJpMVsiU7rVVYbZMOXqpAi
sZ1jWLQ9OUcJ1dzeONEs38k6QkNBBLJo3mbhGbuLrPW4B5PSK1DourWeNNIPpP/n
16eB+gxsC9+EAG+BvdJ2ozrfmKWFPlmn6qsCQtAGR9mLHw9+rUeiQffDYD3M+/oO
s8+hhBGBsU89l5tlJopUHqWh9P7army+ukssalC3Dvlx+/OuqKfAcsEC/+lARSLc
xPGTrw8sMMgByR/xNy4nvlr2tZ+qmhFaMjAYIOXD+Iy+RLFnBgyP4wcJvTVqWfpE
nTYVwrpVlLFxxhUvwUO+qd6bIEfTbdKBz3RUM55JkqWsKo8UtNH/IcCk3pktk+Px
+YrOwbncN0olWw1MWGHolwBhcoedQ/cCsRsjbxRsvH03nrFpgbEob7V9NXDntaeA
2gl7xmqnvjV+jnslTn+j4f4y6ghiix2Gj06Ay3e1XoLHsCBgUbVQwmx0MND02E2Y
an7X251aoFCaB+ASwaMgU94ncrXvEgq3j02n9kCpMwI0g/T9GSu2sFc3WoaGko3V
GLoIdOmyEkDBg40uSzd3+k9C10NFFDzM/FHoJ1QDB9QdlkB51JX+muuQWqtchXO7
Gl8FytjkSqVmFzjyktlm8HugaBvvSLVVPJhpG6wFniCxlYCgDCJHkdXCjvtUWcHx
7JC5t5R3e1/Ql15pZ+8syACY46KDjZ4oSTShXoWxS7LptJxeRV4Wmp4llZsKrEs7
jb1e5QVhQWT1qtVNDcBcP0w5AAz4eYVydLUHsdWyxUyY8SLrpVnWRhZMrEz2zzAo
mXfBVP7Sy51Dj+I+t5Uewo3BNj1DxoFkWYg5kdQ0t23XY73B5En0otUnyZm5R7r1
CibmZihiNoZ8YiXdm1ALCtJ0TNWGsMI/XM7rVzMCnlFF/yTl1AVwBaswGynoCPPT
bgq1VCJ0l5hyu9tBV5vAdbFC8xnup23i9DYToZDXSB3R6npq1hbGXHbhYLEadzG2
Kdo/h4tLFcsmmi8mYJzbMLKhVtFjfiWKzhQ2Ahzcb2EszeBrawfzU/yElcC6yJ9E
j4fK4P8bkOETC7tz6QGfUsz4tm8EZkmFtFNcfpYCwcHLi04YK7rhSGJItIBEK5a7
R1Dj7jCWOZAuCgME3rTWvNKnD8arYkMo9Y1Thx7pLhC0m2fg+yt3Dc8U0nk628UH
MHIVfFszkh+ylK3pMt89258VvbHUtGbPBxRwrDXXnOP2pvLGy4JUrNofa51ak7yl
piOs1N5rx0tTVBSfd5u3ZHv7NFiLt650FXRdn7JJTpZDEwTGOmEBXFW5L2AhM7zK
2wM7G6+26JTTIovFcxDijenDJ8Bu8f7Crq4cLiG8TPzFBFmiXhqkXrQ91gLbwe7I
R+n1D4RrFmYNFHxihuOjND3b0bCDCZqRm/gfJdZLn0Qd3hAqteC+eHXKzcrkVCdo
NcpE7/SgqjTBbzdt+IcDkDOIWGKlpn/FQh48u5TJmMRt9lbOK4F4uNc9+Xx1bqwi
a+bZqasMINrNZhwNNcRtuJmNXkc9ocj89XfJ8b+ZrwkGISBN6yFDdJl1/5CXrtxT
PJQ4WYM0vEvLikgzWA8BhBPATMrGf0LugDY3ClmeneyVV2CsX+uSmg0Yz0u23env
qEx4P1wFdlrum0aaDoM/6L8RafKpjD7LViS8430CrJPJ0YpQJONpRJQTb23zfp3f
p5zonigIBWDznOAW6kmuapdgqlVdttVsnt9EUXz683JObAhJN4LtXZlr/LWUe7ir
gaXgJ434yUCkIxzPYA+WW5lPghZO5wBdO/Z0iRdKrVQ/7Tfe7jBm4gVBrxeMPliY
FenFCdKFztcf3JnRMaOFPdAUIsjammWA28MbgtynKd5YGV9lVRSfW70Pp+7zScvJ
c+oVo5uDgET10q0z2FnpfbYoUH2hfzGP04mN+imWdl2kX+RvbkUGFC3shkDwHAw6
7kYYR9K10C2aNxCq/3jog4+Kt2FgKe2CGPtbCMc4954n2Xcv1t74q7vDzmsmbwHO
nMOJsM4fv5zX0MyBMw8hmXjCdkAzKn1yT/eUAPf9XJ8S0feQ9vPkubB6Zr/YT5N4
dbD14k2taLO0EHpp3K0LiEQA0zTMP23U5QcEHYswBo8YwVuJeWcNIIFu/A1lBOUL
lKfQEPO4z4SGcFN0/ND06EtGjMS+A9CVoNzq61SMOkV2llNuniaL1lrS2y7sVwUo
cOuXsn5MHkyUlSlpH39rPDy0leJWO6asDcSIIb64y/nPB8Th5r4Y7QPKnHqBRKsz
BNsBbKYaVf0zijbJ0JMJWxdC0h/8nce8JEOzZAELCXSOTK+gneJiB8FpYkNcXa75
Y8MpZgSiyF9ndNg8DpciTxpV8nONLn64Omz6ACXDZCtjsftbMjSa1Koij5aEheOw
IdLF7OCSYIY1gmbv8I+mHeywq2Zml+6PIdn5Oylg9ITi0xVVJcgPiiOn50mdaBic
n/uu4gsszp6MblEhD4GkV5MjVmHIEBPDqPGccr+lfhA5EC/4rJun/omQPX12LBIl
EuL1K+qxM/JIRWNKzJIeUJ0v+BpAs9yUWrdJ0sU2JZq5mR849hqDDnjPqipHkQ0v
HhPJ4HDlG7SSWzKRd57lAW68RRyTQ4yyfvpbY5rJ++m1m/o0xRU6GcLLlCqDI7E1
QS70P6vw6zDWIgeMJzWe6GCLWNAs7QHPlQcGl7J82TH7WNe7LCmjZCfKO9chixGQ
6up9/bRwpZW1FhJqFe+0xn+uZF5i7tmF+4iDLT20W1skFmZrJI5L4RP9+FAe3wUL
jqIZjhyk+cJgn6eQY3g8fo7kVmUz8pKBFfwEmvzhXpx6P0Fk+9pUATMF1A4suH1g
j95Lg2t1ERqu3ZBqL5+OE4on3K6XzBnDkZTRE8Ej4iTZ5TixkFVtFLs7kJnSyn10
wlqt7Keb2nyGFlINZ6tGFvgeRPamuraJRsJU+NoJUdbak/RYwQX12nusb4Cfz5QK
HLdmAp+2Qm0RlgP4zbqzpKtEpblMbwIb2pI3OqmBV3HuILFgsKZH7SzFaVMGBJ5a
kMxcJguTD542k2OzCbOQuwz6VIlD9FZpO7vJaE1Os8QH+s2MGY40RE9dPno54BTN
IPdsb9FXozJX+LaD6DHO2o0pUF9I9wp1utCNvWAkaYtH45RoPgbFMoPKqiVGpndG
SmHaSP9Z4nGgQoAIub5m5zhOn2y86fossWtdDxeBTgmjEflkZGj46qDfj0fGDdMI
Vk7W2qyKFAF/TGjZrpriaRPNxZ1qHGRh/ucKkNqVZ0+C7rj80onFmecCMATr8hGW
cZ5fr4LPUZen8V7mIiH4cwG9KfmJzraNJreU5S8Vi13ROVVuXVc5CmMYJSgGxD3g
J+4QwKg6/qPh2qKvRCP5ln/yQ7tViPPa7+gLg4pSSK2UTt3TWEfgCTu9LkP7bfM3
CG7uT26BGDUSnaWS2879ih4sYDG6tbRaDSn4N/yMmwoTGGMZgtHcKApRQ4sHYy82
wvAzOD8lEta0fslktOWJduLcc4wDEP7rXU+iBXx0Naw=
`protect END_PROTECTED
