`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hcKXhJDZayIND5NAIfzVevpJKzIcVNXg//QaOwRS/kcKj40lMG2Hvk1DZawfiRcK
qWhMbMtIY8Cli+vjNfLWpCL2RIMtLo22IRETrwpdDYj8u8bkJrVhuEOnbKSgMPLV
YJ3IVpDf7jpBKKZRr1nST9jMJW0i9vW04qVzfiMDSJ+zgqYAQmavtWIwX20bqpBV
oHkVFGqmm1rUGMFgqbP6HuW93KEmR27uNFm/pI9abhTm/gDy5FbUaD1+BoR6mJXL
C9DAXwG2JZFi4a91BM68VPgZXez04IlK3+SlJAUhF9pwPEMrTCycCpJN8bsoX4p7
2TO1Zere7Q2ThmRFtSiVv4vBUH4Z+t27fogplQ7ezFOKRWnenQKJItPDfTADdRQU
y3BAXj+0NQxLNGnCPuywNWBdVEW1O2gjIzEeAfk7GhOFKuy6jjdiXgBIemHyARcR
TSS+Ho+W4hBiDQwQFglcNMmJ5/FeYm9y7HVZ6YKy43WGt8UJc7b0AsAv4yDXzged
4HSY3K4YHhnVD8DNj08mOA6KcXRB2d15I682g4+i6i4v1qa+MYY6JZEm+3BJd5HH
`protect END_PROTECTED
