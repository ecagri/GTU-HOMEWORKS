`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
00yPq1tdFtUp2BN7FKzHmPPz9eqi4TC/ytiY9827IokeAo/xks+La2bddL8RUi8T
smQWh2gkH2x1wcN1Gdh7wP7qtB6skrTkdA5/mLyk79isCKLIB+zOWaNBB0AFYhnN
iWPqqJ0fDBrqYFx2l+z5UXKKmZTJHByiEKUiZC5qoeflFYeHgsb2HdOIJgj5xNhd
6gZb/XwnMwLD/9Bss382dViW7+j8Ns5HMqWkdFyBRv/wlXDbB+DgxwN4tDZRLowf
PXMWQPN4wHv1jqxjqqXDRBrb6rA0QJmG1wImcv+TlOzyZA+XiO46nPvqFT6YlSNF
sr7cpaJdJFanw8ovs1lhQ4opsOEaAMpLTy4FNconddlLyYzaPOtc+UU06n96b+eY
0ywh3AdziYAQV/Bavt8EO6sWuqeE2xLEIaNN29Z4FLcn/dyTgWp68VUVCfCSLzei
2Nwlqy3u9Zo/m8TQYYSRHfIsL8ss5JJez21qcsAqy7Ilvd6pZd0USVxy04VQyR22
ML1ZaXh0GRsUEHNcMlbRHdJ1f2NZaxrM8mH6GzhHaS0/VHe9Xqb4rITNA7p7aVa+
IXvQ3uYya+QFSlZ0aQRYnqPsqivry2BHKZT6MdNNFmprrFo9LnUohQ779FvrrOzF
A8LSX7qQ1wuBvrgqXCRIPTYAR7yh2mUnBiu9Sfzhg/Bi6Hs6QhAJ/LWYgN49i1b1
Xnw2dZeXVj1mOtgwz5VuhlwVFxhHSMJJnxtEwQcIMzOHggyxVUVxkWML6TmWTyy+
qoXxMca8dORXGyato+8Jo7MULZm9YgtqiEfl3xVdNroZnBoWX7fxdFUonGQ9qeSV
/1pWxJEnHE/Ze/ePgJ1mRP2+/DOsil9+XEYBs90mwpsHeUqJPH/ME0jPJrlyeqBk
38xoa5bmvXJ7ypz2TGnQlxODzGabc2BMoNL2HgbCjrgIFVhv7GMXT07WNVfs4UwD
O7cDwowbFFmXziOzEv5riczRuatfZM1VS9NhnuUPzTqM9+h08IHK160zlq7Wmdu7
x+aUmcRkYUULPABno9yZtOzo7IxyMtcJURfp4L5yXoZ842UMqn6l5diV7sRNN1Wj
TcfLDE14QELH4QcNhAY1pWy6iyMu2vAHBGs+zgzez8ehtrUzR1OXUF1IYFBGOv9B
7p0HLHlcRBBSHqtrw1WNTbGIhSBpPQc9cIOBdDkZhhGKUuYubDNZjOS2ksNzT6sa
vXPvEhBH8EZqaj0mMNWzTrUCCEVuhB6aUdCeFnbO27icU4HiRX+rpN5AHYibPJyp
qOD++kqJxghT1Xvc/TMyZKK1I0hvr1B9L7SyO7wwlP4sJZsY7wwpVA0vTs0v4bSw
Mq7pGsQpY/7TE6Pb/ICQ7SMIVu+8bAbbajs+vI8AM71idaCWRU+pcVklXUn4MBSR
2LaNWg8AEpIYLFeWXhFKkcJbgYaYdoN6/jF5qOVupO/DOQL5Q+NQE7kvCzLubTpp
zXSIBfcNqeyDjhZ2sZQsrE5Xf07YliCTc7JPrsDGZFV0k7qw9RbbPSRncxxFikQ8
AmINvMsOVSVwx+Lh/Xzcp0dqyg/MuiZ6MSj0JLg7OcU/c+wIAAQdYgUuk7tjF076
8QrAuwJgeV+zJ1ArSoVfpP3PI1cQk9t0WwDqrwLoq1reTQ/E06+DXsYNLKGr0Wi5
XagKaZxA6LBF3L7XO5QlHx0chjH+qPiapfIKBPhXXw4QOTIGjGB/3zuB61N4l2A+
+TOoT5VkZWEeVA4Q0Rkxu/ob/A5JS9+xvgR2T948Ky6LdqHjqiT/CyFWQJNDr/nf
jw4Oc43dHXObzFjvT1TxmjKJRvJ5Aqmk6W7QFIIEw9kmFknMQ5SDyeUoxkUOa0cI
Xw+AcPpN6AY+K9xf6g+Y4pVB6iOItQnPLaONIkKmnB/RdVg4TAXopNwYoIjYZPfD
X/SH13LaDZgxTCNrl9WUtpX4vNrzu1X/OInMyVS69P92HWLLjCGdsYGxEc5d+3Wk
W7Zw2K4tw2tLlzYXrNIRhBsO2HwB7ZR0/h5ZyPiiTWc5zO+0PeVJaIubvsl/D4VM
UPSOpSCXnMJHQEpaJPEAZDBHo+aeRC1Nsueudmi54v/WvbVLt3kWNfJBG6gV6w3U
xA5koxao77l9ShiI6z9vXxWAe751hploeB3R5Q0CBnc/QnKAXjik1n7FuFTC/G5c
qje+ZyttXogOp1dyiS48yskzBpdIB8EUMiu9kMF6zVyQdpP/y504EbfR6AiVI0tG
lu24xDCFFSV4KVHRLNeTo+zY0/qKpDL2t5EJMSSY6V09AoYvxOfggRjlePnF+h2e
TJPDJP8K2a3UeM9mVgAhR1SLoiYcGkkZE2vDJo+m7XAPOFxd8mfa8FBQ4eiWVufs
0/elFDIzJMaQyD61qr1HfSnlKakPkGCZZLPeEXgjL8XYOBNcRS1cR7jS+ijIu5Ki
8D3jjr9XijbFbtYAuSpiSoV7XKUdtol0cjGI2hAQ3+fGNxoqZcVoXCaunkE8D6je
nzzY0W28S2hS3lrvIXmNEgWjU0v8TSriJL11u6s7OziRcOhNTfOlpdEG5iF6t0UF
IDP/PQnbb1LFOH2lfceUsu91S92roc/67i7jJ+sHol30Adv6xTnI0RZ6L0ePk0Vc
BUuJABChPcLoAh7fRV4fYtZ2gFBqLxzL+W9qkICsS6kgjeC+gKHo1Zpd7q9t9o7m
2f4I2tXZzqpMqQwhkYuL79mQ9zO/CIdALBiqr0t0KwhDd8StP/mf/EVY0j8zFWMp
nWZmZscwBbh1iRrnFUCfteturjqk5R1aZ9I43GbGAd1LsHouzHj+HigsMzyx0TJ9
qkoOjyiq8uYeS0GK6yfxEW000XW2UaZXPYs0QUym8D5jGDtZIbnCUSrRj0VW/WlA
Feuxq0mb5JJB3BarftOLNTt4F4BrvAwfYrSItPz+NGhoVHBQC06Rnp3pRYXZiT6+
3jkMHgx1RFDqacaXdqiCJnOY8k/HDVo2uK6E2KJpXbXNLncqiJAsGueBsaKuZzLB
T4yMMgpjm107wXNgaae1o3exy9dZId2uJEeOpJBvwl2QzD0OFrVwC3ZwcvNDRAZ4
9Rdv0cRnJYsaBnJGUx+dHrSL0eCHkH7XGkVa+vThPo9kWEOIwggVZ0IcPnEJ+Oox
XMn8Uxrls+0u5rbNNOLAdZLL95n+BRlgUFWUQSWBTXITViWGNzgQSQDiW+qHCkUW
5Dol6rrTFYlZGwl6lk7jgULHrGsrSP9FokvlctJGpa/IiLbCrTr+Z67nxxhPkUQr
XNhC2VPKmTChZ6/hxPHOsSFUs7Os5dtxsMasdSUZTSjtI0APWewnOzr6pOTrUo91
L/A6wBQsZmP6TvhCCADym7VAwOa1jCTwzIie44sl4VAJyiQWvXwlBuiR74vSyIPm
hFsR7MXWTIMg+HJRS0oXCm6IataEzCLBeVvBdAk+nuHWZ4/yNsY0ap0vx8bAO12D
Jyr5wud6lPbg9Gr8xaNs7vk7XP0PIkgfBxogiZUKClf3oyux40SA+pXDdclGYSlq
OlBgF8U+VjxrHk0Aid/tYBuxdUr0JLSfbwJ1bqcytsTnCfHd3tLevsnTfpMFaJx/
A8aXl4UMpXFrEJJTMLROI9i2effCkVkXQs5GHvJT0MqlsgqkCSoiqC7mWysn6x4O
ZzMGfEC+W8qboPlv0dCyHVUasNExuwIFlSkmNnsdpuAcJ4J3j2HtZZ2/G0TjiCcq
E2fpFa+FIs+JptASscCAmRGLx1zAOS/f4daAqbR9GTUQks1zcU1OOaKPRskWR9ZC
JCRvLbiF2qEwLjgWNS5Ii0W1eX7admkXLadj2fmaWyRfrDMH9pGuvXeMUeMz0tUv
1b4b/DCNWsyeA8xe7BmvAdaKmAFiM38//EXLd3Ba0Tgiyu6O0vDpSrbX2GjA7x4P
PhcgftB9t79sB7ldblIqm8+zHBKMaGu7/txC4Q518Az9BED17QoNqla3U+g4+nzU
R/cCmN7nQrj6XEefVkqSMkblwgLNazr6a/rCi+wRYWKGjerH4ugvniULAdrGFGp8
ivt4ie2s8fmY6mTNSJcldNVq4Bucn+1liLG6Q8FHLk4WnqyrX4AqmCisCIxjLRmj
B+JtSZKUG9TvExM5yUrAnAaAD96euyQvlcZaLgoJdnEOD+IqP7GHmMMPbJTSBhO8
X3w5U0vRc651K8rQKMgD3LnDTOb684vU/CdSu3KivEFZhuNrazqykccz03RTXcnS
6cgPE1JK2Dcwz/kTVqMjqFhgnSnEcIEuZWZ7IGTC8ZAxzBZ0TLLVolbHpqxX1q8S
sRj6+6Qxm262eV3YbpVChC012JVicQFJZXVJRnq1TMkmOXpCFlOVSD/LL+P4kpIV
q2eW0zH8TX2HZu4MCXcLcu7XsShiT6sGjIKerQrfwLcTqBIgwge/A0GAekanpfnp
aqBtCms6HMgezAZOdqeOC8fg9YP+4HGg/1VXNo9vgFS2wJP3ckv4rysFebHtyGa7
9eJxbCKCavU57fDT7MwbGAPOzBn2B1AhBHqMJf4gdIqXcfgnZwD+0ZofwjMkruLs
J17IjI6ksHf7x85nRm0tYx3C2721exavoNmHT4cWeaen/N9/ay4l2GNVZfcn3vrF
5quZH5uNX3UprdSIqNafsC7FmV3b//ryTdYQ/ew2RzEI0Zpl2JareRk7L04ZvXRg
jm8O8U9I/jL4sQbeODq1yLHNeBqFFDbetV3PCTArpKWeBPTuj4gUSOxo7qJ2DMVc
6aqOcfQGGzh4lkRXFjI7VQ6gZOdYG8culP9we26NbnkqocfIvURYQ5DfBA6lrytE
Uk6QQyxLEc5MKAw/HAve8MISOCDxD71QiTtdOv6tnYLxcyMm7R2uLNvSCnUEvG0K
x2sgInbw2lRsJhAYBfjlo78S+GXX8+CqCEACLao2Pk+WGu/yMCmJQlrgP/vtjvOf
YhEUjjS/et0vpbZFXcPCwTO/EhqjSYGigJg5zt2An+452TZfZbF4xkxMclQ2CT3w
2ICVN2KbRPxfHbNZOxOZpnYyE/2cLKGzpECBO/B+eb97yvhq0DzKRuMiabmVec5A
QVk5PNILTfvxYbDu4/+zBZt1qEHrI/XuCdLnVLC8zDey49Uhsr9hiw+pum5WhAO4
AaxltmZL59bbOkAZowHpJPW1wNUBruobNE/tg3fcb+AQnMNV2FUspweoaPbllvof
+/+NCHpUYql/3ty3ytXZ2YJZQvQJjSGNAXXZXkfl9a4mF+wzCV1R2/UFKvuJTRMI
tCjU49g4tG014oC8PMVU02CdmXf4BG5PNOY+SUbAO3MStahyo5KgB0gLOfdeRAei
UuxClr9iKnfYYJiVVLFHfMkHFqlLNHmcDM/zYS7jUNz1ZX5pRjRCjWVreWDvF1Qe
yySn/7DY1S3n6wNGFC423O/NUUrvDA/o7UYYaGenKms3GPoejBZUJ2tAPoDHyL2t
VrPuykold+mp4Al2Y2CfmEW0Uu+9VcdCeK42qzv3uqGA42UsreNx1rk7ROQ+LGqd
5o98aMJPccbrSRW615iuZ3p8Bvs4v7LC6QpMbwuLXpctjUzzeK+BmjlxdGTIEPXK
QBGGhupoyiERBAV7s5UVs4jDjao5eFEeTKwXDOFIAe/L1ouo5X6L28tNI6YAM59J
8A/UloKv/Rm2xkOmDcUgJEInzDNPsQIlY48NXD1btvTzNYsZM6S0rNWKxLfsUTV5
5x/J1aeZyBjh4B6RBIJkX58jM4v15cUIcON2sIFtgUsGkc/qWXUvYwkxcsp9U3fz
flvKbLdkPL+MLG57EHuJ5Q4YLKjwEj5ZhvNze8SyMcMEroarrg3mWPO3c0kG6oYn
FmsTFPzyPRs/6UyEq5AiKqc/WBR9wax7Xjn1reNtoQDS07HuCo7ElBq/oELvgywE
05pg/HePgz6BFS39OJgu4EYHkZ0LmMpx3xROvpUyghpZPgTE9ttwq/hVkCLgR+MI
2iqPejHUEATe5BiKJU0stJ0dtJgePYG19RYd+wl5qjEVlGLZWZbGGq1FCBCLYkIa
4Ce87BXk1tCUvQBjzjqooY9kLQvAG4JdQZC+KdDy1p5ICDBiPkJSPeO84TK1Vj5r
sjE9tOT3IhOyq+qUgfd3WXEbOPR+MtwX6JU/3FhncGLrsZh8EzDtsovzR6wqgi36
P3dWhrPY3YiicBTBNOPAvQO8h7lmUR+0AhtEgxQg41TFgN3Ji8odq+akOHyX4wX8
P496a9/Bkn9/LYIkWpfq2p5CRkGz5df7AuH0648+6wbhJ69D5Nm0rqiI4dzcsBID
921q1m7P+BE62OgjI6XpoAlnaGwzfVRYIdq2R7Bx+wXkTucUL1ErkgFGuWOY0kVb
CiFxlrt21MT1ZX+JotRxczoSq9navLwlmldUA4KnjEpPgjQ9v2sR/H+obayVj/8L
SFsqM0EnyoWzruFV8X3BdH+w+Y9o2gH5duwV9cpD3SmRAx8y39xJlx5QlNozLNpN
AY20ybE7TgM69pDM+xhSn1+Qj5zFrHTdv5t4ThEvG1Q+NK4K8LB9gAzTbE5RrPe0
tn/rDQuuDEErQdySSdX+UgbF7zXblNwwl13IkZHDr6B6Ivo+oW5phBAPUtMZRvGT
FOfqyk6KXiSKR7iE28qj7zVn4mo+oUkgZTYqK34uTTqRwdg5/S9SJ6GdLp1oswHR
UYfJLb7MFD3HHvUYQYz5L+N+ItXFtcihBDvCfMoj97IYrPRlkAY5XmcFv88YaDlN
w6QH0kaJnVv/0XebJAm8NUNdHj7KruuNDgoR/9GXZjQEvOB551Vqf6r5g1FNwbHi
m/+bxIWtsgJthtj2h1DouGLJrcW7We1kccbL6w9sehiQcdEYG6Pl4XuUmGQQlbEK
Q/h4ZFr4luhGCigLwAYyjuzWDM2ZMSDph3qNeXP0i1A8Vtiiq+wQM/OdiFVE0p68
M6IBod0hh6FoPVSOYnnZsm7bw9UYtHnW8xr4BQFO/KAUBmruEw6SynZ4Ei8arNVc
yhW9nKkYc1laXJ16MBJxkgCU7wH8Z3yKzPwBm97uoEuFUAAjE50aLawWigdrB4Ks
uLNQdnWxVB51KBdKfDEi1DucQlPICgJzqNTuekj50jQgHwmQSbPtm+O2hj6ldEbW
0KR+f7FWnzb01JcfcqVjRkmWQR81SPIhA7KDfuB9uMo6oUkEVYSifL5qn3SEGfp2
UTWPEgse/Z6c0gdpZ8uVmPIJUc+QV6ko1q3eO2wUjh6SEQV5IH8vPDI04kpB3lsw
rop1da3tQ9Hu7KpELucooMIIB5geq7Xr1RkmLpYDHVcQDz6Sjqvv7s+zi1oC/FDO
AZv+EDqEw8OynWGlHlZPPl2GLNNop5z8adqfuRPG4LmMbT68vBqvsr5q9xmJ3cSP
ntmig2NtPFnXjL1H6IumMcEl6HOpOohQCHYwtG38L3Ehm9/gpGXJfYAvNAVxnqR+
Rm//AMzvsjl1nWhApUni5IfOSXSNAEUJnirAjUYfy+NtRbiJt/T4mUiIX9slaTz8
SH691bcJVWsdenYw2zwFkW5PyE+ooDAxcXlfcz3PFz2hNWcEkJ8isN70wjC4LMNJ
lH40UZPFpQYKFKPx3DRkK8icpivmCjhFkQrfhHbN/WOhZvrCpAwvQ2iN+/mR1Fpi
QT+Zwme1rWkd2Isi7HswZ25XJTKsrsb4CvPn0vDG1JPGZfeKU+0VhFf5Ke9Z3pPZ
tz3Jo/n/Mya0dvV12vgd50iNcCYlx4QnKe8SpvzmOzIfIqVR8M6GQ1IKBjBZXDhY
AM6T+JI8tYdb9IcUrdn5xhSG9KQJtaeB2dBzMMQsG6NzQH+xyTJYxKbX7UByqVMM
ZaxbjHlCcEc0hObTVlBPzW8P+BiqXdq/oxmzhRveOKIXoZkgdoyFTrNeNTaLGu1N
zsU90aFy2rOSqJ1ddLu6PPaLwmEYru9cWBRNm+NgEnxjhz2j6IHjcR7yKl0o1Lzz
LxO7T7xTI1NkyP7RS5qmAxA2jOz66UrPz6LEapQWS4osDpF9/JpgbEfpKsK6rXV/
2fYGdovijmqpCO7bp63MUcHp9wSDCgrwNWmGyv+nzMILKIFG4N2r5LyBaKOa/MCi
rWir5z3yF15CaxFjcdd08m70h0xyrh4vMZPLlLL/XLNUAeLl67OSRjEP9I3aHEi9
X4xgxYDz6LMFosc+XOUkKMJMMqZas0WiqqPR1RaP1sKL67wlPSwKQR7iapgeq5xw
rYul5AMmpPbMBdMdo7G11pvxGEZ5Hqig8dd9xydtcootvQT70jQIQYEwMIKn3TZp
CR1omDWPfzxNTkF7MMn3G0KA7EWdCLb2D9kMzWsIvTaR2VPYGV6gfFEsVfGD+wEz
x/FX64t7nwYNRNu1+xacgTxYtHC+OGv8XmkMpbK2CjSJRO0eYAVAA5wAa7YuWgQy
b/4HUN5T/ixRZsrL6Xipx16BxZBeKKNNFB0XrSrOU/IIIfaFz7WA5cVJaQxjNWXk
/1t/Jq8ZsYOVk+HG/kW/RIx6NVcPCA+oqhtddYMYH3fTfGO/CidBQhgS4U2BYkud
rZ1r+jkVRMJ9FJZnCzTZxV8uQ9bstVSBW+Nt/sHMGt4PGUOPP7LdxdhAAOhbs8AX
3ARx1ph9M0sKP3zs0nkH5vkjWkBqHy1M6m/+e0d0AqTM9N2QvaOnTzxkFrbalSdE
J6cf3jedxx2qmnvt07KXP7vyDLdLGaOBCQiZDQZ9oWsCszKQVcErFAmb3P4jsniY
UJq9uKfwMACJoW3wdmsIeZdtu5bckt+A5pm9LjbdMJey8vGIqd6il3s45B3+xFYu
8UovLJy52iJgtmnixWJ34/6YYDLb6DhtxscEL3JREQU7WikLYDsRG66CV1MJ/Ng6
iVs2lpHfbia+040I5ydajzIyGROPfos8tPXq4ImzibFqZyVr2a7fMWRaVELv0tQ4
JnJ3VhsYHsFLkUcGoATND2/uzWSWjBNBRaLEfppBt5TmBj1qOzt+Zs6z+8FCcejF
POlKLzIEJsKtz5CaVvU5rZp8Ze3w6CqfkeU3IDZnJtiJuyR8Wx3iGXUid0oFyMZU
c7XQTFKkUuSb6Bt+MB4y4QR2zeUInp7gLhZgb49R12oogMZpGsnurWPIO3QJmf0e
VQzi6cN8trF9Os79bkAAg0GO9qZ0CpIIEbyk6RgzmUEURbbdttVqXTgn/HE6h73J
u0BIEAl1W+2dmVSqK8EllPig2afZq4FYH9Rs5djVVEf7YrQ/JjvhaqdQhlyjjfBI
kxi3bL1Npa6/YBar3j0sjpAqxJgoVvsfnq4zsvb3Qam5L8cvsSL+kbbTzs1J53jk
hCY+4nLB2l88p+eJgXDwdk5lytLKq3o9ZDFVdaJDe0y2ie4sE51Bhk29lYzFyNg1
p7YuqSuwsoT5Afw5Nt252Qi9mOdakQnmf0L7C35pF4SiCyyg1d02ihHp32L+KcuA
e/kameX7PKf/MsWWuJkP4pnx3BADPCtiOHfVEcD/y1X/E6PAbgRV38GCDetYuhLp
5jDbJYzi36nqIrSNWbmRv7gk3y87i2IlsJgTJZ8D5OMw89FP0bZhoBF75O5RmhRV
9I4Hhqnh7chgxLOylD1Qkqnh0BhCHnJwCK+TQ+slYbNCSf5ZWaErAzWxhJN9oK2c
fpsRymW1pEu8ItMywVx6mM2lOUjwm3epdtPZeMfUpdALmWA5bYCeLisd5t0+LJuC
C0+V4YdV90Jo4KJ3VBwvHEiFMSeRP87o4ZEb9fut6KNAXhioZ8XD7BKLAdIsIIMU
fffJ6siCKvG6diol3k2ksooEAkmU2+v97mrDOhrDtJ9bWuITsTcfA1vHQVyKW/5M
vaZz5jt4cDsl4s6uw/QZAnxKjZ5Tj6+37KjLHft09aHwKaC9/DhZChWxqQub2DyN
53bGQKVHSZRVEpdlTY/PnaQV3Dp9uMufLPTRctviZ8p7cXGBGrBxnqxjDFQMdmf7
/8d3/icJiuhshWQELDWxHm+DWyxuSWBr06jBgTTR4/ZdnU7nwi/Hi/d/YE78lqG7
xhV0c8/wiE+9Gg4OBXoVh/YzwttbRmHuB2dV+WSKyW39rJik2wjzYIT0Oyo1QFhg
nY7cT1+rMJNtE1ENn2Aesepf48HfUhJ4Q4LYcuqYZg4xIFRKBufFZVwi1B/VTm22
IKsgcxZnv86g55UXwnz7hArloYfeukMOpOuDNZakXDl5dpT/hVGB+okPwv3pGjJo
YuYs3Znnbs7yYLINmtXkvx232itfZMO3bXcXzGmn4lZbABBX0ysDxK9dv5xURemz
sP4oXO8kU92Y7/22EzX6Sg+6TquZc83f31N8uHM3QAO8YziSEijs0FB62a++Etn9
kt5CG+xNhPL7572MEHhs+BBqKwXPPILu/LMFJHuCp2y3D3Z2zgwNGroZqSRbHAqD
vpT7IdQmyOD/2UpLyJXCbj6XFj3lvNos7morQ1aJ+wgZqboblzUWQ8DlHOVDQ4c3
bVi9RfCe/BDnZc/+NMBnTi0L2KOGvsbNvtrtb4xAErrDXuXVVAqoFPRcXJ9DHNtG
LShAdnV5FdCmrkmWyqeNKQotbzYjaYHnKWGi46FKJ3LRmEhf7t6eSzevkSjXuncO
i9Pdwtn5UjfzgqjeglqWAjld/BJjdCNTKmKnMazF+IlYGMS+cOXxMv9Dumruoisd
K7jwo+QPkOasN23qN8uMl4pbr5o2zGgysNWRqbnTWciCFMFc9OHqm7AP1ua1wrrK
ytoBi0H7nhr7QcwAKZ0JtVLqk57PNM5chF5V+odWapEWSxYqoiT9Q+pvYlwGrw9D
A65QQjSme+F7otrLsgdZthO7DVpiLVdSlJOAr4xDe0za74L6DXympQ0XSm334LVE
tC/u1rnFK7b1GS3zYWOlPLbDP46Xo9RFNwc528ge/1mJpzl+blmcpbNWFizmpyd3
UmlZH4o3ADuRUUOU4AYRSqV6mVwyOqsQZsTw/NM4Vxz4LUSChh6b/erwrTha6oYu
GT8f7VMfVhs4in0xw6HXUBBI/t+RGkOVi29U0nIhAQRpysJjeLBHt0yuB8fqrj9r
qMvMNwpcFIrK/Kluc4idqxEae6Okhm+u7ZVrVKkQV+WUuzwXrGS9vZOFqaArcgr3
L2yNs+Gd+XVYDiwG6t5s4XII114e7dCWEdkHkrtJ+kazgph9hOcYH040GYIgVG/M
BnJgv04dpWQ6GO5I1gqq+TReWWW0sfEfObDXzRgFFMDT8epSAp0JCpWVore2Zlxk
Mn0gDFGo/sryW3y8Cx9XDByn8a19VTZPZ9jxiGD99rFnugUTX5mcCufNU3D2bRYK
lOnt34/q0y6iC5hXY0SUMMLmKem0RsACV6raxX5I/wCZ+TfFIWEaNF/pLqj3LEUu
7KQpu3RGZm7zdpfKNHHtVOJ5kH97eQEPOlJTjEdvXfwCOWpaGdyRbzVvfMpX/Lv2
LNL/CsCuzNBdzkjOjxgUh+eynMTaRexxxfwbuFiUzinTOjRm49sc6T01jPWUgxCd
2rkOkzyF+cDepyU6GTcRT0NOO5JkU+d2uOXKZOEaBKgwNJJmTk9E4e+rQzWw4shL
YIDF3zUiuCR41nSe4uXMHv2rJmJb5YwVXM560kg1sbqmjijxRQDxraILY+ey9oCo
SnqVBDCOrtd4I/7FuLw3IiVY9n26JapYER9fvFJgTj/IO4qjNLRNXAEWnwmRMQYt
rVMScSjIArLcaXygFL1HnZlA/fOXzswUE0VUB3YF0ZBsP1ajkZv3ekSM8iTAVWoX
AP5dyFpu/QGWO+yVgmkwa2HDkj6VLJWF+hRRAsmxwxb3TFj3aYRz+m8b1iWKXqdN
Qo0r50l1CKtOcuIaxQWPdGFjx5kmT5PMT3QZmD6ilyE4ybpSwUpWI5XycsZpFveI
8pOn0dxw2buwX3A77qLhee5eM22KO+Gm2bO3jND0Ji33Ms6q00/Hw7iFGMTBIO4L
mKipN0MdpKJX3oMhDXOhwQ612v+SAbHHerRONp23AH+fCFpW/EbS32vTuw/KxteD
IxzyQO0cShFMht5XYbIekOv1vuvGMdCY2jGMh+kao57dVbKvLTV8JZLOZxgpn1w/
IeKfCGwX3NTVjZu2X76n/0XbpXefy1NpRX7yWX8Ch6dFJFaKth9CLDSJ1YJ9EYn/
TOI6ynCVeh0O9JQYddp0l98wbmJ9V+I2NNvduVp09DrEfL+S5DsOGPAiLFo/gNQT
4+Dl819MejjouWoXqRjvj+OiuUz4yE6zpc/HI9+RMkwEO4cEjYAZ1jPjYwSZqmLO
F2AFkF00pgr0JCJpAdjBqx2IaUMLB41VhRG9OsSIQHRkvy9ILVhY4aZPJllzNRJC
ofRbIMvwr1ShCVGeJ42xQjMNeJ45zJqlMl7W8ZXc0w5kehT+JLLtTDVVibM2XFC7
DTqI24j57aZjmjGMAvzwqf1nRtDuAFyom8jeowsFmdI3ZnILS5UyEdKgVBWt9Vs4
3nziYbSJP3SmcWviPk3EahUZmyO5EqRyEjHqTizU5l3Q7j8jvF2cidSjiZlRTig7
PiwfPwLnKCeRf+Mg0jAuYmvfhFMGVTJIBSeeENP9rC5jNdByKfL0nzLQTKVd8dw+
X/v+m9XAEsbtCDZ3aTcbJqZXN5YPqtsW/xj81ciMtx/R2WeA+gaZ3E1nMwB+ocyq
pdAnEQmyieLZDC07svtnoVq7veynKVULZbDHg5LajJ8vIuxK+bJUubEBf17nksUW
00Xc3PhGTXH+SZRsC4rZcZpC9/y0gD2ui7/jSmPyCVHS8gZRgsRwTf5b/YqJynUa
sEKRpZDo3irOWo0J55KtqHoWvGqjbT9M1STkzNXXyNXRqXC+BR3jCzH4RH8L+p1N
J64G15GrOzT31K3eFwZEjTivVEm+aK3Q1oVfGVqAuuZO01gqlp+MrBEyRwxzZScp
A3N2ePVQ94nS0/CmcaNcxGrwSOZpm/ztfuXQrmc8DH85evy/Lk8Wqk0SMtkKBi27
`protect END_PROTECTED
