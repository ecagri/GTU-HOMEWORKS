`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zwUWx6WTS6+t1MbfjoPHQ3ZMNs2Ho1l2VJkVjqIXS9mDCXqtJk2+Fv/EcTtJxB+L
1rJTamSZx2t/guIq15LyX9iEJaZ9xNHK7wzSmbi60spkJL4aHIc1xq8UsI5aLMZD
DtRasr99mNkNvup53Eg+uY9R7VQX5mXuiFI+3P0stsalCRSsEehuXtJhb82QRpA2
yhDESH7XCY0B4DvOBb+gRbbGGn6GQwbhpXS/hZK5mTbBuNAOXLuud1rhuMXzPZZm
eo6x1+jxfKBh9iILQy55OAVjnsNR+MO2eb3G6MRENGrNo+AwKIe4g0hLJgoFo6fU
Rp989wqn1msHvhkkdRyfePL3CxmDbgXu8NIVpuTaOsYawFmijsNRKUD5V6CrG6M6
Nsny2FY1k8tbpZy0+o+AEP0ombWJ+kLyN3Fb3Kn4nsmjKpUfjnF3yi+Lt1Wa5WWO
shjR2Vrs8QObWXDmwKPnPJEUrgj94SNwFDl496ZiXX1/MViXleclaOi26NZVWkDL
++uQc2Iy80+oX2JjFXVk3csihDWU0XsHVIq4H8NWYS3iixhiwGCVGrJZ1vxk//iV
qv5nleKUTQsBdWKFFm9878Io3sA5EDfFT76RU3SMdKjLT4hnNSs06hxqh9ra+uNL
MYyMgj27fXz6Y8WSfxjd+sFq0TdGFJOM9UPQRhjwdno96n2IsTiS2VqZAtqDNGTn
BUQqohJ4pZDqwqsRqs5XyDBIOwzIGZC2aXzejHsMnBbGsWwhKqLhqwW/8+mH8Nyh
VbHP8LAy9Y879SXZJTyJNTjv82mtyiFU6LKktkJ/cfw+pWkUiwoVizzTDe0VfNtW
/u0Gn8eWkd6Cxer1SN5eO8TM22MbKtBq/mvvxGdQcAoZdy20TwcWhg0HnYRkpFDL
`protect END_PROTECTED
