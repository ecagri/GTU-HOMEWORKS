`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I0gbhvommpsK1AJyfMPh6MluvnixVe5cr35i/+RkjsYL07rm8qi7nMqg0b48ldZ4
nJmcnoIECZx19RTLyuMFDzpII0g7oMX7DnczNkTmMT9XipGAeHht4S9JxufvvDpp
/7QvaVIyiEvxgkZVQK/PQ58Mm/Pcg6F2/zUGEQ42XK7chmYwqBD41oVcShnGK7vP
AR06pG94nXpsbpoJq2qvxiEhfDv7kmMBn9kTOUF/fHXR+ipLAsywjymr6n8ThvMW
rja0VwqC/Go30bzShxLxGAeqWq/Z0WDMbhgc8J51OCocoFX33pmygFlUhBSvxW/D
ypJtkumKmwGt6hTRheA6bekHPApjC9rHooI3uzhsHafIP1mPIZ18EMYeFLs6crnf
KNp+BetHZ/J1UFI0DOBywWgq6fwM9GyFxhdwoeSfgmoMJJCbJwYd5DnXmXlxvRhu
Gt5Y3o4dpefC2QjwpYOnhfPcsz9kHarT9ZA9bgAnXZzDoIJQOu+L0A03sUSLMZQh
LyUad1vRb3LDpD2bBdj/fc+IzNA/To4lzKvZ5oXVqWOycBO6tkC7QyQ3GYtJxv6C
vkLRMVzYW6m4xdHiuoPv6w9sXTi1HlI1uXHuYpTTu3AD5mqROxFHK/RC9SG3e5OK
bZERERfm6FOrCgLNnXcVNAwgVGFDf51uA2qMQcRnZ1OrdlUkbUgbLov0+qRgxJAl
9YL39jdg0oNbf41Hx2xXfMfnve24hWaOUFvaEIjBAwmrECh7A0uVPfslGD92B7Hj
YU9L3XD/3aXTKg6c/DNMAodyYYznhIhPpZFJHUDhpyCUEY5DbZrI7uFCxgnmHseB
zXjiC+DHEDuil8MtVaL1yVc4kiewePEBHPcu9evOXS2e/q1ARqGIf7L97pNctK2z
zPJjfbWMCOBzepoYn6p97FzOB4t3xKmXbc4rdoc7jVuRi3RO5T/XdohWmLgRef5g
OEBGophTw7ETYsdmbAOVvXGCmoHRDbPdizjbJg/h+t8+hhX6xVoJZactrI55qGh/
s09yDusV5JKPcY9RsRM/oT6m27UDNP7+K0kpkzJk+c8DLSacOFSRYigDqcRqDupU
72rOLhs8+Gh95gojsgMe7T15UCfk+FDnGmMJJJ3teNUqjt7mr/tA2lNBkcQcW+6L
Erpv1Xfzi7FBUFzXGUCSbt/+4i+2Kejhj32e2G7Os800QFibtKe56cYeLlKCnpSB
mOEU7uEDB2h+sJ47jZFH2Eq9gASChXSDUzBJcQuuvMIJ2U3FB+vYazcJTrbKjjev
EuHOMs1eMi/r9+LI9RZ0Cm2lLYHqmCR9IwSWaM1Fhy+p/WlZb00+FAF5CgpdwpQy
SLBE15fXf3mu57f9fTXKNi75TQSUXA3X0hhPk2CPlZWJzbefqt6NSN1bW+mCud3q
hLXJ9WOJMcXhC+glr4NcmIEEpWlrj1+4tGh7x/gu3kah3FmOn8gkPqbkHpOupXPZ
bF6UchDJmS3ey45E/pRfY+lfhzvp5Aq9yNosPJfym8FuUlKt0YC23tofiap3AAhE
i+YTegTYHHmHCnwP0bFCzWUGkNr/ie/fkxorVyn6ztJfRUw1dKnMOATLo1U+qP1R
atUO8/I3a0tZfHl8j38j3km9/ZuJilSImE4hqnTHwSQ9MZ/6ktRAZX2Ng+gmB5IV
hJP4kH849Vr1MN2l3BHmwnmdhoxUB0Qctm3aunCPQ9fXeBpuu35TDeczKi9ZEyDt
IWwruKmZAu/EtLwDn0G89wXDZ7AXvZ1/v7pI42jhx1cMROJfuw36ZlO9bPSQdKRl
8d77b+CBbzTb//csxiCYGPm3eL1jChuWe6/FrTkaO1catl4qUuG4fwbsfYTOJUl5
mxebMQ3NIV1dFNQTbS+VJ6RP4RR2QD11PRJq/Pg6V+k2fLVVA6nFGoX+/g24wfqY
6HQfeb4qIcFo+qNzaxxsOT2o34afflRND/YpTNUYvgd6eI2Mp3AcbXDEFANgrEeJ
XECmBQpzbIGGkmVFVbemujpCeHHIA2rrKwT7PCsuRcWzyBfDdkPDiIjUodcfVWGq
4IlQDHzlvP4vVtagYVaReQ5wA6ubU+CKQs+lYRFklMy8o+qoa/Ttrmrfnvb44Jfd
opF1sXWlCfFzsadNcBJat0zwPr+1WR6uTdXZqEpBinoNEy9LKrpgcRI7zKEFFPq0
Mmh6PPbF6AavgO/FgyoKP5EFULqnoLdlOdxQDayJwlxFLXQRcgs9Jix7TVZmFz3B
+pl1HCoGVpriHMjHZu4Qm+q6+s03dlJc1711ujcmBr2XQAA674qQVZTsbVTqkvrt
m+nUv45T7TcAcvKFNsC4dkZRnmyYr21rAwURp65qQLpS73PEak5e9fUhDnCE6yc6
kaLsYNtnASGS+i1Bpis3Ps4ZolnGIijeCIjADbmSFNNG6DHd5hRuUi/Q4vkScfsK
UZtxG6MHQCC6jUFAg4Mg2QBOMXgadjCEnrzFKKSSkGtX5HFE4zDlt/Wh8NYtjJUj
5NOnmbAu8UoVeSkgkIRQ3QQnQqKXToNvZObcLzdBbzNcp7HMnTyDBAOO50yLPIXi
8rDNYgWJLQpHd1RwUoCJ+I1GoScVwhAHqtdltgxgS8c9mY3MYSnaOYWPdMzgr8B8
RpcS9wn6no+ERrnzy0xu3wPW99ZTZgevIR+b3T3NihSsFzxtGvnk2ZnnaUSvFlnn
GgTjt7qoOnZFWxVMNK1dItIzwH8/qrkmYyeDk+BIj/qMjAqWn2yX7NVSsNlAARYE
82+94x8CQ/ImYTqA0l+HnJyVS5HfN8M1KNpeCQg8x4MlOLBq05Dyr7WqP9A63wmM
g0SuerryHAYyfBWDjBAaiKmy2HA7WInoILkYt5Uyb315Q/WxLBPprXV2TGUcamaN
fns726D2ts1d5Sti/U940kwU5olx+MCfA2cQk8DThnktYmmaKiyYx6FW/2J6MmWq
X3vv105xOVRugYqGXblM9aRd5BJ52zew99LGcX1kTZZSCx9LWSgviYGBK6ZpWlT5
YgzCvhrbXAKOd8qp2JM6SYXCatN4S0EfpsJ1pHs9DtdVY8GfjxaK1R6fv3gDh+DB
GvE/nCsygiD89eejAXZ9Bq9N5jEPV+JLCMRIYWnFocH+tiN1pkLc5o5rGRauy6dR
dL3E57tnxZ75uuDB/a50DeyUVij4vhsfBJaUGGHxbtYVVAqKdzXbGYrN0RtSZlOK
zF/1mTpsteeNHYOHk/inK+OO1+ZGOW0/aXls0U0dcxScBBSyfDZxBOixirfF5qk8
djcGoijUssOwUYYc82QZjHY2UMRZDKiSkR9aacP8Jrx97mcTRJYlKvMY/QJHIv1B
rJJGWFc46tXii0IfYJF52134St36YCHkZFZDiIpcAFfFM2ILP/9qiXeDsbi2WddW
a/WU0YRJqi10HmAplqP08Y6bVxwyUqudF0V7eTM3RsFt75KT4pmt94nUFCcD9E5A
Av9uC0Po5dUz6n6fMSsjGpn+PUgQHFXAZ/MXI0i+o79ck2GBHKySd6dVP35e8XzT
xmqv88+yOXUBgFN77j33zDUyMQE7aA9Ik4EoB2xJGgwWesiyujXNdv6yShLiAx8G
kupaV92bRC5dgAUZVwMFz5d1CFccu+JasPk8nHproAg9PxNVx8VaIauORwpNyKsQ
NGnVpwIqlmQsLza68/gtmGNYF/5EYXJGMpMJ5qei+j6hWBaZfr9gHvbKA0YksOcT
0BXUv6kRtVu3G638iC7OVYZ3ksNaM4VX0HH7uM1KzTLurf0iATbROt9a1aNP5HaA
vBD/KU184Wxo4onz2Y2Pu32LfFve/KqJx51wTY/gtH9j1Rwcsay+STl5/owNOgXp
tkr5LVAmad5GatHJiJzW5PWwDcYvOFOIwlTXy4/4EDcKm0acD5zyjbedE0swEzD7
YVYoQLLnIcMalR7T9Xh7ANpbxwRuVaR9mhYCdVzaymF4OGekVChy9opgBLMvprnw
pbXfMZ+AtySMpzHogRKNez6z0Bnj9CrwbVeGoQEyjao=
`protect END_PROTECTED
