`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I9s7AkIw77rTC7II1G2xAZzKK4JCmgsyN1POOx/KyPFj8u6IkqEj73MZrAqrAM9D
Tp5gbZW9D1G+rKCGNsLlj9qDfjaaOvH50WgtS0XN1lo0hlnJyMIZaxL7uS58yc2L
eViVyeipYqsKoXFcPmMjupEAzXY7gcs4csOk87bBUUpTwzBz8ADeT78mPoro1R64
UtleZu93d9XSW60I6s4otC18I4LVWA+2wQ1zJUvJCjUhFR2tQRVPsah6faYORu3a
mk7PEhziR55i86QT1WpuXyJs64XtnmBZ3w42WNZpkdyaaZSEYBtU7+nffrOpuCIm
2M4NHjN9xv5BHiqRgnHE18rdLESsrHG+H6/V0OCbX9mOCHDMI1Pbeo9ArsKlLrGt
ahOpwO+eIui2bpVSaMGORVXgLFNMqDTdlqyjzGxQxnfWgJHoTCWrAVd5TM6aQdH6
/9qSAqniIiY7qZgnjkTOkTL9q7pFvuDN7BCdRPup1H2GtIbvZFdYLQZVl5cq/tSp
hvU4cHyVYDygR8W00JuXhA==
`protect END_PROTECTED
