`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wMpQMTh7cuun0HV91p6be6GiavoUnh/DqPUL8j+wwr9QjOUvpyBEVQY1vUSVM56z
KNmQDp86/lpqgAjLt7aNPawM73B8T00K7fXi3vvIg0qhazY64cpDUZlZUTm9gejr
M+a24dh0AfDgZcDCwwVEEhRNUolrncUC9tLV0gztQg6FclLJ3mjF8uy6RNrCfGvf
KPNU68SHcsV5bUcPK8yyGGuJ+pIUORF+YmmSwNZf91Bz/IWCqkyGxOtztZ3nhrQw
P0sgwdW7qzFgANzAP6KPkPKMZtoQO+RFQTX++e+zf/KiW3/sArOXlGwNduI0KGsz
ylO0ucznmWmWCJPXAnbsj5aOHakPkjXZ8BtAYaDBp5FrPYJva3p8oaEovFjXjofO
PmZU4MZGXdQnlUBwsF0Y7nOx6+FW3WG3FLUbL/2iEizGJ5WAp6k7kjMSB6vryrNj
x2PAoblckV44WVAy9CKCd5yS7VzzU+9Byya2+4yLhPnIzz+6o4NHmtK/PEbFAyYS
9QKuK7KJJBHc3XrjL10HnEtTwO/McX20GqIEEkUoFIn0a8LFjyKeua3ZGLTh0yBG
xRWeHFOXzIFbuCQJ9ZgJtMomdcm4z2x7bmoVn4oYHSQF7TZwuHULEh4JorcY8HQJ
fWnWN0G9hQe969iTQIW+ByyeIz4fuIj6PlUn+FGzGeMr3POos7q5ZZL0D7GnDyUG
+sQN6X65iysi25PIswdXDSaOFW+1GZ/6xYYxNZTRzB4bAZDiCGA88vTPtDAzbINw
RhYtx6nnZJL+Be1Js+t5y6QB73SooOx13vgqDYkbnAlPKLC5lkng0xY5qw3BaAEi
oSWKDHJi9luGy08jiJSPuiLc05HK6XH+13xBt3EZGeCGPjXnd7cuSeq/MOEMJHcT
k0YZgYbPyu8adpPQta73Nlx6C8GURRyFQ1W5BVnYZg5V/W2SHDbnDncrWOLkK+VC
CjquRHTcOH6KVIZ4TZp/NAvnuj1sLBHxNqeVInfXznJwmR6TjYNodb6sv7S8H6Id
2y6LxqCL+EciIQpI/zLv8u4EybkXP5flYAYBg7OBS7tfA7zoaTwdi6Q8xD7qvQAs
2WcdAf77gOAZj5xvQDkXjvruxJfIHQxhpSy1NupXzezutQw3QlTTRMjigwVtuGDz
zTMfZTNcjcSNwgc7HWrSHOxWVJp27d9NBBMPSIB1cCmrXXP98ad9CAO9J+Z8kM7d
jQwzYe0NNl5iI9FdKl2dZOE4G6X4oyDycA2GxfkKrkpNJc21trHtu88l94WP80y+
BsJZ6yuxHl57wLZYK6D+sujGEcc+NaF++cBnlRq69CCyGNFU7n5x8qduc8yoTiqW
11Ib02jotP/kg7FG+7LE1uFAW+NOxyWxolVIkMZlPJgD8YR0UQAC9yh+Mw27kSmD
L4DAxlPDh0A2aJAJfVfZNzhyom0/cCbFSIWkPktx5FJvkKcSFt1ZOeDoAL2yxzNO
NV+1hvX5uiMtd8q8wlCNO0NfladuRJZxMVQ7bRT51sxd5pBrkElXYRW4wRYIQxVa
3Qq9EtJLz9oswHVOTozQujJhsUIhH0mCrMfFcY61wEBaDKVlDKw557EEjpdgt9mx
WHDMEl39LgROtnmvNDW5KWltfKe+okCkX4aEH8wQFqWMtMYzZBqFVEArSUXOpmyV
ko0TrLJPSrksTzbUB50xDweKL7c0ToNUT+/zck/qhjQknA2nYTa4ZfO7Gw1YHtJy
XiSEKv0DBPcfL1V37FJMqh5VNJopwxiOQTQPVsTk5kH3KGX1dhN4XOa5RMG3S/7e
GrHOzT6GnNU0OCTU8/vEqO+7x99FSOrBITc/AeMejTrnCrOWdQl+kDclOHyl4+7+
hSO2KanryFiBdU3jtWBPHT2tnX+PCMPnEACnAx/Giq7lUWlHvF1ODhPm06infAmL
FUSswD7O6ipjuv9ZHAWluoInyj7C8ixGFvQkyEFJN6UU+dGdtRwvMW7IB9xNiQZQ
7mZpCVQl+hXyDmcP3CRxTlMIce44TLRe/RAONo5mWbKX9WAZkXf4vpCCf3z92oyC
C+J3I7S//q0eXIokj9GWzd4XNy9ou28TkFss8EQ3C5+hIMglcR9k7qsoeRPr+UdW
GuK2I12rmZnGNnMUTcEWWtXORIPJMLe1iaAuQswMy+9Qn/hOlfGKqAbRQ+EgUBiy
fBDOhzEW6FjttxJ9zAY82HYjOA9tY5gHUbwF9ow16DJHyWOin4T+HGGLaf6LP3L0
9LZKR/SaETEjiqnnmTDrPejXvyy+xIWxhnuKr9niFydRDAQ1CZAY9PvL+ORqNfg5
IvcnZR4QjeQZGiU3YVDBeKwHlrUvdEIWcIPG3PQjHwfkTFcgCJvHbdVprdN0Rx4r
C7EzvI0vFb1eTIj0hCSPB1SYezIWNzs9f08gJQfxbVIQQdIbx4KhyITL7r4648Yv
U/GPXL5dSe42FxjYrnopxLXfeceouDrpPTD6KSvyDGKI+k/Uz1x/n86XcYsy3AB5
LFaVgIwSBqF+AIteyYzgegmal0XoE4e+YKWK7OIE+1pgHDG2SReBip18vp0FeWY2
wsZH31wjP+Kqz+prIt89/j0gc9ygqMtW+mr72lVSXCSp5ZQ/1vNWR0GEU5UZ25Mp
kgGYg5KNjPuLzG9+skn7y5LkkLk0ZWkwkySAheIWjjOJaeepUYDx3X+BZsuCv2Co
A5ztOIc+2C9rbJ336RQRXKbLqkczKuda2pR4OI8VFDOvvhKcvjqE3bzVzYFnxCZ0
mslJFwoMPqBHExh39HYqS4R8sMR6flKlI781gzXTiDee4ti/zUnERlRjD6kFsLv8
at+1T0G66vC3uoqwu0gN86hErp8mYmXYmsyVZK+yCE4Uy9DyX6JABU7dYbi6RkqL
3qi3bXrtqYjwS2eKcFRk4MBcLVaWjlTrm1S+UQChxXUEa+LgGFRQzAjtEykCi6r3
g3Zq3mJsEWzEypnf6FvoMzx09hQGrCOTKb+E8G4yumagfNZptSOQkOnh6gR4ZWw1
Hazdjg3dcOE6ofvfPvjhaXN5RD06FURoPPzbGPInCnaXI74Qw0JuEhvYiimHEJD4
kkxPyNhKg/s4YAe0CxB1x8DV8tmC1VR/Jl8poNHOcSwhwRg3+VJdo839KcS5vk5/
hWsvsmb+55t34M/VPQs6NTlbw8ab1lWqUpU66CLUmHmibp11WXNf63pRzarL9EDS
5W2G5f3EE2yPKh8Fwm6KzK32br9n2rzXt1rzypSfm607+5LHKGy7/g6+w0Rxk2Hx
H/JRrFYHy3SsrQWAc/l+9PHNbGSrTKfqRNImQk71d423KM+B0QT8be3D8rXagvIL
sLKkqW4bTBQ3S0agu6vk8Cmgfzv6DHpI+l471ArlcCNJPPVY0ZjLWlmSSmkjUBIL
+ReXXww0O0DuTYqnIeB3dQuW00HcvDYvnm1HX8BzQktv9Dgpdps7WSWPEwlJVQ34
gKiVN2j1tgqT7bHzktixaytjLzynYk8WBzG8OTXXTAwknmp3G90c/Lc2pqYNNPm3
f7ecpQuYq9Nnp4Hknmva1+7+Xv8dgw1ydc9Pakxfz19D/ZQB23a9UgnYxI1VTpdZ
x9WT9bQMkxjAmXUZsRP60Rk9BkJjK9oo+BTMARzVU4EKVayW2J1SA6gGtjdmzxH6
Ntsh6dXbJexNjwHBaK9jGvK3jjYY43+UoLFYvmMxO3oEZDMnaCHUU77LJ7qiZCZL
OBJBoiuRaX8BB5K/yWMb8ZQjpUstYmLhdZZg3xbcQtsZYAo6BA/462oJOclv5OlK
k73URStp0pxyv3yMW60vEdWSE+2xsLfPmgA5W6suHGbfmDI5NJGLYvEkcqX2ViIQ
VHJyN4+4+dEaxvubux/1JnnwOrOkL+tT7ZtNH+KBE0YVtd8KKM/SxOcPtFeetO3N
1AYQHCUcmI8nRgDYouSqExxHvPdUFeHuvtv8rkILLWL4yajjNlLctFo9NB39RTtg
OFdItAhh1L0OgFYt/DaUVdCv8Vscb0NpfrZDySo8zARdtZJpMry7wPmPfDI0qlDS
/de0JJweMefPW/Q2tqzqqeTAn2fUXkrOgG67f4dGqx2c34f1TejpcvVYXAUC7Ojz
ilQZ8lGmiQLkGIuibECmTs3y8mC0Aw1kRz47pRBvfATnWDMvMlgt7CtNoqCS4UwG
V4MxWxGDzIMS1d70EOx0Rv2JLEngA7f3iiYSsbl29JBbHSaiys5kUlV82JwDbF6W
tV8gyk77Va4MtDSSpe5YY+DyGE44kSlXKJ1OpNUuD9y8oP6+5xjHrRyxNNW9VJzN
6Uute0q0K52L78IsbC8Lv5gAERdhrbUcmK+nY0G+cyQCA2HH93DJE21LELFoRvvj
T8IcLo8X9RzDRyj7UXPedgxDnLjPApDyn5cmlGi/ZCf9UO0Xr8ZjSSkBE7f12gpc
9od8T789ic6yIj1fD2wtCinLMouilSWv2rmdZ9iozB4KCXn7rtJzYV582EuwVINS
5Wle79a40tYDaUXvAhCobfTMfQrx8qMvT8J2frTT3Qt7tsgw6VO6YvK7xi22JySB
AgtE/IppOZajpM7tjAPCZZKAAMJkK+qBorccH8Ah+Np8lVNZCzlUhgoaz7HJfxm2
yw/LUPqx48luCXY4Zw9Ztok9T1Lwl5cGghDgoaRr4scrBEFzI7lC6ppOu3W2TO8c
gPfMwZCXE36hD9WYJZQbAXcJfCg/YLtB6NfjoFaMUs77mIn/qA/9EFiFGV7/2BdU
Sakp+waBBbzrCmuCDUMtmJ9Srs8ZSSS1ZLZHq4Y87yDaLhzpAYkSeuOsJU/UOs+O
OFrXFn7sGDrDj6276KBWTHhBwLTSg1dr20b3IoW8Oo1de64Tu+qDIF0eDuisfhGL
B8csxWEC3met+TWmiqqqC0THL02RnIM47BxF3YbWyHsl/Of6/EJvEnB/e4XdnZSt
OD2GOI50mPIwvgx5F20gxcpfcE+VLNForP2kyfMHQbIxHO28DIa9uGFpI6a5UFr4
pQRtmfbKmDOcMwP++YRuIUsr39IkBREyVjO3raoibHyfOvhsBJp3KpaxxINerb+w
07mBkT3vu1+O4zIegzlk78JLqMYpLVG/htMoShAGOx4KlkiL0sDPsSJ/btJZ+vb2
uH90wXFbvVtX0a0yHT7Sgekc30VYj9NqS3upQKNEaxYb0bkuprT4GAohZSao+jHD
/4gMKtnMezeFD1c2UkaYYqnL9BkXVzABZVu+dab0lSFQukH94mrY7CCYtFp62VgW
E+k/fQI9Se1PtDR23ONC78yxEXH2W6gA5sUM/mPfeOgxSshzMK4OWbTT0GUE+b08
nVBJkgAN26LHr6B2Kg67bxOt58KyWfo7lNPHLT8mO2Wz6CPfTQRNeNoqT6rTF4T2
1GmdwQgKKM9gWMEpR9qLCjRAXNNt35vilLxsgTB1ILtFEwFf5N3bnjVZyZqfzsap
sutU2bw1DTPFtIy54Rm5hqxTiyxUVW7IRLcvvU0JxDIH4zjyElKaGLN7W3pmZZcf
quzQQs1le+35iuoq+IbkYIZvhZeEz/cxe/JpY/YzHbq5Aql4gaCHrN+36NeQaZZf
lgpV8g6XDLJhOjF0NolHl+luuFCH4X9LqEA35fBMHdSlnVu2jnV3MHlA0I252J1m
dXJEDeaSUqnvLtia9JF0gl3Uj/gL6lw8Gqi3ZsF2zn1SZwMh18cwW8pf9oToU2RK
D6S3OWyio9uOFPvVOmzgGp2e43nfVyqVGD1IQmuja+Lz9/LUNLmcNizE1oWiZL5H
N5ZN7v9pPZECUKVLIFtuxrV19d6Fw30fDqkqdasYA3cNdiJ8crsbxxHzw362dRA4
+OVM+kbO5uKz862vAtIrZ2LkhdhT/Yx5i1k3Lg+Ixnk5UgyGxFsmCow00ELSK5VN
tONExXxgK5/CMRSRVQ4IVjV+iYhVQnNw3BAJ5OwTLVupeKLy+HlufVyvISxFPmin
KBCl/4/yP2Z4jo/Ee7ajkE1JO/0CU7BhaszgUGb6yFJgcfZTAUEse6KRsggzQ5aF
K1JCbYlFOJvqzPN4mxGgjcqGZ55ofgnqj9Z6kJnfshtF2n0cDVvrm6QJ8LYMa5Ed
Tx4YsUBF1cqbiPrUk7VQ85sRb1hlspYuyoskZD6m7AySExIu4dGyKa8nRL+G86UC
m9BrV5xWZgTi4+bciZ59cHMHLMC7YHDZLPZ4jwgSY7K8LJytEBqL57nOhZLONdbP
UN/5mEPpQHckTlDBs3ZFyrpk0FxlmT9lBkF01RFu0Q522Uu924qJ3X/2bSXyW/87
KbtcyCmxFNOGPqC+lJM8vjw5ntPesGxMTQhKEgGXFWN5ASWMbwREXR5K8n+mPDPQ
4zrccQgRHhVUp6HXVLDVZVbmHZbbagAqGPNv6QSbGPtNvv7IhHL/4DqKa4Un5649
fZk6NlXwuMU80I86J9eCtW5+bVBwZFP2gPoVyTpWujYQtijLi73wRO2elWmV2Vgo
d4fRYLh0o60zflkCbST0jc114mQSQJtOcH3jRGbhK09mU5PwjxIcSB702cpV1G3Y
J2PdxoOd8sTC6QEVQore9EYzx0LHdvuZL2YrsRAkwOo5D+htLc3RhkoQvuoTgW6Q
2JVowNyE175JXTzdzrFv0XForVLyAHRGEnwHHS9MNy+9dWmkU61iHxydGyhlbrpL
plnKuzhU36o9i+FP8nPzve6jZTUnUeH65TI7nefzRYcyvR1f1CYwNHuzO3/fN6Ic
jxxGXvm5uIuZNlCEIoQyv6rpjvysos/QuWI+xjfHSxliBJp48lPrhC7AfBCFJjKy
9C1f9Ou2LuqNk3PpC1hOAwBh51mVCjh//ABHSU7aWKMfnRHpUcGtHe/DH7oWLwCf
sRgBNcDcX7TWhNFJdXeyFUPIJ5RxbiQ3816tSb8SDQOoheiuJkuqkq9PPR3v8s52
3Xz1EALtqMhin9xNYIluch2vVUaB2vmhOJu3NJn9tXdGGKODnxWVfQmqvQCl7Eyt
+CLkPWE5oQwOsD4UrVN1/xrGEVt6Kx5dvCL/5wm29ctik73oyTxKlYoHadMTooZ7
ZhrlkzyOi6Yy7sFNMWkn9V1tzYtP6gYwORk7nmcZTSXPZa3LUn3F1QYsT/wCpaOa
doe1k4RSEGldZ/IgVHc2xM1eMc5gMJ46U2S5UqOOy7TO3gH3ch7IONIe1XrbXqtQ
nPLeDVN+2eVpMXzk345oevY5AsFvovZ2RrDumy2mIM1LoXA84361ZL0sozmEpNLD
TKeCCn/OBQ+h1Z98s/3oETNxigpFniSgF3iTVtOnBvYiN/ImRuOzPQiMDo+kS6EO
ivO2iqF+baf2tJHeNRYFFJZD5evpScSGi8ZCirURuVEkIKawd5l+U5ndrrvsQXKd
8Vd4DzBg1ykxYGrO+7jtTaInH4DKNgXoiYRn06b9QoxaAqp+Xlmiw0fAe3guhS0t
vbnuM0eirXwWS5eN1Z16Uw9ze1+Ld9L93WekNXdBQ39EMoqmd1SxSa2wkoonvF1V
pc4KXGeZvzLveBTEzmPK7LEIXFQn6XRUsTtI1AoSypoaR4aqznjs/P//n8luyC9p
pvtZ6TSavgflnBTZC9iNs3fLqOKG+bdltuzQ6YucC8Tz+ty9W5sqHe3CdAg07+II
/7K1gILC1o5WM0l2YiiiMyCAO2m4dkqc6mPC9g8FSxhMblFVM5l+lqWQTaVAAzYu
a+jq+ZOagSBIlTh8R+4xHfsH+4Cz+2Tf07IDClUxy4CZmIE8VbD1ekvd5IvXSDkj
ZtAi/PWozOt8rjbopgZPWS9GFxlZ/rxJu+s6ZlBkYI1RQ1c07qH6ELdkKk4I8dlR
p+POvJUrN2QUWl5DYPAMNFZIp8xvLi5q5pBjSw7MNd5Qv+2lzEnrQB7G5iKMmmWE
LvkiiLtuaJ2FymmDLvVjMT9gIOUXpjNv7sr+bPoaqGrGfhkLHlSQFaTN0afpkfHd
RXaJrp0djhBQnxoTzNwSFXCB/vWGlqx+rru9eSV1JKtDF5FvQArS9uu272wxczlI
a1CHl4K0BBYvXV8PtYJgiGDJpuvP382lpoTI00xZvchkvJAXwJbssP4llOa9gSAV
1UuzXdwR5EqbHcFKPWXbNgJjgTw+V9wqlSgEvcjqQqvLYQzq6+AkP7nXqN9w1De8
KhqWwl/WH+G6i5g/z2h64mR+eOJ9BmXgf1Ei5T+1WoIC6ImdheSOvwIRgiIBk/MA
NIcNI9nSsdQgsw211Nt3LD4CwhcLJ/BB/EMIcnwsCRXF3jiGe8enULGMa9H8siWF
LuMVeFArYKeTs7MjIdG9JvkcOgxzjMj/j+xSy6KKuLswdRyYf4SqlljvKUdk2vRJ
Elotrh2KQpQffJNWV4i+0MpeYsdITfyezcHuYtqkqhB6mS/TZa4AEDcE7p9jPFi6
3wJiublEqfG4/6G9KiPAlhkV2X9qd2XUFcy2Ge8/ecueHfVwZEpATX3CeBCNImQW
/s/jx15Ah08s9FspVpjq0qUjf1icScLjVkN0lUmGMRMWqQjlfdlkPg5eynR2/D3b
za4eQCBGPdTFo0iyqpio+ryHvPvoss7Txu47vKJSU+ogqJDkPSMtweeI8pZhrGl6
4BA7C5hNDP8Y8zUoZqPzJvYefQ4lAdHxmPD6WBul8LpvNcgBxJx5cozSY1jVv5rn
KTGP82bNZT8HDpJD/AxE1cZUJ2JJlrXUBl8ZVfgDz4M5sK3V+ZeIP43g4PH7QGnC
rWmboGx753mFovIfDjoKuBQXevm84PaviN8Upv49PRs+IUGA1RMToLqGBnVkvMxd
xY9uvZk55XxnbZaExXaxmotFs75mnUW+I7fiecnBw7/dWvy5RtTCOzQAPSjKHN4R
14GZ8tw67uXtVRbZBJ6gFlmGybLRYapOOF5jZT0LRdy8yggo9UhsvNcVGbHtov25
HpBKewg2JnwnGmhZTrQ+rxpYGTJ9dIxnMsIiTmy9eC0L9uLkR/KcUrG6lc3mvAMi
LM3B05UrM4JeCkk5Y3BxHTgugC4QuTj7Fdqm/+ODHUPcOpboyGmnBVHYk6fUpGou
OnbIYB1Gzo3fcb0pgw25jVvvMoNjsqQKDdYST/cmqCYUPmf1RhS6vqAbknG+Gnrb
y9n419nU+6F0WFXkEJAJYxkDMPYX45kNlKL/BIi985+pHFGCd7VG87Dz1Y0t3ubD
PcSX5HyS0guTQ94DohLcAY61ebtHid4C2GMZdbrJLnigSIedi01Kifr77WENI8Ey
iQTSBVJJzF6FqojmboMRADpbtEL65eA/gu2mJYa0yoQyVW1vF7vCwCAT6JeT7P+a
mvvA61kYpaLCNihZ4SE+qpK7XYkMDApcl8ZSr8gcge/evACLFWHwhZrALIhFXBXS
Wd/uNZnZOCjMYGg7qP8e+A6WZBQPRminKyYhddQWL7U7C5PEs71y/cQswJmLJTc8
DSk/A5KYHo2DaQbp6Cg7tDSqmdWqOoInIMZcsutOFbrzSak0/uJnolxHa5ar6g0H
5tZc4tw7yLYRXI9jlcBOhsPsAiJi9y/nmFzaf4c9CjKB3zJl3MAsYXn2gG4TNljm
RIFGhmiB2gnavcMuepHtI1BoUS6W2dleplYP1KWPXoeG7b0GDHmy1A4dewSLiS4C
Nd8MRRTgJmJdwAOs/hC4cddVwq7ajgRj+sEGfq01Bx0Qj3pDj2R+kIEHI14mGC3L
FefHaIIB62xfwEXEETHHvf1p7o9RoKbGibZ89BcIPouw7fP0m5OTm1pSmDuSXK5o
EzJpil/XSigzy1FCKFhvQFuzpM1rNgFvgC80sBuHMCBmf4vC9wey/wjRG3veiuNb
G4VsiLINaVo8nTnXTEfCdFTw/QdRltbdx4qcF+onszbrQPW0SoJreXENTJs8Pj5y
9mcGoGxE45rLOi8CeFPZLXIfeR2AXKx9G218ttF9caDAf6XCBFWMD0wPhIQv/uPn
5Swr55TLfAvI9feHtflTbzszbAs5wELga6U0m5cO5H5OsUD2cdHeYQtBg1npf1/1
2hvY/C28xO1tvv3lhMEGSaSWEUHS4FJRwA+f0OID5ygCvCgEoIrgxlBW1Gk1+9oZ
19sRnGuusIEim6+QXEzFGyD9Wx4oi9Xo2AboQ6M0ZqOFQKppXH48VF2/cpBAUYX2
48tD7DJsYRcOLCQt40sdDdQoId8B5I5l0Qm5qaT24ILJJghQYXYMSZ0cV76/qHra
X6pl81d1oDeLNL484kenuZ/tPbfgQGQ/Cj0/1rYgUqHsN1XB5w3BXzUUUL5U/6WJ
WmvecgOUtBMD3HRQwyCEEc1KoNdHKr0asPI1Xmq/mzE73fT16M8VBFtvirbyrorz
PXzMkxo1Ya6lRZRTs+6vD2kgSoEazZvSgk7FB/39q+9HudEgoq1qW7PoHv9nhGOU
EWaDEA6zHIz3oFAwau9b2K6OpImJxa/ZW3y3tiK+nvsyJ/Awja62ffvTfIJ5Ka+F
/5NP9l09pj9uBg5RKkjCmIzGX51Dvbvu07wUX4tzkC2PjDWNQl263ez9iV4ixFLB
ARXN+0US5bUt0bqVbnuD7pKy+3bR6I9j1Amtilm4FEfdbBKm/VMOuA+4KsCulPj9
PuMmJigC9B05H3xm5Owu1ZFhfRyd0gSMEBJGA5W/3jLbxYUCkMiDVcagGfUZWGRI
P1VTxAIS/MtQpj6BnyTiGrZlJjB90cVhOnIQh4NLcwJsAjIhacq2yS9H1Ar0QGoN
em4FSIOVlw36wFlNJin1mo4O4GZxrdbqNP1BL3NM+suW6ufZy4DXTTFszGm//ytn
oGz6y1xS+W0fh1YjCh9fd2jZ+Caq+X3xp4l9DcRu+JJ2spFFwZfv/qpqWrlIcjR1
Mj9lGTU1g0x/4OusXaGGs62sTRIwBVO9Dlp1e7Wp2Gd20+2a54ytaXmkW0RHG/np
W8CvfV007QDZdKtEVSkDm9MCo/KCEN4uZI0aVANvMT8+3T251Mv7tmSDj9jFGnQv
NH6j0J8M2pUp0BQY9uD1/TrLjMcrmOrPXLPS4v1Ylm2TfInQVHO5KBBGLGJZP3l4
HJKKV5jRzH+YtxSEyc2nP6np84cjS6Gm4AhTJ7cN2fSJSa7vwADW+05uK4C/gVa7
nTed279GtBtsuLA6Auzg68Xltzqgzt/Zsi0QgX9S2yt398n+A385X1E95FwKgWgm
2zD4PByJs//XTRiwvrxdJ7+QQCd5b/87PR7BLC3gyTxmHht22CuoFtKc5/n0thav
Q1QdSkQPzNcUzNp0kctb2lyizjWenR0zMKRIBFa3xbR73mfr/jJXvZYMyJcrw35M
Vx38piv4oyuJSHcwVxn41mBwjwQkeIINH3Gx7f8rmz1iHmnS07rcdsvCZjtgU4PK
Cjk2XHfK7zpM78LtFVd4mh8ihcfAxWnmENa65tFDPhzLpaH1PkHGnGo2GsogOJ+Y
wSssredBGMJpT7E+H7mtx9r9lWjaJe4C+bgvlwJfozGWRElvL8Iu42BrxpBnJBLr
GUD0AplQwMDhZRKD82aiNHQOURUwlUJZG9exdDQpVO1SVhaJR6k4WFA6khPJyp5H
IDZ/Ji2G300kTUCYzJnVz8AaECOglRD626pTGopFFMkPWtKGGEKdrtVH4wnwkYLf
fQ/L1P9/Z/RSDcUU1WI5oj0r2FEVQI9o9Jnsst0lWjySs948vqspC31zzUPIdUKT
t/AUENXjk/Gv5VVQEPuOmVGMa1swSXB4evyTXyPJLaaapTiKBvwmQM8ACojxTozr
gihb8hp9BgR1so9DpO5g2YHzg/h4ZBQ49YyMn1IyiQLS7nycqI00sSeTQ39diqwZ
f4tAS0ueo3CDx7VMLPGglachQKpIk7S9wYdcaBtY//HmIgB58CiOXJnR2825i5gU
dLGhfW5LkpQo9EGBtrkqWx+PwadZRLpKssuKu5A78oRtim+n9wFSOAQYjXxx11jS
CMJXijZikdWbue5+hnWbq+TEMG6azd7v0x+FOrZx6Ffil4f0VeGdVnbFqLZ/v+Yl
kZsENM2rrj9yC3GnwWhro527qYCDjzycj1X+xMSDW+GGl4AC12kauIxqcdWc7YAb
CAI1qGzyQC2bhMiUFoOY4B9aNDKhbSOwY2W2TedmXMbzEyBQxClpKsljcTTL0B18
aaLcxnsPJMDwaUcRsdp8A8Opi5ZjHaQRUFVX/LiTk1V5LwJLkH0/yoQ2URwfoxGQ
mZhD+ismtLcKfAQSPw+WseYOYf23Rxcm855XwtrbwT47NgNLIciTxXeU5bfLlT+a
Kcim2Bjch6nYdeQ/rtxmxU81IQ+OhO/nsVxW3dBbV3a/CeOYTTtl03uhfG3N0/qg
kJvBoz9q/YtkxQ6+yBUdWSic6a6Te1mgxxt+zEwK7nERBjcd0Osi45+7PUYE3/W/
K1OTI7LYoqTDowg0N6agBVOhu0M5Xf5Vm3E1ipSHqwgLX2cLmBkNh28Eq9hnT6ZY
uqhEv2QSWc7jforfp2igzM4tuQlrwaSySdHbsiJRAV9PNFaj3E5JIwKlNUgmJkPQ
zv7KsfAFmq7swS6LXhO8KHo/O0L/4alJVBzybhoN5ojyXU5nqL1BE/YNcKUgPcgz
s1ZBET+czD8OdtPfF2Bur+Z/88Q2yMK33vtE4gnxE9kVdmldmo8YNPVwi/Qa+fNy
IJkaRvBiCYFdDC2lsebdyAhA0YU/+1bsZWoIn3a1fOXtZb1yni8at1gvfLlXQ5dK
Zcw6UzVKFDwi+fg+Mb2yf+2uCDYuutB1CQ/GVj4Bc7wV3dYflp+aR6uaf0ZlmnHS
eQ+u3k2I89zK6kKYql8YxGt/oAjM2v0DgslPOcM+I9ocAMWbc3UiVEOXgYZnsilX
3hhPnZtPb1T7eG+AhYZKsrou/PNVCwD+AbZNDfMbm+INb+6Cdlyjtb1nPPGec4LL
cKzJbZMp6mqib5gPrX8Phx8y07943ATpn/Vl+8F8f/XghZ68diZ+d97GkRhePR1S
HQnnxh3KES0jxtACDWouDim7w1Rm9iqgrSluxPxPvzN8ySZmz8RZ0layaLSsP+9B
5+4/34vTjWydDxW3UhLGiGkhfkU+f2B5HBiQ/iu8vc/MZS2g16Bmepdlm/W3XHpj
omoTcgIoHXQz6keTkkitt04zuDZ8dj6KLIv7TswFuleKgLcG+JqvhixpSUQTyLtF
uf081bJhOPHq+9C+/FltIq6TlHY3tELg7DCyHO8NhF1u1bGk1WDDAiwl5dkdf3F0
D3WmhT3T+yQZ3pjmHrYXp5mZB2Ay7ea48vhuVwtsXyYcaTjg7BHuceL1gEE4/Tt+
63/diSBgZb1qTPRZBJzDWZCYsGPh8QkX8aH5O0T10sqSXsSah0HQS+V95sGNWfH7
YUOYyAof9+BYX00psM53+5K4abL4lnIhh+iXf0eoCRcsN4x5iZPnFPVegK9lFRld
mjtMwv5naXYruN205xTxtFtpZ5fDP9gWC1L1oHaelU8mDKTSAycGhJmoHMjFNKNx
Q2E8ce3sUIb62fm7ocPKz+RpMMbwhBGrb9CeuZygm5EfGv490tilWfMgNRxlKtMY
h6jg5mCWkEeZ+rK7OGdX5A+kohaDETi2Ce9er6fPb2gO7pl7Om8+p32wBfC5Lfzu
DFFGYGpkaaWoIR/9suzF1/VRekSp8tteqm/VuSONwIprWqOQHcfm3zBraihHiRRb
tDps2DHVK76dGUR44+3LDVSA1ooys9Tg/4dmxOHCQ9fIJyNWYNpuCCyqYVddgDWf
ABcEpLQdesbPltb45YQ5C7gXye3epnk2Cl6KBt/hnz+skkfZPnoJrXsHkaghgUTh
vycXeIxtkQTTqLt4qTZt7WePq3tjAT2wTobl2beIbfxgH/iuJE4WpANh2/CJQiA2
BiImVpm37MD6YEqNSMVOMSb9acPQAjckU03zZY/pLXApFKYSg8iQRkJ607FyaHzd
Dvpj6OWaLYegDsuzOmtYqf+YpBearwSn2W3WRXN6uNAkDpS1opHJW78i0Vm6d1pg
HdxdIrClVvFK+t5etqacIWt2QfEKAdSbjFaNytvjYU0vfOK3QVevTntpQq22ryOn
TmLE0QFCeW8q9RbGZ9pDhVgCMRDIYHC3dWoHRPMTkMgOU++fZf3Ob9g+QcXQ6azb
pzE0OcgzEB8ZVvkuX4S/y9IoZxAYIfZQSIGiql5nztbzw5Wbl6+4681GeeWKXGhu
V+0HXVVfA6nhFdAH7ukNtY4g6QUuFvgCFDgSAfEqbEM0aANGzSuAhe0u2IM/WpKV
izleK/5PkYvjX5eIuDi/4r5jni4LqbdNxk7xJXp8uPAMPs0GK1orD3cf5aShwY92
hawLMyI8amsFKjQKALWsVAphDweD6Lo0cSmtZ87rXxDpkg0YjrYil4OaAk2pgIx2
JCG+oyxAhR9SJ4UZJth7dMXOQ5BCOOSO9dkFDVRYD1X9lgtrQuU6zh42f9UIX0o7
h6KgJVxQcVi71J5quSATlNF0HUuQxHw3QLJMvDi1kHungDhD7HqDntxtYP4i2vM0
bsV+9ULk4cXFzm7XDwHTkerqoEbx4rXQ4c97dCvGi7xnkG2Boy3YqoE8LRbCb9pn
9K83KK1u55T9dwSwUencjon4neCpmEKj5EkPMWvl9An9ZVKcXtklFWEuARCgHRov
cNuvB70d51uePWkL4e5V1ZvLlczuSAs0wn6OykOJDVtNV5xfe97fTckFMXLMpIOg
jYa6UZ4gc3h3MHfg5Z8hzqW28KJ7Ezh/3+sK2sClCzK+KPzq2x4YRsCbMNBRbYdI
G8UarwJrKouleUgPPGCM16r/AyKbWgexGMbKV7AHdd0LFbhnELZZhu9JGdg/8JRT
b8hLLItN7pzCBjgLPjnz6S9yroZejaipdOPbILIL4BPpEJxTZFwEok6YbOKbVObz
deNVad2Xtd06A2sxsF7I8LGc9QK1H2byIZIvfQUQY5lLJgAWEDUjkxu6HtpkQ7xc
oEt67s8jQdf98gBL6TKqiBvxyqeW/u55nye44DT5qSCxixj/36Q1MqixJgoLIGdj
f1InKG6Q/ZZUZVkhNZra4o6I5YSQlTnslX5olEgOrvea2nqaHYCcfICYiYkGSjkB
6nrRU90/McPhLvac76+benJkD6GKKWOE2LQMtAZVo5cy4t52o7VH41s2/7SSOuIx
oo/I8/R+IGU0nMT1M20fR1br7Kx3uZlkj72jswY8fA5tHEk5JujySEWgHwkBvRIq
/az/u6EHPtavpGxo73uOq/+0Zp9KqgrXguFWcHs/STW7w9ZH/KzGUZpW2cTjXHPe
+dfnvHBAb3mTlVLUEG+5x5u/sHBnirMyys/Uve4lbH0WjzJOdqCzwjWcAu6lQBcA
uJEb1DHa78M/Xbgx77NUaHGmT06DPWCsZKd+byLFhwXzYNi4wmSfXiStKjnHDX4b
gT+etd+DYeEiX/QYS/Rxau8eufOoE/o588/e+kfoQyeARisof/CkN7gItXGRCJWr
4hhZd5x8zJas14Witzx6k0mL7ZFtAIDkDTOwG+NVzjhKrLipeB5jCkePbKkpsoUn
9ahbNjG5Jm8d7pAOBWaaU06nDnpVh4+uiDxVxNJIwRM/Lgn2x0QGZ0szmCa4TYD9
6fVxtVeQFWR82ST5uGVMxPa2eibyDy5DavWBQiAnNEYFnD0eMTmV3G/ety+KNL7s
VkS+hukn6+Fk+cvNrf95/hVHBvZNAxMsIxVbhTMdrhWoErNdH0OXHDdWLhOUgT39
H8xPxgNeFVjg5IIRgHH3G2LTTgaSYE0xAYqmB3o2RTg/w/GsESj5ao78Na9gkvgt
rBn1E7x1tPnXJRohAblbbjrg4xCul6p+O8U/S6uyHABNamMDnTFNFIJkSsMztShe
d07OInuZZ/PNR2IqTmuMfGrPgvtwcjgkaeZUpDNNEYc3PWhfM2BD3ozfnFccwkPJ
Rcs3Y2yDj4oGZOtc7rNC1evGVGvMXNhMfu92y9QX8mkG6hol7tn4PLBSQuwkz1Ho
1Q000OQB/Y972fpTAYhU4XNpqN2gPkLlCVx0HYgYJV4jvebzHeIwpoz811I3oKCG
pZ2236B3MfJ61O5L5lbaxwSeP3ZuEsz/tWVZZJaRiMr88YJnYOa9GWYfNONG88Wr
oASz+E06msVIO8c5lA2xnCanlIanSgVSwcpQHt2YzDrkefuvwe1vCuUxS7SRWBYe
ZYxmzXOvHkNHW79GYCcIJ8DSqO6Z9zIx95xJsmOLbwq38JeS53laXXIsfGIjWD60
yuyDSHpAZwRD/vR4nJ/ABtth/rgHDIDXA6mTaQ04tNvOi/xFSzxgasIJa7MR5i+0
/6f/kaw3krRqSB8bl7YnC5wYGgbF/420/hlfGGaJVsJwitYO8dqzSqqLhb+l4CXH
snYcTcN4OlQupq8lRffxpgFzjLIbWSOd0rckJSMQPcE0FmFaYMslqCythp7QXBFS
KxLWDjUPn1CgM7GJf+r1IRyoIMABsspWSksKspwMDw1R5IDcEXutsMYJk0NvgSJp
hlm9w0FwKSvudmr/u7Br7DedcW2XT/U7Rs/Clx6oScSVl+qdz8zvgZlEj9gYCmB+
ocSPp+5q817Z/hbtRie7fhLpXOxfuEu2KjbsJyi6maA8CGIwZNRkS3Oxvpg5Yi/O
bTkBmcVvo2Lb5RB1FQIr1DGkRI1kbRGbU+NHQ3F0lSbiTiB4JUIybkkVdp67DFTM
M2p+3Z8l5CefMb1vsAUgUh8HQoSH38dIiWDG46phSCfZJbFMPASkS0xBlHN4IB87
ygmGGaNnpNbzbUfPpYe4tdNp3JNY5jMLOltHsqZqs4iomZ3xP7S+PXyggBypzoyl
mnZnYlkwcA11DO63h8KZdG6KI8MAKzYCjztW63tpO16fPlFuMzlrdDOduMT6aEh5
YOiF/nyCv+zEgcC+Wkz7+Cm+B1gr5E2ry4wc+13baOjiV5zt2G1jN+44qVu/laEQ
GEXazfNq2ib3uw9W99W5hYq7Wt/90UXoKihtWJylnKIM0vArm3Kv2Zo12a4pWDG8
x+JsZmFIUAiXKvRi3crKYEu8a6ouvfjoYyywtKWfaP/iTUAmRrl0nw6ezJwzw8/g
mN/PZRE4TwbnyaRUHV/iO+yXw9bYv3wJyQC0YX4N+EFhevOKYJ/qEUiZ4tNR+WtJ
6io2EdDEgGxipq85XIhLysxCmRLQsbCYIMt/Mxf9fi+wSoNZ2G4pCoIacJmLwABO
sT4WFdHjQ/w2Td2zhS9trES9u6g7PTDOgRwhddI5pUC1nTRAeJNhUSWW26qKatJo
UG7KN7dyLwFAwgJSl6wUXLfSYaXjt8d4NiHh1EFtYBtJiBajZDjuzt+g7/irXLVP
0WJ3p17D55vQSWY9NMV/Lcqj8Bf3So7lYcXsBev12T5qafCKZGSNJrE/tprI7x3o
+CtHmWRIf2xbwwWHVkURGDRmildq9kkDTJY3Ah3Kmi24SbNb0cZpLdSDxgbFarrH
ntE/VjAL7Fl/NSl40IDcJWXJ72Wypap2Zs5xzmR0aLcTlhlkiXLjj/bBN4kMj+G0
YW1n1whBnFyfydi4bhw7nsT2TgGJM5Wqm8ZlzziH7fLb8VZjB9GgwQTH28pC/l83
uLq0Ey984CLlaJ4PlWeVd+ljASz162aLMNcCk7cZDzP/TyJieWnmhaTWAgNX8ecE
nfYPwfx9AG4EeGkpyAKSCqcBnbkIEI5YvgkxVK2DFcDusr99YP1XCISq6q/v2PC+
1MvXbmK5J74/ytsMi9KgXZIGf7+0JPGDVPBl2Tmpz9pTaNo/18WJ9lAY42Ro34vx
yaUxETOjfdlN740HoRHP5UakALq59d8zSToBO4bFK78vToazathv1sGjDyQDl6dN
lJb7TU7TmdzM3KTvf5KlP3jm4phijLbaw6+wqEKp2js4S+ux9oua6jjqVBoqhzlD
iRWcfDXafknP/F4xzk2lmx9qrVQnFc5SKlBK5z0WssbBmHIauaNiDqlRsahPImXx
4B0pb0Pxo4JHIbbRLIDBTAB+9lWDKu6RVKb1lyIH9M7U+W/L7A8GZgerl0klJgXm
TV/991LB22yaKuxGSjJNCG+UTZY4ooZf83FOkf80eRA6XzRmsIF3w+mzDZn1Cxt5
m1pytTEBbcmUNibE/QAIw0V8vW1RftwoRxhb+Wn6lUEjXNPXQYsGsjYJHSUsWgQq
uvz3VQ5RRKnE/YwJVY1yLYw4utCG08uvsZ4mkwPb2sRbgjvM1dF69iWTIlWsj5m5
WzlRjPq/Y2C8MOVOo3b1OK2EysNMEIUacWTFI5ZdKcW5ySA4ZQuu6wzbjV+Ybs0Z
JJbix7UEzgmrb9pS7b0oYguDOqPZfSAGNWhtSKoFsQgMKdZfGcDL5Ch6Fw0K84Oo
8Cjzjchtxq4stdcxCxxJhSuYJ9FpLrWzS4PLbGyCIo6Vifkipz/EAFW6+YfF+iFw
j4eNKitjt9U6/hwnxT25F4Awk4KV5tPrGF0/La+IOujWW+OlR7u9rZowpG+HHu6W
cW9J7ADBXS5s+vfMFeCHNxlXOyHQtcRbKkVtu/1IjV8W0PovzB7GZtcPEYIWYCXv
B1/3kuChfksE7U7SMqdbQWUc7UNXHEtipfmPBwciLP5KribeS0oSb1ywaISINHfH
nB/6pttzbeJL+hPORuiPh6tWm2N8RmdFUWG5tk2M+bNGcfs0TyBsdFtEVZ5sYjvx
4/ielOPMGZC0naX4otrAqq+t/PkSqWdXXBr+ntMHYWYz4npLYyS3fa8hDAOa6sCj
Zdg1dLTnOwlQvUWF9jcGVWg4jq/j+B516FIKuILF5BC5PXBn/DBRzQsrpNIorJYV
uJBkxLzEjJgxKzrB07CXmroJGJ+IUXORCZ5WUJ8XPOyunXQuG5vSCf8pspZljWBC
RW1Ii8ydxWe/rX6ixnSqAktir6sECmJSBA4S/2V+bbyJXqgCELpDPEFooglrfxpm
h4DbORh+89rcq8Fli49D7zoNbs+xZeSyQXfTO9lUy43gy8dLO2558u0ot4t1y9Ms
SDXL4Imm7ejLLCFfvF/EOJvWmQ3Sd+Y6vnr+CZAokxV3IdjPg3Ch53CpilgG9/ct
DWxAOFwYOHTgbp812+LDGwHAsOhw+2DF04fedzcWZyoM+283InakPMcpv1rC2hxH
xBfiUhSIFJdCOPXNjGQmY1urPhOwt63cdt6OSN+JXFZ0IyobM8tYKeI2PNlY0v9i
8v0dvnPItoPXnc/9cTMRwxbh9qdTzBJS+/roFptknQNpSlVSricI0ojBwl/yDFe4
flUwHmJO8M/NvXmtdtbQPKz9wdzeNao76sf2ngzJBmq8Fh4a7a+eN0KtdNK7cpjO
CpA+ygBLVgaCKNwBu8RXjcbWQ+8D1MKPl/u+n5YQkn/i8vwRsj6tPptHPRg539ID
g01hFhy4aeKDaKLC/XYVkHa+gMEZPlgjyuFDfhn47HCA52DmjQfxG+tLeYUvaPk4
ix4fn8naBIhjVOIrBgofQxEZFXYJj+jaymsWnVA47WNjiWDWMVAFuGZewYG3AAKO
0KRWybmWyewVrLhetBg1YJwErJ305sdvxyood23MmE9KL8I1cCQWLZTfJ/etQb0n
DXO9AU9EfgK0Fzj64c7s77Do21sejTeh01wphKjCNvU8pd8d1+5VPggnBul1jCKz
0kPblq9dRcwLAUYHbTI+/4wacRhdsEVma6yJr7+hV8ro/aNwFsNlIrJ0jrxGkVtg
hNCPemVt3in51rU7LmBvzLtGwz3ejz8ZxgS53zFf1915acxlkUA5pFkzx8sq4Wf2
su51DkM8JA5rfLW0DkQiQhe7595jGjO7m2Sys6lsBmAEdLrbTRdLG8UOSZJ2zcom
EMK+NpnUtxdTP+HzY49kSgJLE2BIGoKPiSdgfyA4Dt5H4O8SjcKorBLd8SvewqB1
wAZnyukF/AyTpZQwS6APnMjy69J54/X03pPko7X/UrVbY82v82on3jzxy780IHec
ajQb4E+/hwN9bvxvqsqkvElSKKGz1RfVjTA+k1n1Ls3ijHZ1i8d8l7zQysaUWFtm
OXDSDdR+8HHtlcpTmyzMyTLMA9iHKKE4ACVcjp9amrbWmdCYzSs5LJOQxKas0NQT
6XGGnBwePTNwlAUhWyq+NNUD1C0FDtMxJGYKCrdclV2VdWjc0AzugB9tYVmQ3mWg
VYddurjP3NB8Ws65UWi258i01e2xZaoRGU8HZnwRfjOQv+arm2lN2G7Ki+aor1fP
GZgsncv8BoSkLUd/sbd/MX0pwyKJPMUuxcJW1lrwjpVdnhgShhpRRIyE74DQ68Cs
Ml3hN8qEJW+yoSjROpxzF2BoHxHoY9ga/ISzMfrEtRYzx7xefBeTAlVxGDeF/bWh
flWod833H0R2z64lsozhtFFjarBduUzBRvNeB/06DxLeg25H1MxIFIHnobIPG2h6
T8Rmkmsws1GSgONQLruv78GvjdGKRscu7FYtV+Mmb+kcsop/1cc5wtzSuiNIXtGo
q6ql1T9FGFNiPfRE3bYpkGAGmfYIgwIidRyG85fT6m4Gidx2Nd+EJ2vPnxTLOxvu
AACfRRzWuU4O7//eM817tXuM0H7sG2W63GDqjK6jiy4veNfQWdBL3OpbgGIQ0EzH
YM0f8cvOL0z9MN6wcpeJ5RWCnqSi7NDRLyPDs4C0X8S8a10BOiokM73WyZIIBpCu
LcnpmoK+ByDVSjnrp1Mpm8Y+QTfLwKzTX61QY9zw/9MqQt0ERW8AG+UHrN7342sa
BYfCZVOhyNoNpH3H5rAcCfsdbunxDkDg0rK9vVjA5J0jojTmEkkJ1ShL+pXNYEtz
Tjm4jRzHponuw6fpsq4mirWAuyv53gxGG7+XGr/6KOKAkqY4rc8iSJfkbLyv1Ve2
k78z2339oFC7gw92WHkY/b43riPrQ4CdeniAii7sxiz6I8zFNJS29g0EkMbyMOWs
6t0i9b6KN4T9Qn2d7GKprUU9i+/IUUzKrBcDSA1lk6d10oWrnYMvR5ItcmhCdfMw
8wHesq5gUYq5tcwHfuqQHv24zxCopF2nWaF3spKTDPjd9IsNISCiHYnW6H8DbGTe
8riDwqLy7TM64P72DoID7olP4cP9lxdt6Ppl/9/TLi+hXO6V+/FOHYTYZNFliwFi
4Ht24IpKX9s2W2JCLVfZT4I+ev8ZYoVZ3Ztr27nIFS2kz38zYc1pOJfzD27+VDdZ
RGECN9kyEdX5fIHSwEEp6fc8YoEYo0g8CTpLWgkYCPntuDXjgULUACkc8zyBVxJt
pw0tJ4oedxsVImbPQsQzpc4J/6xYFf4XrC500cDu2eppTQ+xinlr6xWTjuMY4IYI
xNeTMugXUXrscoI9/i0ofWpVdOD/vEQ4+iVO7pslsK5hIYIqChSKN4xDUWlEk5oq
/ErY/8H2fLF6W1Dj9r0UtmFYT2CfPXkuH9GLaGNQiHwGkCLswmiTL4JlmYELYC4O
2X0OYqs1Tc0M+PmmBRYb7LL+BaP97mu3l4yjm4GMbT37ZWWCl5OqeaYhjfpgmUCs
AZAj7cqBY4mrU4BLoBI8gne3GojWOMT3KQr5giF+UuArHbxY+EQieBmSUiZJ5DK2
0DmGOLTJtxvmc5mP+SC/MPG9RFfluNhu756SjKm6T2rktxgp4MN1TOlx2EFPT979
lEZmjCpZK5UzYPbnSkYCFn07la39tVjvOedO9sQHjsXFETJU1wp18ggPqCVWD42b
OictNf19YZ8vg8RpSOHqkjMAe9n8L0NY4SiXcAbzgAmPYeO9aLdAAHh/E4B5q6i1
Q2JIEDRm/GJgOGo83Bl5t61xUbYve4k5UDGpuo7D2fy6f0c6rcMmHrilJdWdCaL+
9cuhPfU/Iyu/MAar/0xCY7LRl+j1rUXPz7a/PFHVmZXpYUAAjDA6lkfZjVwVqRTU
3CyN6TYsIPYnzbBfSaV9uOhBOzh72pOSh6lSYxc6SrCAROrBn44a7z7GQ1GfiwtL
S3hew74hfEc77mIFV2wC8qK16/rsk4vfYJjzbm79QtUFyoeKm7d15HQoglmfrv3p
KRYjForf27HXtkII+hKP8wWRa1A4VwRlAoOyujkuEnjPeWtqhJ4ZnJzNRdIotXAi
TM2c6JG1qUkvSLdXmj+g3pyEhlhaJpS3mF+doLkVMSPRV9qBIlvxkQwXKD1EQmiB
NH8Pac6l+biMrGhgw5Nw1EWYHT2+VZ6lOq18Qk0PHqoZpimw19LAln6kRP6/3vmR
8mydQvFcKI21bhvgFqG1DgPaRGh8Ne3Is3t9c0aFQ/KyoucErGaH9rmS8hgH17Dd
PTbwvQRg9cILdYxzxDTQW+IUTYYEMWqHMXyuahxjWbZPDawqwiUkYAct8wx0Xa9A
UVktmkoIRx6g7s013cFgvLMP9OkuPHcJIbjiaontIoM2QX+JbOFAZi56jPt5vD3B
zhDEXh9U+eAmgcZPWgEEL6eeADOiaZW1awgd2paCa64qN9V3/26y5X4JvXgj4i2P
OIpACkFbO7QNZYcl6UK4q7MV/mjm+H1dKU8RmKsmi5T9KXpx0TVwGBVHtQ00+vD7
os6L9cieSESXOcHvLQ7ZKMT8XCfoh0C7zlds4yObEqFK+NpacTGeMeKIgs5U2iVt
XYdKz5LUmOaTFDMkhFxAG0d1HG4dGKTaq0KHKe1QRkn6qhdQFliwaGHGYqrZXk4d
/n/ds7U+q8QDZkPmbA9FvpWZdzOOLPJtj0uMgvnSlFgdgMzIHyBNCqmTqZ9QPHJC
xBBTh5dd05ERH17pswLOHedt8ft32paTsFBYSAuRVt5NBuSL70LV+g6svl7B7whU
osP0ENLR6TANU/5S/4Ty9s9BOS0FhWDxXg/B5EsDcQd7rS4sdgLGcQJ71xaaeGGZ
CZeyjFp1/fP7xJkjE+sSPPWTyXfFfizfJ6lsZ4BwV4QVuot24PxD1op3BJdx1vEG
bU6tp/k8xm32BZIMPU7zK/+7uh26Ik3JSllobMWLpIOKyawkDNXnAPIFbGlXeCJ0
P3r9P3ef2bJrEXLDT899+1wRqj84Z/Ly84QD4u1amoRoaS7LvC480Q5u1jaxi0DT
CWxJK5jwYLfVAFVhJTmFZ62nrbjo/dEWQprBSpmuiXwC1+9wEfwJ6CAJvavItOGm
BZw62XUZpp0gY+50XHTMgysJXM/0FRAvSXtXQ4kwYpXmv4/8onWKTj9FmPMeddaD
CRl1zvCqSAdh9Clhs/Fyh3B8W42PMTOolDgw/F7eW6UhQBJ0ER2HnNTyNMHNpxxi
7Ib7jZOdKLcB5LYS5Eva9EUg50XEieBj70hfePn4U01T5CvA5z2f2cW1osxy2yJR
lcl1aNyoEiJ8nEhfLX/ywWxdop0DKfL/fwlTjTaPLpvR/O6qbnX+jZHL7msOvbtf
mhHs0jDqEQvfSgcDcE6ZkaxLCwPrU9t5RvHqReg0zPCTpkZLWHnZK4VY6h8AKu/l
f2P8T3QHJI5okdPMxgRuIompdOW9p3hnn+JzxMeVge3+lVAFJYq4X8iKVuCisF84
dv1Zrux95QWvHpdmJugoxhdRxj3bDs8fZP1XazZIoxlGSyUJYjobqZv+B5VWy4xx
SkX8aggKrn5Q2nv+FSNQXP0NeMEEpIq88S8POfjx9Z4Aw6hDMbD8jmU1gTun/cwQ
jVzY01dzduy4/QPmlym4AuQxqg+y+2vOko/DdSoFMbIuNFnhk6CSRD9+7+SX+ZKN
DrmaZuSbqEtZmp2MpsILw6XCJkBch0DSv0lXwxEVFRM9xqJByBoq7ub2ly1RytLd
7xeqM0D3aB/rLlR0z+BSlxQqHeofJ83UFC6o8/8x9jDevjZjLBgZ2F9DDmesDmE9
J+MYq7tTk9v3G1furDqVvGVq5HAgZrRm1JGwW7hNBFcKOfphQfx8MMOJyO4+5bOz
jHWopUDPOaj/RS39Uqfvd4yjeRVjk/gnM7K3hMkREnW1ypm2d8WLJa3D7z+89bj0
uBOc5JW0JFkxGSu8ehRzhQwLahs8Xkv/7XCTDacfF0o3dP4/JJrmEn0U2kWFMb8I
88psYNeo50yUZ5vpu1y4sFzrb+efcMno/aTDV67MECQeQBLBfB+O5WcwQ2dajz5c
vgiZ8uYu8bs3NBDOHi/7tmqAqpf+BZCCauLeJ+we8sGFfjJBPId59/fqTOsAmw2j
vGcGl+D+hYi8W/rN2LajiQ6uDLxgxTxFKbKdDwYqHy6y0a9UXF2ytnr2dDbFTDqW
DHPWT2+Sh0qZhj61joeED5z3zJRGUWFgR5bNYUpr1zVZU96sRx6EHj6XfA/iyOmS
t8VAPQMD787oNiYLEzhofWs9WbKTnkIJ5MYgmZxw3iKqC8GXTvVDH0g8XoZOE3rk
xbuKWyRmXtP7azgHWnBZq4RvTH2jG8rF7f93P/zJFzEHZhapshvj7qp8CBc5Zy/j
8twgYZy/yqwJuJTsrDpLeEHXcYSBtw9JCCbPDqRziymHxuWsiv2/tuGv3ZjLCXI4
GSsjgiI49yLdNUdzev5F/zthYgxGrK0RKz4lzv5itJI432/Jzqq4VyHi1yl6eTrf
IiSTNrD/Ruxzohph81wUguMyLO1MxAuTWlWNFo3dnDqIApBE1Vd60tg8OxIjdsW5
4RCbDOzyweF8zlU+29xc6IpjygTeRsy27Vjo+KC+k1UrqqvHENVBPVT0CSqgDwwR
kh3DbLRpamqwboKQEfdHrBpepV/ZMkznMYwE2GfBZiaXaGJkpIfWWYDRs9niiaDr
Zp1QLdEfWNzGmODHfJ+S8AwMEbTn23C50SvwsHkaCpvum5iNvDNMBRvfr26fOj/G
GrjPsxq+QpwGUSeuNEJjMvgsz03hwAOyrbzWxDCm47947H2rsCLawWL9fsYCYhtf
IxxjNNomKbyZMrvAfpnY7ho6axi84NInlgYeiEsTnPd2hE0RK8i+DS2vVQgFc/gi
o0fSCuO0HgOD80fC2EfCxC9kZc4z76y51i0adAP3rqdr8cNULzj54CU4ZxJ28AbR
U7/n9b/SCQ70yuqlnG1jgbdtjgGkRNlIh8N+xSqitvHxMT7cjlw3ct/8Mg+UpftW
MWIwme/4yFOhzgJ+/VKEezhPDEL2UwHk/9aI2XxjCwVkjlEbw3CSG/4Lta/B+zcP
xSJrDlUr2fcwC+AMeZK8MBVo+C7+OCegvQa99fQU+ZyRVZoxc2VgZXtYcbIw7iuB
vRV64zMKMaNSn+pQeKnNXApTObrviDbEtTJgjcmpEM4eGeqriRzgTUzK2HGZSD0Z
TkEmNhDPVahejCmmJbdkd2wjt07Y0zTFxVCnleIwvMl5r5ZHNHWNzZyR62I82zya
KtbLZQ7d+Jn0is9SLPXi0HThEY4OAKZ1zCX7I4fCN1pSRDx3/PysnOfvYptgVymZ
OQh2/iGy0sWCpkIeb7QVJDwT19wkAPsWoYrlxSFPRknJqdbEEyPgjcOUV2MZyoPA
jGcotPYcgkFZauzGIhDpo7X2tyEQlpl5Moiyb2iOaTwQiwkt0//OfHWPIdanyV7a
QYcM266asaQpKDqA4QOfntjH/ZXtR6fUozrkmx2oMuxydLKXakN+UFN7UpQpgKvl
jTYMZfXKLsXfSAF2MhZaJULtIZkTij9hJnNi07/ayXSRJlUem+jq6sE87ZDjCFFo
4g4RZ4KFL25eNCGqTOLVuidiWDHxBYR1yIxzCS6H5cQ4o4BG4vnArfHwLHyyoSuS
tX34rdcTI/HLCJN8WHA8JViEfyVs1hli5shZh06E3M2+WUE0yXLC83oJTZpORQT2
UOee+JdRCZOKuUa3rOGx6Z0tQHfwnBMep4BBRO+KyljzNCqZdLWHmaE/q+cpTnlB
0xhQb4KhXEJC/cu/xfvYTlCm2WSDCWJGyuj+EuhIOEGAnwJtfA9aV21mczwIGG/n
7ly6ovplJCU8tzAHT/ygQGeAdYGQjhGq3s9TAIonkvPW9aSTmYNCvdJOlYwuTxwo
AVXS8KBqd8DfHzCYhyoQvyhbYDPXjOx+Jw/hO7bEy+rZUOC0thwh3vOH6IZWA9RD
MIo+jxNVmDwfYIpNeyY+GWwpHhz8kNu6X5gZR+9Ma8niN0oABUh9q0FT34894gYf
5uVq8rNBy5b3jSlA9NM+xDdrAT/KiPIlDI/xCo5+fjls/HycXbKlk7xYJbxCbUy+
kUOCzAxlm1TrCGYfJzfKOxNt8rTp8DiGFbJY77KtV2aeJkYp0ni2nU9uLryZXhxE
/xAlehioG5neEL8G7oTyHdEIrtu4NmrhiP0nMtvdO0D7SSx+H68rRj8qOItp/iAQ
ymP6hkyaM4mHQlpF3TLdcUhjqcao6O+XBbW6v+25MkhfBSWRnSTAJUoX+ivMIxxX
s0OcPKJXQuH3+8eglrWWLcLdrClprGLP/5ejUkNPVhZTxBLwHlRoGtu9dkG+eGne
TmvEyllKt4MMGRFrydV2Zk10Wp+B2HoaoHRmtLpGxZ1y0hkky5+LSxYX86DrDKbJ
VJnuim/qRKMOPO5eTTH0JKJi+cwUoBvDEIZPdb7YbZGZpHK6e1MF7Y2e9t8Dh8v4
WWbs/VSo+Lzs9B0i2DIjGYB/GAco7Fsb+0DUPibuyygJg9F2HeUzs+vGPj+q9PNS
SAc8H+17G7swVGRwrFxW7FRgzvkKashqs4RnXEurfdNNwKYveyCe5TEKyRSMNgAn
KPH4JJVOUwFktLBESHVmMTk1BdBxyolbfkndn9z9MD505jZNV3WSVZ5Da1p2+z0N
sX24rigPPR6FV1HUri6TO1nZiX2TWg5hwN7+AMkN2uwaa7k4Gk62d2Eh1XZFpiUf
7Vw+URfSNUjwFmut7ioZCkdKUkNTLwv0bNghBAAQONMaolEMDakGGGiFIqkj0SFz
qGkEBZ1OwOgwkaGoJa0kHWzuJB0TYt2PSYDQZDcbv0jyYORlIWsNR0ConfzmSTeP
ubHYEtcxNy39FSAiwifb57ZWw1TBrvLhwYF0rzY8cBjIGzjIdgKcgcn3IfYdgEy2
Uzc4gXx7jAUh1lTFGJWUSsCyv8fUJ6Njx6jomlL8qJcQmAbTYSbkDeBdy3jW2vFd
Yi0Lhnnk8g640i2JYg9jQjnB07OYy/U83AdkA/nXfeYHwiYWvSRykUWsxu+0BHPd
0B9yHAXMbZH67sZCjGXGdtjNLpTyU/v5zwgnkIMLUgFI/aM2Ew8zmbgYV9iKltpl
LbDh/JXtPpMqaVECl3dmutfeuLcN6RsbolrDVRuL91eFWO3qSUdA6Fs/lEOS6k/A
NzXmUiNiuBJAeo9BNhN+InH0q8fONHPl4NlrjFexy+auT0PJq3gYIbLBAlFFdmHs
UMGdLmQQohIJhZQmG7gQ842rmyuBvhWgQEigtBsAef3oObHk5hTEYVvJ2yITz/hv
gzx92lpJ3IATdPQqWMNBXdT0Q/U/qEOgaYVz0aimaSHaPH78yExLbXebNmztVswp
8QNnnYJD6kbfAgSFYnNPO8e+0VABlul9ovRvU4wWUb58pRM9KlnF0BIcCygeW1A9
Q+P3ILgbDOWG1et6QNBUESYb4dU3OXKOo0W6aLz6KtQn/UwztftivR/BKN6behr2
RRsLCV3544LFGyiYPc6UVhQhlSAxvsDlf1pEERViqkxFMKXb9txhv0IYCw5/SP3t
bX48F+LD+b/UFiGHEmOw4uIEMYkQNrYLqHKx5iZ6EuMWZGE+qI5cZru+lfNsWAFD
i4zxwTbU0aRxiLbxZ4pyln0pgODbpVbqgpTGvN4XQxUeBMwaLjYjps8OOcjNLaqz
QSQ6CCWIuXI0QFc2cd5NtAzhXFMSEaKAJBrRzGk8Y0/Q2zM3D5sCPk8upKxhkMfM
cew2uFMfJsbQnLwHfcwjuEsR2qZmUtJpDV0AA1zI5CO6LR3lzZGuyoVvRGErLTyI
yC9UMSg/SlGkDUbArgzRiMCSZI3DuImbMdS+apazA1IpaCb7ZOwgNFJpblr5MI62
nbXf8GNmPQtYkaljndsE153JGrrU5SslBr627c9aeswGljZMhysVqx0A5NTNBZJK
r/pYQCqxFwSx5SqsMednVT7ZiTd53G3wHMIdv7wLCZw8mxP8EIvZPO8AY7INr8sw
Wd+0Tos+CPjTqaya9E2OlMcAADtJsvINjB+V6HFIBKhF/P9+OUOGszmrxpiBx7EE
p7BfNRv9QqEkjUJm+OFVlVETRiT3VD3mEZRatlibo1cMJmDmjP6vjH4G5mytHE9p
95ru2aR8VhkRXrUiDrC47zs8x1ook7CXUpxkO6YOLS5rVcECxvBY/rkuIxLW3W0B
Hlzzh950Ast4+ZoqW5Dgcdsp+I+SoV4q+hRxY74cAcZx2WuhTCLuPO1NF6SI3hMW
svUNbu+LH+L5/bgd5UzqwaFeoKs28Rbiq370912VjhlEXzM0eLa1Yn3wT5Z/qX9N
2SSy4Ah//dnPAVLM+U3GV5G/oMlwnhAfXdJz/e5vD5REgUFxeJ1b/w3DePD1RYSG
jMIoTWKQc/2cKBJ4wZX398yxu9n8LNcLz1DztrX0YKCN8we2oURDaJahiQvYDbaU
2Ecs5u5Dzn4Pu9+yoiTcHtpgef8AvrSaswzStrJKDVaZjROiXQHKIJ+sQGcqyk1N
+xCgJwBfh/Fc9w/Q3reNUNltxkrnw8YPKdBmxAnXGWAJ7fwy4L1Wu8q5aHWL5HXQ
1Sy58TAdslfmDate2DbTiSH6hXQ+yLx7WG11z8yb9oLOHA8ilJ1Iw/Rp7GnlKeH3
4u6qUa0e4Yr8XUfMhtM/EjoYM3hb4ngeTWgoj9wCXHiXrAGBcnUr+M/TptPKU0KG
Hnl/Y+ynm7IDG8iHvlz8AY4tUF81x5u2pO4sSQ5zCfb3+f8rk98UX48Xi6k5mD1y
IghNWBE7bAy/+jM6RGKUznD3UQcnTnbt4sAdTJMyXr28rG04dzwGzA/mZcLH05jx
USkE48roFvIN4T+wiDgpg1czt8I3ID8nlU2gqqzgWf0PM4xLn6OW8LKNezXZoj3x
Y+laDmVNXSTXwZAehiOBsqUjCA9i9kK7hlzo1RnGdDBsS0Y5gQB7TGbzInJthRp3
V//2gh2D/RxA2QdRiNFowZCKmTdlzN/tumj71UU0RDL4gw4WC1guJmdIDIDPq91W
KqJiqzWuBK2+OMk7PBYLSEI+6EoUrCDqgtNK9pBgiW3F3V77DLBvmqePRkh5OlRf
EZwOAIU3MGdZkKhNl/fJtRre5WMHj3ItUKzcK3byFMunCMWT8PNb7+i8/MnLTkJd
bWPnzLZz0X31fFxbov/lA1rddfPD48hvRhAO/EnKwdwmXINACgBAXHjxj1/4HjV/
h1QC+oDTHwasbPlqy0Orwl+INLlg6eDDYYng9w6xxpg3Xwj7vwa29KSz0+dpSwCQ
oC+4gNBG5Qqladanwp+Aahc26ri6+fkWFdSm4Q/RUXaap4x+Q1KlhyZ2Qe3fOdwB
17UT3ljI+wwpFFgRgQczOAYnZny1J/z6lbbpNOz2HtWdrGVCEd0aAjC+vqg0542T
NrHDXhJvLs+ZmZydCWWyd2lVsXOfhftA4vxib+BBZPRs9vPPGwxufkG16GKKRa53
udlQnC0GPxFL0jg/U2lsVDWof8jPLjJtXtiJ8KxzL0gIUIXagBJLEg89EtSxCHEh
kcUqc7oBOns7m7spLW59QaGly6e3t6HK9UYhbpJRqC/fmmyhbdZAnixRnLNwd/vI
/bEjGyRznOE6fNW5SmdeLXWMAG2O2f3mSO/cSt7sNbCF6gBFBnaxwujc4MOu2Fiu
eONp+zYB3AyBaedma4cmb6A9ra0lC/UiGsZ3i7HJyFXeMLFYDnyiRstgSy7g/eOo
m/HVYuTNYpEojszDqovaEAPCTFobLDkQM2Qfvng+pIcuI3p5YhNaIgPnDhfwrejL
FPYkSVxT78x2tc/yOK/EYCbpMkv2BE1EiYFSbC3u+hJ1sXXHBEmPLI92NE/Rd72w
A5aQQqq3qbGA1xU/i3ZjutHlcGXoPLYJa+MWuWoweY6pCe/GuAetmfsSoeUp5cuI
0ER/OO9o15VkTIqsGXHoTHVv1uL9C4a5YjtFvajQt/Bghm44eLQR0NHEc6bU6Urp
Zk7k2/FPDW8ziMl0Te8kGJygTDcq9AaicFePm5TJB6kWKT1qypvPJt7sdW2Y7r+3
D9iHIRKyBzfhnGzv3hH78xr6vxZJJxg1S+AtR8ytVZPyoO90Lhc6YFlL2LTF7vDq
yr55dQFQ+bzCC55RZzvs1SDVtDI0mgiTcBjCR8nP/SIexmq4FCbbcw4vj3cqhAHv
NDfEmxj/G3uCh5L/dMLTxXcvtNxew463/E9T/+19vd97bZfnOmyUxbRc84yDcWxY
YqkirblIR4mpjNUyv20S8rb9KxbeD2GBgL1Ew9WCQEN4dSAdelOEcdaceB2Xxfg7
BC1fJohqqP4g0aR4SkNNJnc8yLvj5KbQK4RsZ3oXl1K5W/KsxynEvcMXY4I1BZEK
ZKUoCZ5MxCedr5eJSY2uyfp8wS6+WkEmKLxozVj9CGH7jneanmxi8NGvrgnPqIUu
ZR8t9Ip4uevLFeD09RaD+5tCLnBpGFJDqcCkMrKOEqqSM+YRROnyIH/XB8rCjKBK
Rbt/CVoOoyaKMTEmvs82OJPbW2AQxKOVPGfO3B/KxWh4WEMDKm+9jwgO74I43sf+
WHXCRC3eDIr4J9XxR+L5qY5ymlY0I+YwUT7MhOwB38T7dVriODjXhZOqHAr7lip9
5gPugmbTuoR4+tFcgT+m0b4cDQeMSSeOx7dRglUG+3jC9j0qJq1JKyp0AoTOxp0C
ibix3cjiWEoAu0nu+pPz4/5wylSX1e2yOxGwCzW5Xfs8GOcdUtkSrz12r9+ljVzi
DBlanRn3KJMShuQva0Ks4lcl9ojCOTLQQwv+llSZdJG5sXGcPRV+6SULr5FajfWZ
aEPyzTJx14Bmv/4RNTug3stznHm2bYxNlXfGftT/YeWlo8avcMobwW3rU521Z5XC
0Db0l7ZE4ksxutECKDY1Kj/rxEKSSDcixZzljva22LtwXdH+uqq++3uh6ha0igbe
21NH8G7hGkkXMzEBz8msJmV5VlO0QZUkhEjNPLOzuFPjGAD19khH/fqIQHK4mVLF
We2uxw1/PiS7UNjGU7eu6s/3yLHdpl+8XE05ztU8Cvd2vsfNdKFR/91Zg7YVts6W
PUWsnjNM1a7GKUcYgT5AZhCcatdYpWXGEljwqsdXHHsF90kZDcVu8gxD5kdlFt0C
acU3sZWmlB4Xw/GR8nBawDkFOVZ8tvwMfeGQgsig6hKSTyAz4BZ+voFNy4gSlV2M
1tTw6OSTfGcmZjM13PEpDKyBE1H03c3rMbb4lma4TPwjKhjh9CsGQ9+cSjLymy/j
ReTZbqSodMGaDtI+LcKYaQ6d4qtcZzh5bLsq1yBujwoUeG64bIZOT1B2Q0U18VaY
AN/3KTkwo1ep8hS2lWSA8J9ud0pTfA9vKazYQ7a+UWoDXL2Pk4Cyw+0AtLxl/I9P
U4RZ9hKb9Uiw37Q2yLheqX4ZjFWp1W0yrBTYoORN4AceoeljDKiZdsMjaL1mF9X9
1vFVfnEWSpGECfWIm6PJaJW9PHsr0xmsJNo+9kTHYoAL0fklE6ZstGo4vBQ4cJjH
VGVerPaFTjn0Y2MDnqSnYoec+DKxD+XOL8AWD99XljDSKURNlLo/Fci50NLLsJmd
BTeRWTM/gTvIch2g4ezgc4M9IW1Ldsvw2hy5A3Xh4a/Cu8hf2cmohett7rMY/Qsv
rLahIFU8/VAIuKcI3pfZ3A9RfBSbSb7ESvu6jQQNMbkgSaAlnh1hRfw6VJ1UVUda
AsOprQCoiaEYOIVbSqbAiDXpFZkHX6U/pszjZlY/birxChWChiRhEdmB7b0HCDUE
NwoXEWfMN+LYWlOZWjEaKodc2E1ChlrhX/X9NNl0Kw/jzZuizx3yfhQt2ouiR0XC
bhBboNCiOQ3J9lKdb3HFU6RMwqkpZrvLMlzZfD9iqQe3xQgffi3Q1jS7Vp0dl89Q
XLm354AK5DIhbM5SWxvD+4ejtzRQo5TuHcGC2U+Saw5hT371snC1i4+s/xhJqUMC
dlcPP1junOFJP+nnMv2fwNVnnSEhmRUevr5WRFNympR436F7VUWb1ZurfFJJvp/v
4g63ApvvpJFqwpi4K2+xOpXce4qzG7bcMxdB/+BBCT6vSiXVt226HQmCE5wGorA1
AfXaUf+P1klinTslVKi4+T0PtruHAnaxZz+U4Zw9sQYMWLZ/7mEPWfrBFoBzBwUx
LbVc1grIzbFLMFOqEmQe2DMu4EcQ2VL8T2TRZIEdTmM4HA1OPvVn76cjsa5TKlYg
+Z3LFVGcr9/FWHASVoyrzvXgv64oGABSpSDdw6vNx/lOcHuOYfGK+XzyUUcn9A3E
rIj4dsUwegluxqbae2w0AXj9by5xMxoXOo871oMgW2Wem/7r5D99/2cA5biLMSqO
F1WslxcLxm36d3U42qGpDndzgO11Pa9bZkVy8ryP4/ILfNoSSeJn0P+8/6//rTSn
XJoAkGaYbCcuG5GUTt73klangCyDIyv1ApaieMlzEp8UiK0zBxJcIxWEZ4bzJJk2
Fskvc8Q3XcuamNSnGheGSoC0lwpBmg/DTNxamAS0QQO7FTxzXegb7qpxC72OOCiZ
EtKAkaLRP3JRblHsg6wPkJ8WHK9f+LrytQyfflVQJ5Ch84UO4KFfMTn4aHQuIKv+
0gcNjCXyVfrh4/6Zkd4NDvkTC1f4B2kGKjXmYLnaEismQ2JHlDu8ehw88kk35fp+
T6L128/wM4gn09K6VHQhyW/aeTALVJKm4+dQsICsZbqrtD/t6rrlEB6o0xAoRHbL
YFS+izUVE74bAmIY/xImzmwLYYOv56mNK5M1wdADMHSdAxKwZXmkNbbntea96hdm
xd/FML3qPkP01TqKVjF3VA8jVWsDdR354a7MyxAhytrPgWtqAbNFvs+QU1Bkvgn1
OGb7RuUH6eXqSMI2Eg9VQztNrBPrHZ5mVOwoLsHHneALiK54iri5el3DRR6f1yzJ
y6CBi1LV/L/XFtx1g1mgCuuX7dBKHkmU4/L1Hr79TRiPtAW7q7Q8+W15Q8mP8NiH
gIHWPtYaTSq7r56gfVY3ac+zBTX6F6Rf7hNv2xsJWT1t3PhM9piUx5gQRZV2I0jr
v+j31GlQaVDmzT+BOFSJQxa/F4BbGGTgIIWn1CPd8PY9bM7WCzWqhRWRNiDla/uA
/xQjUBMfGTo4b2qkK9WUgYkDHX9odDXhbzBhHEiXgniYiWl64gRGU2jrrziXiYR0
8AYwK551azpz9IMpOXk6ZggUPnzmyJwQc4gMGdV+m4baR6wESn9qDPZKZXZqtAJN
+FxXk72RUvGKhAfx6NA82Bqu55sboCJFxCFOHMzwrlWIDp53+VEenOAeCMtr5s0D
Pgc3xAtezfUKVmc+r6+1/TZWfT3DWbJn99crZq2QVLiTmgewJlyhOHfsrCoo4rD+
VI66cz1TKJqM7Rn2lY5UXMTyuBA/qmi7kRzbFsNpezWyZyYcX64TMTyDjyA7sOmr
N/JWNOaVBM11D2UCgomqsuiTkjhGZEbAzgSFNM2lENNfNnGGp+9ERjHQ/aGnPdjX
cp/4CtkUXfmTXkwEDfNjIxczRpXw5Z/PPe2Nf7v1utwpbAd/DfrJC4SkQ2tH4eBQ
wGWp7elR4XCHbCA03vEz2+YxRMdNlmy6M+QO/DM98KL38DcHrHEuPOgPNrx8w8bw
H3NYcnt1HbVNxIQOb0f8jbtVnxM5fHg5AnfOGYQfTXL0iFVz+gkMzUvyu2EmqeGq
r5m44q1DODIJU17cZ3SyDQvpUqXSsJOOHlWWyRAUAehlLS2k6QGz1/vHR789wnZL
7FXvvW6QA+VQsmtthoRRsrG8gRbDMXl3iUGFpBlRgSEvv+yrbLDBiFaHlk8K891c
b4clostJsHmtdayjEfqqkBg/jVdVmE5PRueEy6OBO9QVPZDx4XFrkTFc1BzkN3Zx
epg2rek8KtSE1Ly0JgHJe+AaGkstDA0QbNnXwHkujKvgKW/lR6s3JSrIpNb7ECfw
aEXjZuO0NjXcPcNM7JmQA4cinF6CUGCV+Bxcn4sU3LN9S5DPAD6CeEUy76qpY+S/
HbzRmaXIrDfbkt4A7nO4IY37Imki0KvhUZwSHqu3QaCYdTU1d167RYgrk5A2lZa6
Cn1bbBuhLUWtt0/bv1cRnFVa1XJYOov664t7txlMpq4ZW+zxtZts8NlgnTB4Ioi/
oqTe5trIXCJ7SAMPBvY5soRwS9HXpfxTOAR99FsKjjfOvH02B1QNflywDTs/9KdY
XWsPt56iySWNA6PxswSbyMIG4LlJQy7mK5DNxnUmmv3R370kbOnOsmn2Ya+JJi7I
Jdh/fn+GePpGYSNY8lGSLBWq2kL1g7C4jRIxSla8UgQGibe90bYDVWmIvSx5EUMB
xGnzHp10Jox0Ojcf9blFufz6opJFSanCeTToND0KL89tAT73i5vlmgBgQKOe90wP
ZuyGwDzlcyx6ftRcUXLxFnmIog3YDNOqv4wvw01THQvEbnYJafU+41hmWUPXJi3+
P/Q+kwkPaQ6Z/rgYHunOf4J+9dP9D6bKcwuRMys8gkC/2/uJrveTBgj7ULNvztu0
cscHOgRKWdutRVA6cixaYMDlidtwgGyqKDNgdNJc3aV4txk565azoceH1iXfqEkG
ehPuS4Nsu4YlAhjUPKxlQFia640Qq58WYGlFYzO54yuHHcpgyUHn8omb0b9HvH3+
W4giUrtr6MmlbcEnFAK86Ote8b/nUNQ7lb0/pQlcFR7rSdc/sBl/4GriptVK/Rzf
VYJQA2yXXTJ/KMtLO5Uct9dMHXYzYnI58VZv4wl1jkliOY7BNXxPAjzRFGcNJgdF
ZfDfXpzuD6TsO9hc7S2dOLa7uaE2ForkN+MAzHmZDfdL8a29TXlMPGXfwXSXoIh9
TDRtEKntyBrzE2S+UUBf1hI3s9nAXHfVDhJsf3qO6dpgSJH+80aQ++413s2gE6Rc
md6+OUgT8d0yQQEir0axRDK+YkkKU/w4gJVBKzI+MFUpcu8MSCUXWdKEbu82gr2c
atvEyuRY6+JK4KwWcd05+62ZV2XC0rueFtSVkfnhbjdVo59GigvnonM6dWKoWtKO
Eju+RtmzURr8f0gjy8FzV4UbZEHw8JC2BYO8KggihXLTbNq0IboweGgDi2Tt+0+L
EkwnEeCBXnE8REtTaOlZ5OC24AQx0B0EswfmwDP/EW3ZAgILxdhAZY49D8ODSOP+
beD/48KvPlKIxmQAIWoYMZHoVh+vVLUNe4SHtUqSeFxQAYhNdxJNLNxTeeXwI3fT
l3+8LD3qqj/SG4a9+zAUFeU73naKd4zvJ8QUQJ/DBulcnWY5ccZXImI3+7LyLvD9
nOuxcDbY8bkG/JfgFk4tqcj7M2k7C2rtZVXKylIm3Q47ChVBIhZ23RWNX6oSV8p5
u/1fTAMSEbv6mFv7Ns2m/GVaefozV3ZHYfQrdco02xrlKOEFUsHanIjsQq5k3roc
Lq5bxkqI/4lE1Gm7Ym71UovHaal4SBz6Yg8EcO9ztKzc7rECTv3seGusiyrB4206
m28pxlxrTyz2WBtwo6/tVrPZy69gSSfIcD5UyTGCvE4aop2nF8rpHxvJJqk5cdEN
VrPN9faoAUieZgHWtYKvP6Ktrt19WF0zN+14WQophtNejGK7oM9liW0E0RqeTo30
uB4NVMkpe4pEX6ferjt7i2mVTB1zg2sWSAvg2qspUpbtz7eIBPiTr1xkL5AEUe8R
O6hi/iXWCbVZhoZ4RAisUkb/GZHUMunrnEm5cBn96Hhsu2PqUlOGDMz6ARuuiyIn
/qIBv1HbXfuspZ2ZkIBqkQbXk/N0ArJKi2MqMiKAAHlm3NgJGSWJDkO+nEgGW9Z4
eWMv+KceN0yleUPfnFn50FNVD52aabfrpLzA9cNjl8OWI420Ovka4MWM1FSi5wqL
s7koNdOBhFakacwkDVVZqAxrHkJGXL0MDW2X5v6r9qESCRyph0GlVq4qvRflGXNO
LukEBajiYXfNnIDQO7PPX5XzJtUe06Hy7CSynoIwighlX9eqYiGuVd9LK0jWeTvy
XAhcY8CSUFYFeCGBEq7VpYltBmYkMgtqMCU5cpczBSMvC3VhxW8xL8vGG6TIGn4B
vfn3ORb7A58WWPjx42gEdrFCD+sxuCqY8sTmquTFRZryUCZZBR/rFgB7aQdkEy/1
30guduFzHOEM+Ybf/8ci43o4cYIaJTR5xenQeKUxmbu+N0HoJOVZAXCEVIveEJlK
SXnOKs6JOgPoRv4alhWu474cJ3wkEKZnjJDPN46pduatMSYduQIQxp3qicTbnkG0
T3UscXHweTVOzUC47QHs3eOC5Q5+1sWiP0Jv3qg/SOYsS2q9qJlHhYAQkBxZE7By
hTBn86wjL4aGEAlXkI8TvZM0RNkciPeNZI4gyoaNJSZSJI/qankpGBy+Z3ZZ6Yn9
crNH8lisXK5leQQqTiTIV8+Z7U5+8iDOcxur3p1YOsjnqxQY+kl1iKMdRqSM4UIo
Kx2EWNyMd2eVaodO2dtCYraSIVelTltRB5+xrrzv4K3LELlxVp9AaiM52+G58Qry
+aNWCC0w72Da8Qt0gOq7yxS1vNIrDr7LOYNOimOxFtR9LIENVZPziXEI2Hz02v/a
0/0cPa8RPA76r7fBHc241qQ0IxbdpylOeVmw/PuKtsuDIN/e8NnrcitZae/ZSGQN
AIE3ABwVos9ZSI78QjQon53N86+YW4QIaXRgq81ClZbNjBilEmfKl3IDDiGiz2VT
e/TfBtVrJx4VIqvZIPUwWuP8DQyB6yPVqZqCRW/+vkfW8NtE/FVsbwgB9S89grHH
ksWH0kLu1FFQzve6qiUlCl7lNb6uItnDrS7UlN3RGPto+OW/7zX81R5mz5c9WKPE
G8/fUsBG/xGOEsCBPTEWhkVOGOQl3y4AXNcmx00+WfwmE/dQA4hiXhjxFwQcx6TL
urJ1f8gysr8NLS7dhMDP7zbl2Vl+IeXiH3fMFdFk7+jZeUw5XR/t1JgeZvxSl2+Y
5RDHPEn5pW1Qj8+367H36dPmyKF85GXNnHzTAWPTpMqD9Ty6csm4h915lUN6Fbtm
90QdyMJQTSSkRziGprEvRFcFlw7+udFa3VYYLNhnI/6wU/EcwFf9l8RSru6z59W3
7jQ+PAJ08C3PGh3JfTKoNevniMY4B1+9UI0Q9EKmU/trgSt5YmQ8Mfsu0PDuTm74
kMRbukbFwgQLA3q0RT3S8DZPoqHDyJMZqFzUDMeyPtP1mWGV0yIoGo5gHjbtSM8z
Zmk/5xjxzwgWEa9Pv2tGjlPGY8t1fQSlEVw1pVLGWlJetDB02BQC9J9twukhrIEy
8m8YK18YcCq8tI2BcW6b0HoYiywvlKj/4gGpTUMowR8M/xaxHjW7Ktt63gEBVVH4
XDSZBZYvJwKhkOw2DtsKDxDH9NF4j+PAb/sZu/nNg0KlqzAVqNfoh5Rg35uj4LSo
c031NnBXi0wiM7k+ZF3N24CYxLzrBqtMiqVVcJ8Aod/zv1qH6xyDs/o8Efv7DU0G
c6rZF3uvWBTTOOhGzVopX9GZaENzaXBr405N50Y8akYF7AnspvdmKNnougVlqPf1
t8nlqjAgu3q9KX2qG1isbzyUYXJdLgATbYdcc4p5y4sdpz+fDah/62KWtpJ0/CnF
KphvC7dliXdReNpPnslRB2A4kXrkVlCpafLrUpe3Pl5kDxPJfSuCr2WFIr/H1WgS
1i25dmrVnbixkS6S++6uFzru00/CgYoBodrxH5AAzjk2DTrg5MgfGMJw/fFow4w9
A5eexEYhVXP9UQfz0QzMZWsKw7zlq3KUyrFroWVaLrW/uU2QsmhWhX0oVYbjNDcn
dLShbyTWeejsbp0WbSEZOAjilvSZGNeeNvYnk+MmzGnYvzK/AV3dJoOBEjDPRhzf
FkfEUU7lMiJt2bluo5zb56WE0CF5l+GXry5QaVd84DdLUdSf3RyAf0AqwaRLpMtk
31d4c5gABhClDf6741kwD8jcNBu9lrrQoJztSa26S6JeRZEARk5Qln16GWy/Ye/m
nR2SKHbuksg8lKi0CCR+m79C/M8HtuY7Gk5RLtbpb5l/+VqDyadnoF2uvpKr2o2+
W77ZoG8rQdlwo8XwajnfibArLFvyVngNIM9zXhFRMc+v8VYBWK35tIWtAzNSWltE
NuECEhGTULKAoUYY/IaiAQlAt21x2az1aHjugE+6wzDXB3oe2bB7OjTdGIIivxS5
F/JwTrIQu4jtGKIrv2ZSiteGY/wLd2eT6MkvUtoPZonEpn79mVkTsdkW2T8amsGF
xWAuwvjD+YSe2F0t72E88AyXDJy/kb80O7tjMMpc5xIBJ0yOsWZRNFATJq5fnAMw
78ulQPV/WHqmjqtUMhpbZizgTArUwi7llg9HX57QOidl2g33vM3dI1uwT4Hu17rm
e+ylYvzH/FYwAR+wR+XTY14b8kOIyox1sTDZf5ntSGD6bvVBtj2MkyYZPs9eRZYc
WnUPt12hUE6NXvuadDrSeBzx/s6GTnH6VzQeFf8k9onFU8BegdWR6HbG8UdJabE6
lv2iGc4a23cK7MsPnP5t79XlwB+vIZ3l4FHGzZVP9VpcnDHgeGawJ6jr7IIlaz9X
TWPZNOeDM2NLMuiFkg/tpYrqW1B3rksh3i4QskVeARWdb7Bj+pqQnCOt6dQ0LXn2
xUEYYO4U0gSh45dx0H9btVAAqvsmuxBkcgL/xbawzduhymg/AYIF+K2UHnZLzr6R
FCRK13urzgKVb7wvnZ7hA+4nTGx6+dq7JaKmJ3BrDuGefC6SG9AWpI6kGV4CB13V
kAwBefSBUR1ucsadxl6ckSKCgA4kxDCYcKcI8f5WaDOfTG2EWD9Fqry8KQIB9Vka
C98PRDVloHLEHVblFQ21HQZwMrdyzUXxBNcrNUOi1lbSuThqkDltp6knbSrcVt1a
3LWw4EBNsIxT2Yy0XL/QKO59JBbyQNdOiOQxnb7KMgVhOigzvkIEjv6snIQw/+F6
PpHEte57CM+Sd0wlxh7+taerCKqdUaKALqBaKzMnkxEsnQb0H6caHS7iFTHPW6hP
s4bI0oES9Miij3mZytF2Pb+HNzVuUV7awRuJqqKmn26QCE8ODoJYWfJTuYB8dES/
GhsX1jwKPjfk88Pg0sGQzRl6Lsi+DrZfL4eCY7BS51vOHDHmTB7PsC0IkdtLBeTY
+fb2q/m+XtoFPs1zP2E7dDs7qCqkILaACn+fbkWq5iRmDDTOVAHxZLtfMCmMPS2u
DlXzLS/DM9WhWb8HlGBclmiLRncz6GT+tCnGcpRo44gkOAi8EecJTNmEGmawbBjw
8XHZYXLf6JVQ01ieyPRzjgF3Tu/myGU/rAylgyU94tK08iW98aFfEwVMlSqb+BQH
QSnfEQagIIFfSQE6ltZv+4BzpkdapNysrbHZuEaA204T7mt+IIItg8OImKdb95Ac
nHeDQcQcgU2RAx1/vbYAH6ZfWjWJSR8eJ4dLCNj/ljYecGk69zi041P4sc2Y5Ufr
Vww7KK3s8EDrkFvH/GeHxMGjTBTE8mZkjHGfaAC+mlQWD6wXULv6zgUAp3iW6rqA
ze3xYfurUGzTtt0N7IvAemiYeY4GCgy7AG6lOzJlHW58NzdXNhh/V5TUbdmZUPTn
GIV+4ff29CNrsOPfwIS/fYGFBeWdUAKj/4/vcvxrwNYRZU7+9F7lbLBUNcvgmmMN
5B1LGvU0cc4iV8d/oDasmmJhbK7DSKrnx7R7Qqy5DTTz+UtCUX6CdFruq3gDVDLR
Nwr72SlALopnR8LeWBUWt/7tCNYozIcvgvaoxL1u6jqdQhc++iTroiVUJOqFQDkj
Zi+vIhN87AlZXxofgUHF9C2RhVUwKSD4qla8hHB0bLRyG+sviCzgM7XDnbAQmQ0F
+XxO7mGaddUIqGtMx5nrp1u6d3ZdMmislKiCJYAOfeVOZ6KUTtv9Sj3LR5vxH3cM
9e4ViE/MoilLe+J9j6hghlVyE/j6j1j7PghQZ0Vpv+6cOycZ9kbQ43Pu+DuM7xNz
RcgGKJenHVPudpU5VoLjTndHHjF1IGtoep1PemIpRtuFpONliHzgAjxEO4ix20/2
TTohBMQRnvClYldOol6H2x6Kw2FtoVb3I7ZW4MaVUGB2j2P+hY1kLW8UUkK1JXtk
i5+bovXBtupXmyGq19fGenj++H1bTwTd6UqzihFBwdzeETsyUQzhruiVBumgjc8a
0SqzWkXbnUgQ+EuzbmYxow/R8HfUONvXTl73BQKskZLIukMHD0N2HtAQPBwXQz7B
bkrBfWtE2hEYe6uBek3fD3vF2UhXg0gwYs2oYbWcxhNR1GsXbsajYLyp+e1Xv6NO
7dIgiV2nxjf9dPbGUf9xFy6V6Pp2Dlnb9OVclcTBhpv9bs8C9M9N6DPKUjYG9GPD
CH9VCs+lzW3lXPxALPsChIj8yoPEPde8n4GUbgpT1AFpOAcX9c/LAzInUHXBonfV
ArHF9PPh/Mbo+prC7HJWH0YhdpE1p5GVt5T373tp5cvk3d8oDvRQ6hncAYuRME5B
DMneBwb8YDWrqWcYxo7qROHbA/6NW0CCuVQ98Ld61y4/PHTwdl4vQJVcIUsMK/Af
ooiuBGnCg9QGvQA7Ow6INNGiw4WdxXVWaZkIxHTG+IehoHNxJbn7R3F+zjvgIsfZ
0YDHPoCGo5k2e+8c5KtBUuKJNKN4x/dxQohxLcS20Ec1wddPBbvh3Jg2Jq+fpmwG
XCKmg5KjBCnSEbNiTnX0c/YIzOQq/ESt88bWaEE/NY5zUT4Rmo8gtEtPqItZdf5N
nGfJiHEXSF1waVNOO9Jiq2fXPUknP0GzjITui9/c1rmtfAaDD+MqY5sJ3RLNJ/Lz
zHKwwCXAnQHISrvpl6JuPaWHajE0zee83/XEFf4xHB0vDr4KWYFTOVFi8uvXPKYE
brSQAV/ylHQCapQiq9ZEwK6ktR/VNmhFR9ypxjV38NyJFPehxkYl6Ft5D1swqjEh
ibQp14CRt13lAeOq5glC8WlzZGUZemLdjc9TXBBLMh9/PI8rGaIpckFyGbrAVlIn
JoqN9YX3IQmXpZBvBEnkrlf20p2oUHBs7+YcsHsfTn51vjfKCrKhJLrtUYXF7B+c
3RHYkswdGgxtICErpJORxQEf+Q2v7OY03c7iDKSW63P3X1JApdzCPpuYrQXqwxqA
x2/NkkTr0KgYFPtrlwOUqOAqukKTpxfNmWLf8pPddmF5TYbIjF2vL0ZlWeglA9Xz
hZY/wHo+q6GWLkNCU5W7nRkKThj2Ee+CtUH7EdDw5br4FaDV6EiNKvE4TXg9XBDs
D12e5HIaKvV8yZhBo3o7Ez5O0lPYFyVpT7sgwImIzs+1ccYqn0+GEaml33x6+9Lk
Q2NdVa7kU8+xMJSVMhfLyk7vlUKl1Z+6NaffRCTq07idszrfbTXgHc5jJaD4u1Tg
60FfK0rSRftjWtqrXn2cXuwyKV23t9D5NB2JeC6SAyazVVia22cEhgYqAZjipBy5
l/3TuykCW/UR2OzQNIKWH2nlu/dc/4LNFreFvRzEo74oD7s0X2o3+wurQyv2ARLF
+m4RHcyf09bHuczgB0TpYcsOVfdH1Gwt8rvbx4o7g+KpPInb7CJXJ71DNfuG1CgC
SocEy4f5tb/oUBEGKE19FMvNC5XOD08ueBHcCgfvf54muGq7iELV4y9w5OgtQCUi
dYd3zrzbGRo/tjN421lOXun4+r1vxWFeYc5lD0n/MWasMzLpW+gAECTiYELCUzTL
WiLy7hct44hG/Tn9ib7BF6A63+fx7vTqQEA34G612ZrUv7AQVYbceUs/1oi0J9Je
iNEMMvLvQBqQjwOCaZ5OMWc7rW3je7yg7m4kQDQBk/tMYgmZeyg5JMkDw+Z4KLCJ
mEyJTImzsljuewElDw4Oyamg0OO/GH0MIObeURmTkDyrlqUGKfVbWjUBBjS6Apk6
6AxiFqrn+HPvZpmUhT+gdPcDXnHPq4+bJr9e75iQ2jJjPZdhhHSKqRndB6FSm1If
VJTZE6OdRuSyU1ks+P9tRyejdeezvZIG6pIlpBTob7zTkIOLUMpD2wmkwASYhGEA
0a+29jhVW8VXioH/+ZDZ2wKOoyfh8KdMOjhLCF1FFjZZblXneUzBqyRyoKZ69o7+
+CCiTUHFEXpnvF9Qs21boYMLtzXKMudn0aKWRQMqZ8MzHxaXhvzosl0y9h/434wx
UsWls2mZ0Esgc72/ZLElDJoOci9G5j5yBdUq8ZcFAzaOvGLZco1Kt4tM7eyxDaK/
gTgToKjTf3Sku9tjP1KuCI0wWI/R+5zMnwvZfKYdTYHHiYcHe0CQiwQ4Z0DxBhj5
wnzy9/8g7gp8248zUN8ROLU6ewOT1iv8Ymxsi/kX4fNGtyB3RexeoqpNg3ooqutZ
n3eMdTSOvsdWklabndp9yzo4/nrtyICVjJPAcdl64i3RnrqFupAhNMXHWIGpW9zC
kEpO1w4g1yUL9SSw5Sc0v2sA71ujSETv0i0vNLb7VOy8ucw/ni51p0ugLV9OsMNH
vdfx1tG3zq191OPyRvXKhxoWPOLSs/CjcR70FKeC5k5PLPPqkcZbk24WmGm0+Ii/
3+8kiscVNKw84qLZBCI5vD75Gu/fe1aReiLkOrWWlzvwJ+Nnt0GozaQkyNBwiJPY
S5d48O8ZYahr/KmEBvEA7uy2jFmeZxuRB1i/odT0R6cQ1aK3wg6unDpF7KKKEZvs
u7AV46mcHrzR8b2FNFr6Z2QnbzjE1w6PnPdxaVlr4Hwd7dCJUEy5dF6dKIon+r3a
GxozRZhIRat1H55+UoRNftU46BDL7NK8y+m9m8Zp7oYDv0K6j6FVBBLDEvNZMq6R
R/EAxrWsLAl+GejNoCjOg+bp7rbAnvkQRNFxK96YFDYSBwecqv9v4ZDU9HE768VM
NMECQuFZzts0//3vLP3Oj2tpFe8nDDQB2IX6320aDqVOtCUXFzRbFO1nb1q7dcQC
bKOKej/yOVV4mulHYBEsrgrTJ58kFr0ZVOt8zV5C3vwyhFPp0y6ZD2tH6wKUSLxf
nSwZAEcK4eifAfrIkFoAZiGacNiCJlLZj5Zsj3LGG+3J+6TYwTCOT2BMxLQGzaTU
sAxrDxEpVdfc65YUwYWO0i6OlkkA+ZVvsPUnmjLH3BdjCyF+5JQqafxCrpok3YQ0
KFWqmBbJTJLsh9w0LFEZeOiNuIVyoNNs90n6bzKy/lKGPkHgDKGSBnEOrF6savI5
UDh+8/EXzesohXi+tsOut5oJMXNZQdpBCtrHiZ6XLpKG6onY4tWSXZZ7Qo+g/Vjp
y/GW8n00nDGO2eEEW/cn8njOsKC0weBl8TXk2Pmm5B8d0IM6RC0dy29S2BeJ26pj
tibA+cvax+wTgB0rAWi508/un0ePcuqbBD/JXzHYwidCF4eHq3Kw8ei6Db2s2vb7
IK+3t4NESputw61pyhqsMeDTeity8aDIehngQcQ26dwLoYy7R75W63Y+5dGb5s7j
FIY25y1m6rk3qWEJ4qVAH5GTrJDYQnpb6KalPcDz5eS6t9jBmzz+AOz/JpU924gm
pNvI2CzK6R7IVuh+OEXxROkJYFuxctsrmMWrCVG32OpiOU+FPfcbGFb3PRPiEYdv
Iz2Z0R8vrNXJVU0K8UG0nsSVfx985e2Y8rklonJPQb9lQgcm3zIjmfimzlVmYxe7
eVxqrAc9jr69nmqtjemrfdV3PODV6IqxMKaZ8CuSHrJ56XoOom0Btjpe/Ja6EwjJ
6tdZHfDuKMk4qXRE9mVhZL1Ah5ay9EYBv0bbKsug6hCatT15C6FsylTLlGxjRn9/
CFkihekknyLsP/PBLu7MlYxdMWYimiTqxsF9lbdtQChkr12WGzoGZtGnwSgHVczy
q7qQWP66gcbXfqYyiFP+WU2oPEz6kCZ4YtqMAM2fU3sLmQ5M3eEUcHJeTPaW4ik9
JgQBXV+wy2OWsq4S8Rh9kPCUfUSqHO5Ll8F67KzzwUzWTbauyInlzpLzZj562V+w
e+9DdlZwL8mtB16B7PUqb28Yb9cfp6yfHu6I6SltnJqnRLdI3eble4UwmareNJ2w
htECIz9RaCmd1u3qRZ2qrJDXlnyDmJD4Ka/h1pxPJob2fqzxdrsMs/hJKtY4MPSW
qceqITQDlm/tqF9VB1+ickgcs9wri/FmBqiY9gJElmMi2KDGZtyOedoYcyrWGL0v
G5rxhMc/+96oV+JgERdQ2jI3m44Xf2I3pxCXQ2Q+2lF/lFzOQB+fAMXNm6SFBYNj
HeyeIhvCuVaYl6IlYUQptTOtNqCuNiHBgoz+J2JfVX/VdTkTTrWbk4bGX04D9WcH
Vkb1gE/G63tNTXY131WhzhQVAr5DAG2ssAENqXf5z7mthCffwkyFIfLTeiAXFXIT
5hkNDlnkBd+ZFr93VDuQsmNTegy1U846Kol6351Wta3C0g3lNV/PiiH4msJVXfAI
hyu69sy9ik0fP478Af4DEYclemiUu6SXAAzq0NkB8ltb9l6Dg7+sSHDgz1DHxpAr
teeMQP6kb6uJTxzYRwwM8ggxTKFsGwRXZoLhHMK/0KOaNRx9vft9mnxj442CvDlD
CyPm7TW4mpY8OoABmCQ9r2QrhGD1yRXi9G/wIlbcgvJPuKV5f/R1qNAGICVjJyqu
OcOpOB21R9+2tGOoKY/EpjS20ArCQ8d5vtrEqAdavwlnP17Dp8JDLtlCSudzwQAD
aurBsevLics12dqRzXju9N+ILED+cHSHutWCrpFRWVkgQqy0MTeGFnIC9WLARA1x
siqVIh/bVDqOk/RyFVUGkofFcvSfcDejpWh1K8vMfmWrCIjRx9LZOGcQPUuLwYDF
j9/EYKJT8MEjK1LMRdZk1vVlLopc/fFdaKOfP2DkmPU5OfFr4AODxeudnhfaw5rk
BHEGL2pY90JX14m27KBd3xfmcwx3FzfpjpaXfutZ29W8eogp5klyy2EZ0lUTnFoo
Uib0FxGFd0WqmYHG95hfvT9MLd3dE/OWlHL2AMrq8kSWkAAkICz5a0ohOegFn6Es
12o510wfbtsJNK6czSu4CV27Oh3JOZl/pRpy47M3itaPq0ZglYhQzDBg9r9vZX2c
5bMdWwC9WdBfygyvk/+Ejt1C5+gddnh5dnv+PNGw0qvnzprj6xW+f+5X6LXL7G02
aVL/CxL56axPBJmveqjUlWeBgLt5GHYvbWV6OiyF4nhbjsma45qgE1ZmoOkq38UV
baONGFlRacrXAD3JEtGOnGwqHMsMVJXMX3dxSR/q/rTaEPzQZHCzIlkRchtNPFUI
gMCyXQYHVPO8A4L+jFZBUrOsEN0X5cRW4maWrJaS7ogF8v8OsSUbRYNo1SKt2BcM
karl0dShu2Bs3D3tiU8LYavgc2WwTONuZ4LfzsjJlJWs8k18G4ASNPJGfY/YUOWn
Cl4t7KU6hfdFcKVO6h0Y+b/79wY50bg/p4s99yf8OiZjZuMYGNfshSh+4io3jxZW
AK8lOGGqRNcnWnrX/iAQPBnkE2OIbxILqNt2G01NtpUM8idT91hkS8uBznei7/io
RTvylb5WLKAsOMldCr863BQ9+2xcnwxXvwNAAGARmEcwoF1S4SmQCW7js86dTiPU
J+srn1mdseuQP1gv+UkHZpJZIb6i1gWCy5c0g8KSZbHDu/IzvSpFkDeOQ1b59ksD
5WJN9Ih8zB1cFxCPy3NPqiYOZ18uoFAHyU1D0gS6JlquDw30RKBa5vP6wbXddY7D
cS5rNLxR929JvqfQoC9bYZUPn38SZgt+6cqexnDuk/fto/wjI8qORGp4oi/EOE0G
sFZRlWy7eO4bUNZPT4pr9b/emN0j7o7KUHcQ5UCePc6Jc/YsUJnA7GzWULr+/ROG
AsSOz4S6/jBAapm5/TcwvpKYBKoxwtMsykylmIET6qNP8G2Th8em3ztQGBWHizAM
5cs+b1AdsYZobfWHw15PRJ/TG0IokNdox+R3lKaMnaqGK58ffsN0b4I2D0T5vrxx
ZWyXd86Ee8OERYtZWmh1xMphY1T71jcPGotMXfPw3O1OUTL3/GWKo9IkMrtFKSgL
MpcgPix2EQk4xsXsVz/yrm4X6YrGO5iwHnbI07hSY1D+fG7McyDm0PtV9aSFhR8q
vCuzYfXBYVvqT5GTP9KMp9EIFoyviViLDICo76sBoRs5jiM1hRU9lIEdiUG/j7gI
ULiL9aryLKPJTr93Wo/ifv5teeLxwjhOcguHYqBCJdzzTmFJqQK2PskszxqQBH5l
PFmAAUkq8ibs5n4F8Dp7DsUqopUiU6T5Nc9QM3LXKsmq1p+B9PS6Oauxi07o9jYN
QXinRJ1VWX9QS+BjuiElpQ+SdT0aD8xZfnNIgeT1PlcKtvQtWcP/Ku6+Sr8hVb5t
YID+jnAre3l9AX4BTSbrWMyN++9k3Ter38ZixgGW7/rATtcuPtd+I05jgA8Nvu52
3M8VBqjUZtYwRy8Nb2smOW1cs8P+B0CIEvIims3qwH0HCZz/aeFk4Wg3O8hRArEH
OYWxnRTZdUm0AfyP6D/esSjIztyUGaCFNdXmBuFQgjl7gqYV5j6U1CQbm9zBiBD7
DTt5BD6D4RnhVtJfzBAeuh3UDKjZioOQ5XmYE3iL8tYnsA0fDe/HCqtsH6WbTCCb
omzruO8Uo07hFSe1VHheLVIl259Guo1LcyuxXlADdMmnqkVsWBPdU36jgxcaK9Pv
GeqQe4dGJ4/hn+3z21HhfT6SIBXlF7RTFN5NEF4Iv2pRgvyJu8m2r+JM5esnn4t7
t731TsYJ419cuf38d8nfdLuQoEfo5AL7ryJ3LVbSim8A/65zjg4LUP+AWRdonyGF
Eci2fkZ2+7tC1azM+jnBsmnOPOpqCuBIGPQS+VX2181DcRuZXyyeNbQNqtR0s7Io
aaqy0nXG/59oB+c6pPPeMJEqWOBfH3hAOMSQ7Qx77Zf93WFz9jU8dYRbApEqaFdN
gkULLRxzlbWCso/t9jNO2s5j8Z0Zx2kkhmepSqqIwClNyqqwTNg2PyF97Ez+S+LB
VQ4aOKkUZmkZX8D13BcoTq6eJ2PevTobXlc99Fk3L9bGvsmpZys3GQzWtG2KaIBe
Dfe32nAm6GFzpgTrsRJATm6WLAoI+oJlejcbFoP/bYijrHOgzE8R8gJ3J1YfwrIj
IKFk90q7pqrIVXbiRIDwUnqFW3LNVbT0LeeztcjLssJAaM7/kR4x4U23PRY+58NH
onhnrQLqLTjO4aSLuusKUpMO4uiYHYlM+brF/eoYfr0cAOWNZsaFxXu69pcpODof
8mDGQoxHz1mOFyK+x2r71trl582b6ZAZnOLAxddAmtdRuUyTjZSvPKnV20Q3CzHq
EMatKgq/FSFgtJK0Ae6IfHYCFqXTN/pJ5hzrcWZtBKn9fb6+oVKpZmobeVvBsifv
jFbBKNIT44FCUEsbM5qrVhvzplcQbYfFwavGJJ81NlLcvwC+muV9qwEFO42To480
Rm6XpjeMpwqT6EdED5OQYyxJSKrCNKT9M6vHC3Xfs8c0q7ftyCEVAhLQ4PQLWbcK
oXIbtfz7d0XBAnbeKHsjA3c/7vTdGm2LrZOR3ZcC4JuNNlkpMd14KkEnbKJM/1DR
dndB/qTXzju7H35sPG13MfXlt6xzvACYyEX+qpwXzddXbXaQ/FaAYacrMG+a8KGb
HfW9wziN9gvSHtzBb0+MqtPmPWz1WwUM8Q3Hf7Zyi1CSwgBt0QupKWlmJ7VO850e
frc3BewFwjhc+W1K3jpT02Jp219u130n3BeLg15vnAPI1zciQVE07a8qF5SApNjJ
qpHULh0ij+w6gCSZqz0pME5j+wWmbVv0uxYftJ2KsTd7vgwfnsxt+hd6ZwnYyZr0
WzKo0cuKEg5nAhNaDjmuzbd/ATnnpLcsqcX5JovQtx2c1ZEhBPDHKtU64rMR/0JS
dGL1pTBXzkcdX11cQknNJSGMjLGfBG4hX0oE8x641V1CnSP+abdbGWMS9ZSORB9m
ETOVD7Gat0hN9jjVcEOAvxhOtT/JZcJocAUxBbeuxh5sjM2DLPAQxGoabkhmmMIQ
zg+F56wZeDGqShviS/EJj+dp09E3i9FnjdguX9P0tCv+iZ/M/djDBOmkbWpdbmEY
66xt4j4kLWXomHgiXpKQZ2WWkYYYRfW6CNBwIKU6vTNH5VmEp0iRLgIobxF4u9u3
CnFTPkHuGNSR7HTaLX3nIbR1BE3fgvPVXQAVtb9+zsX2srAzIFJ7AKseCL7liTRo
0Z7ANdeYSpPX+zQBc6aUvn4e9GS8RdmRTlLQKc1JCia8M0SeeKoi59jcggGDjObS
F1FwDXjIHqUx+9/+z+TApKE5zVgB8r+9N6+lDwravVlqTERBiZ9exRzasnH3yjqc
+TrMLOwBBnAsyw81b1a2Kvxy+6opOxklJh0jU9AdnYO8vzAHrNeissOpPsfskUyK
ZTR0EyYzC077K2jMTSLYnzbg38fIggHrgJ4f+W6wRSRSM77ja4a4i+8mGBwDjTjW
Lp99T+19cr6wG/bI1ACQLIP7Jhg8GyNP1ucHE1ZsP7Kch6Qs5Gwe9xWTZoieYtU9
A0pGXvlZ5DW/6Uac5naamfX2z2oKkLNs52nAqqMGS0XSUZzWo1kjd+eHuvh/AE5e
FFZfR6L2a3wP6shI39deabFTGyfE15uooFvbcke+D5wy69/LICqj1bYuMmr8HnmR
4J0+2PaSylUhTiFgpCF0+Fvjn5DpImNVYi3F0bddx60ZJQuash2KdwibugkVdrak
pDSQ60CxhoZ/dGxmOhu9bK4ayC5KAVWg2lgOE6EOdiGHvyXyUDXEMKTF4N10hkdq
BuqZLQNpbvsGrGhuLCtFcajFDAT0h1S6Z//ldN+aBUaVnpcjV2EczWleEQpCW10P
fy3MQGm2XyNaSBtFAdeAXVGqiyULcZdOEd8+GxwzqZ+arsfsxsaXadfvz1ShgCHX
xseiDhcSqneF9J1Z3m49rYR+AAALgVWyLyVQ3nPZu/NWIAob6vHiB290VCANMd3P
8PyUdAVhNJR+BiSG96EYZUaCC6XcOc+kVejOdkbirajZv9eVvLRc9qxhm7q5IkVY
a/80jRF5p05JBnyZ7fZFkyU1Q1eZBOm+mzYUnMGnN1a9QItwsxDp2lc6Q6Tsoyl2
26fiXMcYjOJpg+5y7cvqU1AwXgMzm8jCEElJQEb+MZh07pQZKZDD2+oiDIHi25aM
IW9v9aaSil7Tx/uhm17bS1PCkWsah+QvhhGy3lsYWqGcBnlOwu8XNPS8P/7iTpth
2w732C9/ID/Q7smUruWIctxulDWXMVdQsiGwefJFk8R3sFCA8Fs6kG1vY/lHBENU
Y3ZwawBSSpFZQBlyoNEs7hUploLPVJD8xr5HLqlraMWboLzz/6qiWvbgyvU+0EVz
lMDmM5vEwkpFs4nk/sVhJ5fBjpQITMTBVaC2/lhm92tay4SrNZdGvNSz9FphVzBd
YxqMTlrm45sPU8o9p92uPFS616a4XtUgfwe0FRcjxMqk9WkBgBWTiQo2NbDqWu8r
dAEQZ+N7knCBAOmnDSwfe3GdTi4qaIB2RKCOUPBlTTuqo/JbxQ1t30yMBP77bmTD
7XT7EayXP6qFTkdJ4f4O+iDSWCbLGOyPrqPfNEfVEVZPExrlgzRaP89mLAta6e/o
Dkwanr9qd9jbrm8G7x/Ga3uwKNrjqANK6sGF7IQg8A5WaTo7dEkC8NYRaFq2lvuN
FwSkA0MfLUM9WOReo2rkHHvNZd413anRMaNosyaSpDfplhKoT3oxCg5uszAUhZ/C
WE+ELY7AlKk8V3gsodRGQmX77XfjTKPKi89yyVjdZlykjXJTOsPdvPqJzNMWrrHF
Zj8VZQrSepACEHccGzifcJeK2GgzKVy6fe7kaKelhtt3FSfC5h51jJh3lbUGtz+u
E1r6ZcKX7v7pc60RYm6ULZay0XhZMxEyQRcX0FLVMyRbfdXTEwRCjLkGGKpJmWbM
d2+rXCLxz12jFL3RFHWYpEeajkcIsPuL/YKrCAAjnYOiJc0D7CLzJ7yVOJkdP3hf
eMHxiYPQChIqAUuRyCDq0PIP8lMYOgUr1unxNnBBY9PoJHv+xHgQ2nkcZhGONHwJ
Sv019doWqiGWqfmhZ1HUrG1CBnJ6DIC0u142aoAaWSgBrtZHRUZmlVGLXwULZZuV
ZMFZIVWD2aFXrJZHBdv5zmm6gKlGIqe9yJ8+9lM8kHqFy2o2K1QIexUMBxaPJQXO
7LIPEnxyPKDQkSQ1wDb14/+jrANZHfWBgdjvDR17QhpH8wWK4bC2JVpYgLEQg1uV
MLUvn07uZj3mMxp15WW8YLcQt8jDSz1/yVG4FAvQ8YDMqtf9XlrA9fyaeHQ84/TK
5ePMoF0iwuvIoj/Qm09FmTHw4CsDx7n5i5ef0gKOgBcvk4+HuxanSwOFJRcLAXY7
dvhZjZWSUrder1dZbFnvaQMrLUlfZXUjw0P1xmAC2cxZjFt7Ln2wsCNZi3GYqbnM
nDHYFV/4bZLJRIfwf23Y4UbczV6WGp37lr/55LFRN/KPDdno8NMdLLcoB15Z2Z8U
5SCT32QOO6WtTNT+vMSbxwxRdCpwl8asa2J98JsQ2kiJQZ2du6A90xJ2RukiWTZB
qvfDTMPNyqFyc7CgxsOTCacf2qtaAOOU9fbBgaxX0WiPsfgo+pAdzt/R48RzNmWG
b4Vo8q9TUfrNfcgLhPlvdN+czSNRM+yZT1jte5cUSAIMZV1iVx4ZV35/TvvlQ10k
n+1SapkgiMYz0P+O/zEeTqr4LC4RTUW846eOC36XW2FGrr805K9OXAJzEGXznsg1
kaiqAmovkJ5EwuD6wEL8lLfKRVIRXM5M3qOiUFEJ2gBfMRt+ttXEqlSTbCMEDPLk
Ef/AqdY+RrqZM+PlTRT3Sjm4IzKXPXddEXk72GRhylEYElq1H95SvlOT92j7HTE7
HxHkUIQmH737hOgagd5je5YKcMeYwTCohbexMZxUSH+7A/V3FUhEX5TTlnFgKRPP
tY6QeOFEbIxUz+uv92JCFk/zd4BJNbu9Sg8X95SqZFM0CKphIc/6hV29GjW9/Xg4
fEaFmV6BO//HAjmWc9EKdLwwm5TkPYnmaHHLDAjgb55XUHoiULO9/tbNvIH5BgTM
aBKbTNDdkL1Bk7ab9d+CKDVohnKenSGb2CSMYYtBKrq/WOMc1aGfHe29nBu/wNnf
aBymq4u76CRGfO5FLB/DyXGtP/f/u85hE9nrQUe1+4GJytYrFgzZgFKyUoNMKnm8
uhTHwTs5/mYtydnYxRwK/WhPscF0Lltn6ZYEcptevQORCg4xxUDmSZjFzOWvIM0C
fkhOBgLq1+KoN6vvqAJrmhGQG/sp0rXGqCzLDDoP++Y0yrF5tMBk0RtIt6UX8BSR
bkSUfTm/YvoMmdDP0+0MubI/nQHCxfYjqa79RlMc1Zi4xH4Z6l4nkUK++q3HGNXX
GqQkndx7G6Mbi6e80u8uBvYv546KtqvSl93hw+A0wRwXTtFQiXK/33kc58NZDqdd
eR8G/24iLTNcwUSg40VU5LFakKgVZxYkNJhG34cKBvFezCEiIfXg3pkS8U+1txQw
OdXCZDwqZ9FDt0BgKb5MvJbVpL6v1ZI27m0FIkMcg/4r+WrXGnhWOk2tWj8Lnobs
5LHWrorCqwxhExSz1xQhsXqTHfpJnleLsp4uQgpafWFz6XuZA/kdnC+BYWQILL0F
+hQRhnkGJz3qdkAPh1lrA0gB7nECjBMJbPRXDf0xykhxbMddMOSKbp1Svsgboo1O
0ikIiyXvsCoezkgkEfaf6hiPMD77cDJITiSTt2KcP4c46CBnMM9YjByYWFrh+flV
qqT658760XAjfHi0fmRMScF1E093Nhyi5RgZLfAYmaptgTSA4W8cJvb3uUuIccyX
Fdwl9+3cpSccjTK8voNux/ZR/KAWQnln3g027fnypNIr+LVaXdG1WqUcaPUIyVOv
XeaHw85hj9E//njVaLZqAnafnBQsVIR706LMEwWNaCckZHGOEyM/gb/KlqLFHf6+
SrQQBxJDAv7L50kJ9BZAj8YI98uUYP6Lfn2GBstOg5Cq6X83R2nCPHH8OQFTCb+G
O7x0mThhc9UaSStBjWlN3gXX/nefnQUqKpV8Lq5prbN6muFYXcA09BvsE+pWpqZf
FcwyBsOBagpK8HBwMd16g/GbtNKIuB4b8yfg/KS3QQT9JzJusWefI7nOnEi4Fyy4
bpZZgGCfbWaap1C0Hk5lAQ65c6jAAKa1RuRhICmFMTjZxzM+KFgOWO6DiWmS5rwX
vjjNsgWulfoVoz6I7lj/BW4DDrq0ID5GCUSGGS7aMeu0/kxple3upbn9Qf/yOjvH
ek2kkewulkSdDNhGA5MunaNTMfKgAPHQ/7mlIbYPZ+JPP0GbYeTuQeRMpQQeCj+h
ncyR4biddjdOHOcRpmE3kwldKvwPC847AqKyvgliVubKabloVNkJqpFZuRJnP/gg
d3LOHw+nn+lBjWE5h+2zFwCYnjYem/ICG+PtshWkDLcGvUOzjqQvPJ21Twp81kAu
QMdQRK25k/RvU6CVeXQBQJ47IbVLYnkYmdponiGbRYjo7XcosIPWDNaa0SBrpDfl
SqPw22gTtCTHzSBcVbAgfW1IwUNNV2D2Oy0N0p0fBcV9OgO30R1Y3o6yaVlNNXtN
CPPMGR51iQxB18OMZ9vBR/aMtotCNTYVfBLyD726FxlzpyA77dMZmFiKfTe48eSp
Hpk7dyaDkAuWOjIl91o6laRKehFB+SXfdd0H59/dJH0HGksY19a908BtBJ4JbZT4
ai14KvUbZ/yh6o/w7TEMXKhlFwxxD+8cJDsUPNVwsoBz5tZ4jj9eMSfn+RIJNbzY
Go6+vOLI+/4iwS0u2MOx2hT4UCs6HY+jLYYS87ANKfno7AO4M/XX8D/4s00TV1fO
XrDttoA3WVxv3kvQTX79QFjcxRIqqaLo6Mr/Qq2u70wJjh4MN34HHB3rSyXycXOt
BqOdm0XnWtTVkVsAkNSE8exuLQt8e+eP0AOX8m2e+7krgGxVUf0jufmAwJS1xWKM
E+SHIdpSTDsluhwdcc6K6OyaBUcm2kCDV4rIcp1S+gf1Ph2r9ZM6vZ8KNRahpRUu
7Kqez3fiAzz9mhJ+iIlr843b6QLbmqkk5knEFoMnRVXQ5WtR2JXXIql2WXbRRtCN
clRpaBAZTjj+TGiA5OqbcJTnHXyTXfc0J60WrzAWPAtO+S2Ml0IGL+wjfQMGYD1Z
2e8ZgpFnOGP8R4uJp+DFztVlH+V3fsQDwh1mcyni604jQ11jFEgPCg4TZcrQaVur
MTCXPzlQNgM3aOqNRGbFlJVU0FqM4RiEBnvm4DMzYlF/C3/MKJCf9htwJjLM+yAq
LrEc43T4zQ9J7etoPGz3MEIHaEsseRowAU5wOmSinfK+l53llAYtsNYKKgkSRYko
5aOR96m95o/V4WSHBZRSlLFqu19nJiRZmdz6d+n3fjLqj68Cqj/+7zy4q/GyekzL
nxsAqiiW7r4CL2ZXk0tmmlWtND7w6BXfGq/GS8obsdEz24Yj3K7GJPeWwvx/ChmQ
VaT5BSiJYFL690cMBEMBWYBwRzlOVIJwn8jmg6j/ID7c7uo8JKkN4T+TIzwYOq/g
wT8ubQ//rLYUreeatCKWqdMFbORwqq3GlT16RrBBd08SWqFmmp1KSpaxtn3YY7nS
KJSAP21Aq5WMB2nb9BXevv6PCEw8Nh9S2GeIo1r9ALlpie+/jFeK6BsKaNvux6Lx
0MESSQMYZsjX1q0nSsPrqvM1IZp7O5yfKT1stPwAejKFYm2N02vtvZIF56rLazaA
x/LC4k6dzWNyAuIhkJYa9ctjYimRNaZcejQT3MVVASi+78oeSFGQmNQJwpVSndnz
G51xmQCIL7557AH5U4SAXwFmk51GsF2GXfo+Vy34bAV1+pCWmw6SP/I0AhLyPDNk
cfJHZjG++WOWtxm3LCkbU1wOcXhDxqBQA2+UScTDi0e/uelJfm6iU/eb6wr4khr9
iBDbJXWuWFlQSNibtbD9NPyGuVQx59BZ38ruZY43bWh+A2jKm39QPKXOOChjzAqR
e1qyICEVIRBZakyUVoRew5EjBbuBDIdZNWfva/aImKb3kAumkHs+LVLnNWwZQ/H9
eRY/BI6ZbsnMQpkVbX1QT4gOqJIBjslXiwqCLgwqVMNbItRyrgHJ4NASalMQOfmX
0KXgNcRvYGx5R98IlDOAX1hHFFaDdMSlMr1HtWtyp5e3c9oCM9ZIbgh/tNZjiiu5
G6ECsPq4GYu035gt1y7z+i+Ip6eb12066PVdAjWewS4N1QJ8CGT4tcu1YNTK6or9
z5uJg7nFBjxG/vH8ZYfzVp3q3T4+c/W0oqxlnYD3PKjMRAYAiclEMolbvsMZ7Z2W
fH4Z8znzz0h40TBIpVvZ1mTialcc3SWVpzUMFUFz8spGMkGEBayc9WMuhHoIvm5u
ZZWErWO66TwthX8b5rc96r92Ut7HU95TOJ9wuHf4SvRBVpG0wy/DMeYLfqc/nbbx
Reh8n7S6pWZSjPWHQVz1Iag2xGP3jZ/uWG2wTL6D5rtXDu5sfDqt4Vs1mOhyoCE1
UDIGcfGekxYBj0hPgr1Z4xd7H7NzcNM1YwZBel3gf/YqQM111DWteNdttS+L2sY4
EdqZ7qt4K5rBgk6sTJ72heDUv4XzDvm83CV6dbRrmHx2Av0szLEdQlKOfjeu5dZi
CVO0a6QRemYrKHlBWnT5EaNOi5mCENTHLVPpWSMXuym8YvtMwkL/GtqTX0plDfnZ
bDRXgSbjzR6+4X7+3B4lxUyv+YO5tHjPWpDCDD81oCNmpDuYX+EpSJTuRxScWCb/
2ZfQ2CFgsb5+LaxwT0yOZFFB7bWog8l4fPPjGp6iCa6mlPba5MUUkXBg31DqQ5l7
w/vbnKrvDRN+p40lOgOkV2m+cCoBCYjfjPgNq8qFw4qG/7v5+2ZFPY1JiUUV4lmF
vR3EdhOnco7NvrEl0vZwXB5sYbsdmhszwV+7IJ7y+82AyB1ilIZpq2UvJgoA5Qqn
eC1wOLzGYVaHrSeZxz4ICgIRFIM6Q6gzocNMxV74SWWzw/Jz1COWR8O/b1Pno7iq
9BdEVG1pJ17nIDhlK/PUvmtSIOZb9eOBB2/zziMnYeRvrX4+mOtOehvGSVAzVw/d
l6d0+hvE3/aLBzInHRaeJwCIooc+ff3CEYUDYSBfbKSCkZYDPQzuCnPR7VJ7pfyi
PhHsrmYvF8qCtcaQr/Ys5pXsTp/1MHj8KE5eCqGPDFmIlwXTSdIAB5leJKhlLBbm
fIfUKePLbMYfMOLiU46rHVpIcmSrHKZA6o685SJmmuhrFpRePN8YN/6zAJkYGetY
lroV1A3N+vpRyUz9L/H4tkmiBbLzHpeIcO18y8NTQX2TrRwBTYLk0gHcj92PcyJ7
ZnsiBPV/pXL7n+2zF9zEL0lf9hqpzVPcb+cK64j2QjXnNmNWx6gcWCWCcHhU/dYn
cb/2AsJgJjTaF0C2VFuBG2LRvEvnBiWJa3glh30U7LEuVkxALZrk+nwPbqhPgwBW
AmpudKD5P/2snghIO3340IxaytRQbWOHfrGewkHQzkYsWsf4pm7h4V5PSSUNfxQ7
XuhwvbjvMv/HgB9KY/vuEbShvcat9w5OnE1RAstrLKa1Cc+Z9d4VC4PMG5PeNOho
8mr7jl8VeyaPaocnWdJn0IwLAyXttTEuOCDEsqhDmUQd0wYOOML51EkKRbJacwcs
Yf7iAjShOQDsu565gz9VZmElsNI4sp8992qg/2KGEyqyxcJC/HeQfBLJ9+uUr8hR
+Q5Ti0vA57PS2wia2a58P9KVPpE6e51d/5sJKWRPh4sDpNcXEuhxxXGsONWtMTG4
+fMVG/P37lY3CjqevIpWxsWjjxxaxuLqkFpEMUtUWN2XGNacUCcw2G41mftagNZw
vxsmtrrOKrLjvTmRmR2hDnxB9nvYcjO23fq6oA6+2Xtpl6Ylf/6Ld1l3ywrTqVtc
twP7wxq0RNV0A9Yi+l+bi/QErd2NSjIZZf8SyKrwUuWVt/xRzfNdDaDYeOLGJnAP
3BPj3Sx+hxXAHkbtqM53pIkJ6J0HckHCXDaxXULC2fObdiVV9v4rgrgCWsGu9Njy
KEVlR24yRsN2vDFlbcGZE35x86TPsAiDd4KB3V1jHHKj49v+up2PlAFhXID/xvbp
g3g1/XGi3xuXVVCOsVOg0gUKydGIKqJBye1qWdxH30AVf8sj90SnAoWxqTnH/cxx
zjKIdJsK+Cw6vk6x2WW5/YnFy2PLDflK2heLZn/aYomVjNGgKC74igzOHPC59Mzy
hhs6vkC+3K7zJC7eNuLBnutzFFbINed1r40PNjCJoV+Sfxu7xi25MSOAlPZKV2KP
uIVehiNYHHdPmxlrAGdMHNj3Ak6QJDK1iIhC5w5f/JwmuGF9mKN6KccYXkJx+Y6g
+m0HkLGea4TBB9FdymKfadK6A8B6LJcKaUYmY1UaMZbLvUW84AUZFMJts6a258gZ
/BDrqmsGnzYSueJJy5LCZNQIjKc+I6Q+G0HP+5AjuUuXc9PHmhGEGcS7f9efHCt6
aXmyhSHKotF19Lqte1ch9RsuuG4SMpTd3Q7T/0P2nYiPm0SVLcW21PRZYDQEifiI
qIyuaGZHJdD8mrXZ51Jn1wCNs61HreSmiLiOLbYJqlL4ny1ioOCcNxhuSmrcLqsn
2qmJ1UY/bxIdFqnM92rlwe49/1kt7/Ejs/3JEYvRxhX42lGafrxbm9+1bVWgyeNN
BZ6e58/QOHqaRy6RVZeN5gyIveVZvyTmxo++WsaBsGYFIUrNjU5Ppx0vSuEzqrDA
Gjt7V2faQfd2BQRY4awvgDCWeav1TkZikE8OPb66XizzlDCj+Ml76j5iunmRgCd4
NddKmCaHFQJ0uCpMVgnzNtqcQBQ4OIEMBEKtK8flwXSYCAMzI4holxVc1/Mt+nRu
7nwU0pjib77eEPhOyOi5HZTUirHRdAZb72keAFAT+tEHzD4YafxAVygAITMf/oHC
u1+quL1QK38HtKugd72N5b+60EgRpCSEFfkA7utbrLmrZJN07QxRLXDQOh2jq6Yy
iaIGpahmEjKM8l20hlg+J5W7qNUPi3zEfvMKKjq+2XkC/89WUUH52cIz4PyWa5DF
u+CntHM0ywb64GfvNy80AUQ1EpkXXot6ZYWZ0WskyJquGA5UEjlXrPc+6KfcjXsG
Oz5IB82XxvVbuWsx8op5H2o0k9ZHWd2z6e1pZJ4x4S7ovKUuIfVkpM5UIDSle+l/
RcG1wco95jHYVFrzMz4jCztItTZZkppOGRZaz0Cw4oQbfHCBzBvPPNirfeFAW2IR
c0mvMM/DuB5C2j/6RHstfmhvO4U3FWfnV6d66Qql/axRjgf9c716vs4kVG34Gpox
oO/JwjFlt93E8l7si5hp3xl+5olAwZQrvlTcZQZ2JT+EiiErC1Z1NErtBBcNsaEL
k8cb5S4m7SXLBd7Fg0B558zHX8/125gQt6Fk9C6xaLUOxfJeKNmJ/vjmCQFdRSTz
FML4FaSWVyrpoQm4DS1QcwB6I0+LA/pWKgyXHJ/cBWyG3jyLFNaprFAVjlNoGSrL
38VhRsA310WRm35AZVu9ONVY9r489vALyYUY8y9Mz4nDSSlDSDLMZqiXqrYPiupq
Bw8Qph/HwgRdSbNBBZ7rgvbB07bwjazCmGbY5oKmbRxTh3DoWM+aYikSLYMdeoHp
KN+YRoYhy635jh8F54uXHFh2ZSQ+EEScfBuP6FrlLaicnWRmf2D2dVe/fzhUNAbM
hCXJS9oTuWUOEexvjSReYPY6pGDdTK/hgUqdsg0KUrS0rLjTb+F/M5tletzxEjGB
b4+ihvmK4b689oc5AZr+PA98vsTQJlGUKSVn56ByTOUNA5olimGUuP1HSjy7dbAj
6cW/v6Y6WoEOqVaKC03NGPjSKZTwKuap2FVREXJFaXTRenWfApo+ZfzXbxRR0apo
ztW8VwQR75ixKYwytR/JDV9XPw2St3J5H1y2UX6MM1Z+rkpIz+oF1zx62j6UOFz/
oXV0z7baIAvv/S1LSdbMZceXv58h27aHo3LFMFO9iLAZYizoqe7Qzv1kRLDJ2Vse
4xsctA3E/T6tRScD+IZxlTtGc7/umObMZrJJ+5tQGKinrXzY8wABnlwsOPv2HWWz
eEZAuPZ1zphk7xsjmw4EtbZ4sg0eoYIzj94dcI6j03056+kMvdRIU4NcUr2+wbcW
ZeCdHEnn3m6dSSnvYf6lNxQXOBmcZJMKDCBDYZmo1KmYzIxqe7AbYVkvaG4+ZPc/
CfwQagV1aWUYH1ruBiTjVfr+eekVDTGd+c33vpHwKFlJSwSu/5vKR81/OV491BZ6
vRYyzoWgxSEamZTUIfj+5oQLB2oRT4nDf99AcrxKdM71F/L1DL96F9/Ivio9H26S
Re0E/WA0ICl3XTbyIuQMQwOmGHUGislNfbyRpM+H9+2KmD2EVdHA/qCejWkr62QM
JfkKXKpdzSXivQC4Hef/yGvVWCdxWK8uN7MieybNA8xLeqxHa/pTXJW1d+5H3qzb
UI/xNn/XRvUhAOfRdcY7L0PbNRgYuKkdCUSjQxEL/ncN1AfpBc4KWMAcy7HmrcVh
p/ONhLoZdpF8lMcMFG6y1JO/ad5ydUhxbka1NiWXJ0QT0MNgM9UfoY4SA4ZsG9vP
z3YxWHIyHnaF4E3gKhPRm6KKpFVQqHviN8uoOjkt3BG4az4hP1x2nQt4nkTUyomk
/wr/7zxQuedTT0H8rZknQFzzjsEGrE/mfdOvpcsdh6jsWhnotw2TfMPxh/pKxT6z
zfwbKK8lcUIV7mSciYK5mbX0VT1U0Zeevbyyqog+4kFXzunDS2ActGvVgwWKbQnK
ivGZRcJwsesWjN+C1wqmjDyToZxNKy8jSFFkWReW0KNj457yPhYEQUKxqCcOhqf+
lycl/YeZRk3MI9WGSzG3DKt4BaUj0wtJN06OE6hs6/BlmNrPZmCvIzuAZcv1uwph
Dkm7EOvC0u9hkG3hAOA5WiVzpNPkq/PT/+Gd/30ORZasTtB7M9/FHczUU+PiZCHc
sYf0f+q9/03HLUdxNFOhyuP19fb4G8/R4PTalFiHhZwHSgL7z6he9CN5Ok6J1bPv
UwKowpj0Wmjsm6ZIS3YwJeguEHL1e4K+oP8Y8EppV2ZKP0RheIU06bs3hu1IHU1U
Ef2qH5OVZxSnJt5tIze7eYBd5bfm1GJ9RPnyVuvmZaXtcOxVVlbEzRndg1sZXKIn
7zTiw0WoaLKL6hH5s8k/vPVUFw1hpo3CkoBig6K2orfw5h62/73werf6WGwd0aYc
irEo6PFSn2qxBzLgkIaVrAY8lMq0n7cb2NvREKcwdbe7pi7KuhoycYfakTRpJ8WC
4sGF78s5M/G3CtuSLoa1jw+lzfjCAY527dF8sM8RrDdpVoOPgSuWnI4ECJTPEpv4
Ggwg7NCJAwU+GVs2YIRu1K8eC2m0T0fyzNqgX4KGYqfX6/hPGjI3EZ98X/C8fTMS
IGeqf3JuXSg4pZe7lxHNHw0/fKDCpGMvPFHwzQizwmzv9ebPwXpQtyDxaNDO9CC/
sxYvX+7vomznHvaIUIp/AZXwaNyzcWHuYEJAKzorfSAPetBdK6kH0nqPDvuJsz3c
XlRfRKVLeXbUTd+OWvC1j2xUu6d3cSh8n2BVQzlkRdvh+DGySfO1hXAb8p+Jl0PZ
DGkltL+36i60Cz0tHB9B/J4MBRyNG0em7loqiAuumphRyr8OINWuW13xPQ66mosN
Q2OTspR5RrHAEJZav6Vd5Ie0u3+awTwhIA/s17+ucWE212DIvrha6xgFdU917kqC
z/la3tlbKHffHTzFlS3Vvg0drWIR4aS5ujNyQibqdAtTDHgHNM6SNf/n3iPqOw/o
aOF47QY35+gw5/kBHNAVdHajr0HiPPANJTVkpn+we3SFDmrw/DmmXJ2+3s3jeF8l
/A4dea5ILpI5O7quVSGwuKq7q4zRWAQvnZXJxmJ1WzS/GcZKQvqnTBRIDeV+j9xm
pV94NiVmFDqIELNfwDLMu245RYTglF6dLI11/i/daXol59MuQe2H+4ONhN4vc+TG
3qlbas7buQpppDKjP+rmYL1RXujlcN8op0tmt6QnqMaXmgsRHSv0YgelAZbUASgA
BholxRWLCAyMDJv5xZCtl4y8XQIQafAAi1CKniaq6e8cMyBEgpejZRTzfrgUN/3h
7U5xkiMJ8SKjF/xgiFesd+4U66ZqV2RoIfU3Gc1Go/1IgFbCFPrk3s+PUK4J33Tw
Qvu/KLVKflZEzc3EcntirY7cQbQ9DXWkEO0GVQKNclgcoEl7QRW/Fz0SZOgfT6Sh
NZwy4PRf8k2ZgEKLLWr3eicHk6ZT+cnfHxCaEdrjgYdD/wwm5JOcYWFZUaM+UdWF
JPndkyz1CTFMuPStyGnYkUmxUhmWkZoslzdes6BNWngk2/l3hn58ved/jZhrL76L
Bb+DxJCbRlbGyfEQ3yzj6tbCwLf1VqfvkKPwIowPSd2PtHxmiiebY3d8y9O/rGCg
MJPnQVgqxjR/WW1xWw9uR67oMIXkeJVbu3BoqDdzr6pK4F4SdgLyDf7hfcKfkd3w
sLFyBMT34hLgqbGrAXIAE3KPJrJAMtfBJW56DGOlvyO2zWXbKha7bWp6oDJx4kP+
31hwqJnBJSI9UXS7mwiCciBdM0ROBfkv20lr6oygNZePXCVOzxiJbQSnRgBVDSSu
USUGocDHMLC/nO598fARR5h7U397s3w+PbLmBNh2r2CoAbmuyuP8Ek8xOYP+WY6P
8NcuGD9qNrieQKTXqMKNJtzN3sYvJs6owfKI79Y0vqWer2F1t+PeiacTI66Cygth
oioPmIRu34r8PRf4sZTgyUg3N5Nxz2bYrchrSqU+yRWa76obmUTYBv+vvTj7WVki
tXOjXHiwCXgOQAXjyi+kugZZlQ6hrxEGhjXD7CAxULQFctKW5rYenOUteqInf38Q
1tMyJVziKuA/iFZYQ+PjSwjtEjLnmTxwk0reIyQVPavlA+AZUve43ogGVv7tVkgU
v8+NEAZitSGWof4UD0s9uu91rYocwu/V+MOhCGixCQBp/P75S47Q0TGgI7OT625s
8tOvCrDf9Dls2q7aneCifeqT+V/1RFgbALUNssHXjT8TG6l+tgyP77/FveeujYLe
1zno3kwG+MfunCmHVl5UBhO8x/+I1lTTMdKhDF0BIst41M5B7XP1UgRytDiHBMrT
DP9E48EMmLyc3iKTrbw/QLkrv9Q/8VREREOObEoSQiA7H9fbvSVX4OlVd/DgaTOG
s7CLUu1GbNcrw4fTSDi1zHJIoyrxZNVas75TY0N5IGgpLWYtXWu7UzYTEFBpVANq
MSxaMr26mo2VdkatDqrNcs9Z/Tl/A43NyQo2BkSwjiVBKTdI1v3XRGrvtT3+nTzU
`protect END_PROTECTED
