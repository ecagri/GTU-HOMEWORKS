`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wrLlGmpWFLpu+GMVlJL+Z1hZeaDey1bI+LxMQcg2VJRP+akyiwtDGKalIHov9nKW
tCiFuGHcD2hgTvFDGwPPB3Sqfn9Cuc4Pd+sgDOqJ6ApV+CXtnGu6ZTKoIyvDFF/e
X46a3Gppryu5HsvImBckYPJ+ne6RQ2xQHBjuibHXle1KJOSF6Q3G4YDmdZwcj2N2
Ohz1lJuLgv9FiGqJb40z+x3yONIaUhkOqVsmYksAyn7wBtv7fVfKSx+V3lKP036s
udw1xafVQ8wo5j5EJMJaFnaYPBiU8WyzmhkGbQeCPx/AKLh+23rlhD+Bfu+odYaT
LW2qrrVg/oplH6dAGmTkH2AtbTNJKDDHeiqSmxzNyzWYSkgdlMDRWmghInBtD4N/
8uhIU2vDO604qCvbyMytKK/P1RrmU2i3nclYGI9zokNZDl44t7XD9p8xHu3aTgcW
ONjfUi4bnzOgo+6sFBBaLLhg8ewYjyRlL6MlKIuZI7Uj+pFWVcwpRjanfzVzgtgc
KItX0KcPLHqTkSVFzupeAPVm4zMPBCiH857Uw+z3e9qXyiRIFg3XB62qoSLJ8jA8
ibts5h634EgQhQ16ukh6+k6ze9imPk1T8JXcpFVJkndgsd53Ul8avOyL0sIDkGvQ
C8XQej5zuUpNUoI07BV7SUi3ci2QevEFEZYsVuK8RX0lITOEQOxwW9jLAk8OXXe1
P626yjceTFVU+O2PZ3cSe8IyT8tBQYxOq7mbFqnFAffNmd9EYTbcqSUSuMVetfNp
/MhrTGIlNTwqGTldnt6LP4w+QCtT60QoG4ex/8qlwG6E6czVNVfobfpiQgSOH1OU
4CZyvXqPtFsmBXQLuUqXRoRyj8N7SkDgj06zqt5dcJQnUxgOlsrjIlN7N8oIhX2U
rhQ1qyZ9maz91ACLTs0YTbgdoFvvOl3VoKLlySfrEeirsgasLtNnNRDQ+4fk6m5f
FoQVQaVhYNkuIg8jm+DexrtLLv58OFMKv4rQi4DhUYfxsSJkY0Qh9C8ubYjxzdA/
6n8qEm4qMAOm0lU0JJpsh3vVZW7J2HHpxlNoHyDd9bXu6sOidLPa0GDWGRdOJFsG
z03z2yIBrGdbb7H7e37XTOaMXxzlNpTeuyddnveJ44KNTLIVr+VQNC9VKOUj+eIC
c6DjghqbLCjeJtccFeHqxEx57TJwcvfg+SnSKMhLVuCxx1gAF/asJN79++oN7o9L
h3Z0Xk1Se4LUo0xteoDAmKdTXUaCuivJUBj0LUg4Hrg=
`protect END_PROTECTED
