`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y87NtapMbRnBA6FJzLuJMgUIlTi9NWTI4bvCIhuKnBWzugrpZWAaRgmzDG/SAPo9
T0GLhCjgpfG1XHINo5760Q92So5xtWVdorg5yMYYoddoggZOm0fcWDeYp3R/JuzZ
ZETXlsPf8k2fkKA1JtLluSRKLX1TjonQZqoYV5VBpgx5T7voPeva2f7rSMWAg0sN
TIypOS0YhCZB9rBuYXOaXy9iXV/qwGMQB6avp+pHLMEVjj26NfnuOGp4VQiM+zbn
LJY1VnRUKBoexCa+UHDGyTPj7RxvD4G3nDhc9Lf+/GHqQuQ3h72xtWZ/8ibboUpj
MsFPkn/bLk1B3kGlPDZR1i2Z0u42xDc+zBT45JHk+g6so5Nm7L2LftcAbSA/cARs
MPvjFauxvFcva6ZuNJMJE+Udzo47IQqiHbhWEr3+2oAWr2SZCp1tLNhX6FAkgTRI
auRn13lrISrIbTNy7PF7t1gtmGm8SH7mZHama0IQO1nYaSmtlmeBwEfbmPYCrTtF
Np0kS+CYsMg8DN3Ys0CYtPnQRz0GM0GEFA6j5GPrTETWv2DbuoWU7S3RUN8HAuHQ
YN0qXCmcPgCTaFSViDYd4kSuP7wbI5vyp7cxXEWAShpaQVI3+uIRjm+0ayEYvNr2
W4j+Ss884GskJK9T0nnKhLJj33n4oXMx2h16TfZJz949ZhvAlwFQ9y1vtSz+A5Vv
yMhopBnjsSmHzWd2hxZoqS2B9iQNVDOPws6sFdAPG/LUxNwUzY+eI2WwVedtXXRh
AjIpxAOlT5zalsHXe9zDG/juX5pDN4qZVTmFzWQd1I5CqWbOZP0LZB9bCcQ3IBmY
YYKhE76vPt/pSnwdqzSIRE1cJcKop7Lp2/7E3AvCCuK/SI01LWg0u45sWg4BCroA
dyLkPpmwn55qp92kWLUjdixdxmJYzpmzks02mPrtGKOJmShUSXxABXdMgkrNLRvb
lVWIpd/+FdIXudd0vNfTfXW8ChzEqxNMFnlBELKlYMkoUpwX/Yu/IrZGfET7zakZ
5PThgAHWrVpt3mAjfZ2LS722FedmxbdTj5wR+VI780LfxXJIQIWA1u3Bb88B2H+/
bANO7HheFvSxrXRzhaMmobprWGwunxB72oXxImt9JgEybbpDcRUlEDln+vEC1vky
UWIl6u5AD7/E8kdOr1szkIzksgiSlhNa89Aza0YpmSTTyBmCV/cs7jCOHXwLJ0bJ
`protect END_PROTECTED
