`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a28YXZ5FZfwb5ZLZM1SfL2maPC3kYN/OsVX/TV329R7hiNCjhJLAbujNbIzJBmBh
8yieNoW9yFdMS7oQTqmvY8UPAdpmBBESlk8SLF81FGAYSC+uONT2HTaVLSUb8hPS
4RZxmvJGJFPeYW3WLc724wrvaLz7mKgRoksHZYstZiRAlwVXQa1E2CiHg5sjlxtj
Qzw7FuOZcFFL8WAVt3ypxBAKguI30JcKqjBFjiyhHBqaJ4DZUhkQvg1GaFZtPT+h
JdrMICv8mJ/0iQ67NA+WtshcX7+aRYw9ymymKz1ttDSdr4SEUEiUoLou4bGrvuRk
KE6/IlT1Q+cXIXBnGAcBbOSq+oSr9T4APCA7F2hgfml0F5GSuxR5XZinc7vlGYxw
LxwzX5s7YPReOEIRviFXtSO5IBOqivKPvUruN/+zNIUCsPkdQ97LFxbPqhfqnC4U
hb5zNwMeQF38KmkQQS9qFYT2TJRlW6QWhgmyIlsf3b4CO2TaZ6LB0B6+cIgXNVjQ
eAwvT9ob/qBplzg7z6MXWLF/m7JZkB9se6zVeOIMLtd3VOjcHSBhAxO42fC1txZp
OWx57Fz6XpBMdu6bkExRIzDikBNzMUo4Ve99DnNczrZqY/xWNkbW7m5dorGSFhpk
XQaAtk6t+fO7hGEj9W5gLdEghi2oz3l/uOV9XdIJkzY5ZAikbmkLEVSInVKiMPPs
4DvRSunXoqwfZdV+WUqd4FQeRlEoC3WM9kGLAoi/ttPobq0kg12oz6q3nYYK4tu9
XuNI47AI/P3NuVRsjkMMdRXlBOmhAC8Ps1n9G2+OfkH5n+qIGdNi8ytwgU2H72Sz
tFAqbHruDdNp02k1UZ/nNbj/ReCaYW8lrHBj/yiBRpYx6PxPi10YNu2PqaNbZBbP
eNlMIs2Qa2MjqPhY8m63ZhdAA/JI8+qxxaZYn26xDtu1JrPNRLZ8ZEAzWuXeuCfp
rOFaTHnbSZZEIi5a9h5sAebfDRJBD3AYpKfqdz9fzZ3WUhXb+ypvzVonvxX1aNcG
DpfXKhfmTQKYS3HJlADwo5fszNYM9TK6U4Ej23GmzU8vJsuxRDpp1I5V2w9cMU23
MrMm8evk0/m7nI1Ymqk1TEsn5iuW/1j7tU9nF7unOYmtPAPbxH3zPHc9Q00DAj3z
eP0/8lda7G1SbZZRFCOg0SFqJ/l106ldnI50KKxTrYZ3n7+h3y5ahzmRk340bySu
v2bOftCZmxx7aeuULPSP5AdgOUuDPaSTBAlMTVCj+h8hwpBOisJd5Vf7sCavDiMU
atW35agiccAWoprkVJ94VNmlMcFxUQKsCbjkoSpO+zugW8zTAUjuYUXsbcwouq8c
zT6UftkibtetqRVokiLr9tB/0/GTfWAedZBt4o7fvOxLvztRhtS1LvZA30GY8JGP
uof4Pru+bdLmkWzfZeR1UCB9IRqCVAZy0VaJKmUvbvg=
`protect END_PROTECTED
