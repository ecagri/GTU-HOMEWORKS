`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KbA3PxrGIZXxtjUJ1ggRmaV3QcsuQcL9/gQICMlUAXO10O95LzzbTbCMRQxLWvzD
uj7/tRQ4yy2Xee1uD6AlrBfcD9wC8tUogrKW0SHLltBahjnH/s/HUu4qK8S50NtR
Av8of0RVXh+n7GKYLF53l1E2+TXjNGfllrdjJlMYdAL6YRpNF17S3qhIE/v4qFSV
REy2HgeUQhBNjfBiKidx+YsFZBfS+vGcF7EYDI//yoYJmT6tvvCplR2hN7zfg6GB
SkSYTHhdGIVbXVdZvAMH2qrR1FmIx85YIbTPw+s/wQeY8Ur67Cs1nV/qIeOwKsWV
RRO4FayDL9zLrj7aR9RupFBvbkFBpKn12E2rowjEYJ8DIVsUfRci/oclXup8JwfE
MLrMkx5Uz3xnAAlFNqi6x3lX05CvNRxIF2ek72OO8owcedWTgCOr6JWoA9MadMnC
VAXU0ZfEeBHPMNsFmL7NQ3ALGqE+y7hCD6SUcHbCAlYLAx5wgdgNBJm9HSbA8nzb
hUauGD7GVPaTLCfH3iFaByWQ8vd6l+keidg8re5kAGPo4F6w74/gDRVcinEdiG3N
PkCkOaPbconpbcUlR5dgMKti9m0CrAIFlqBsYrCEr29aOvhRTvvrGZVJyUZFgJUh
L+o3AeJwZHX3zw/6V3Ge6/xRlMKWFjSA2k4s/KfYsrW9Z5sHl+EWYG1o9rbwendv
E9fOls0DXxBvjp4bUevEACOPnj1gJoqY9aFfj1knxPtmehmdBCq0nAK/aLJ/XtyQ
J2+ZoRL8MOmtLIWnf7tuRLe7yxIB0hAHOmiH0/anNKzUCiPWxE+vkMRmFOs8fqh2
P0OntVB21fXM+UZE12fUKHOcplqVRnCTmjiVwHtx09W/tc0tMNMDSz8bS8Hg7rk2
1gd4IQxRfMwl/uHqEI9YAmsHT6kA4jt/H10igF6T/fe9YD1E/YnTS/ds9SUOTCu4
OzAFt+WsEzi/S6sYi2E5Q0npHlJPdSdVfHfphbHRkKmD+grQRqw9cqgM0+ZjJCuC
WwoqWgdpoY2DZaVoTmnx6piZ9edgrbHPiK4NmKNx4+JnX5IljNB0yG8QbH5681IX
9ZeryKuJh+4dz1vxfdLW2z4u5MuxPUA/R8bi9qbk7va+BHpdGar/DcoiSzT7ZvzW
rQMOzxxpTtWbNseeqbuk7UGQwxBDVgJm7PvsmL8VSy+IOXKdPGBLTutYTYwB/F/Q
SVPjyqyf2vNc2fIe8IgzNcVUpc8cxAZIRs1cQDIJs96UU5OQHUj+PwmaYJC/YRQ+
Is8A9VmhcmIXw6MU+jvZkvPTzKjqCB4vvqRBjktsBTQzH6QFxdXctWarWTt6pbP9
E8rKPfllBrY/ahrOW4inuHM3gpxvGv8NgRFMQgKCBfd9gq13I8eCv5nawSKIbg8o
uWJwI+QGFPFyLHAHE5l1mEDK+kWK1a1v6nncmpONFlc45o6PxFAOSd73yt4fqQDG
yETxMWP62kq8uRcSABgRqVFwTmMd0xeVW9T/Gao2AiZW9F1pl2NvgKerhHGDwvdT
P4OWyWdKoBXNPbkVapCc5WEf6uqb2SEpzlhlMXXwAY+wDZxeTspnuSTWbfF39z+R
M83AKbXNKd938kzgHf/6GzSTnwGeKSzkR06RGbZh8z5JYy3d7EFMU0d5c2HGX7mW
dz6aZBf4KOyLe/JZ/uHTMf2+bgQscOBYULQRr96HRXgYdXmdSi5eX/kVD2QXIAUs
7E+vzCx+S896lNIWDURAtAqospIAJn9zOwQ4wayOKbsTHDRZodV34NNnUSrNSXh0
csgHQ/yDSmc0ZzNmGHFw0TYPcVSbogBJsiO6TPRwNIHu/MHao8jNOYoyY0f+ncrM
sAeeeXW8U+kqoFPxcYSJ/EioN3iRSzJVZk1Yb0LvMsplqlFeNyiUGzN0tAw7t9FN
sN8IpKPvRW4Z9xEV3Yu/H9ZhHbN/rJkntASuruNEga5nDaCQRdXPBsXih4+Ubecd
Hnb73oTpsT7W+YDLkomfoWLn/RCd3Ud0cV9oxiDpufKV7LpHW4ZTLBee4lXuEhYi
us2EPTVYe+q/dj5/HlkMY/GAEQxtvEdp6Xc7Og/704GLhLYD5AMbtx00XGM5soq3
BB9LVHYJi+02OzqA/XQaxaziHN9vKITi4lfaC2pCVtIKe2XAThSWM9g7IohL1hUz
ZrEYNlXA0jRee+O47/HpdlL6uvg1EjunghOqvCXyNsSPmABc2ADWJ9B1eHUFyKH/
a/cn6B9sB1N1Xk5Up5EkpIf9CCNO0D4XIfowWbQz2680wIysAC33ntJeehP9Fv9X
Yc8/hyk5DMkj+m2Hl8PzqlMvK0rlq+NpnTalI+dz4vr3RKtXBhnfIN62EJNNOc3v
ul8RlRQTtzaI2aWYEkeBE7VR9JlTCAMwhk1VuA7zqfzzLVsOTl4sqWWEcdQV0ELU
5gfJjrM8GOH7ATDEJv/EhdFoXJP+ItzFJv7nPw6+MYfyFBrIAOaM0iANa8fJJ1r/
8vzA6ox/D7RQk1D3yUFn42yHq0GmWTHbC/5JnRXDbm+bKEIxcSxWshgQAK/NPbJ7
hyjMdssQa2Lfqr7DCUBUyijYhyAk/AJjAiCUcHvR1D56tjAQbq0Z4xrTK7htEjS5
U3K+5qfqXBWqxzi+nHhX2oZHF1hCU/b2We9QilDpwof0lEjeCihptVcm7uJDmGQY
vikEsYRxRbd6TQ3+BnuUtyTE6wJuo7etYfQY5emic/pyuTfbHXyJXplsiHRsUDoz
BSqaVqzfHRfH7O92N+0LUkfljvATwvSoY9Hrm0wPHTiwyXseh5A9KGF00CLLEDha
0/GxvfVUGtM1c+Bvd/QREj9p3k7igMFExos3ieKtOKngYB7L2zpkubcHM+7MpIMF
4kWRKSRmN/j37pQvsGjbe2BW0IJtRKJmYiaV+py3x9oXvxpvNKj1wX0N1ez2xNwu
ELM8sCRdvgkJOVEqSygsVwEBGTUDLGe2G6WkvURaWj3SqK1IrHcJKd0T3Hktx2cQ
PWnULllLvCPQEdTRAgtSWndRJKwp7kefd/qGDOkiyVciTx8KA/j2NFqZdETwtDn7
e9qsFQTviY7pmTyzD4roi0HbytXtKBqRosC2gm0b2wwqMOD3vCYI3YpjgjpIBzoM
LxO8i93FCA6C8AvonBMZxjuSMy8MugqahYcQ7hPV/EJTXth6rbX5zdpNLDHgLt0X
55NS6nkfVz99y/Q8Q+7JJg==
`protect END_PROTECTED
