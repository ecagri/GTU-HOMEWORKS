`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oPChZVy8skuYmFOeVIAAgihk2QZ4D+UIpOgkfHG+zYPmYl0XEx+sKWbLrhVeqd1W
7b7Xx0OdgJEWp5Ir2lFxvjJWD3uivJhCN8CoQ/dbSIgBQ9ZI2uaTO5/E2heGIm2V
mZJc88jhUThgnDl8tS3YsVfBfR0wwZyF3RyMkdfzUoUZPVC5LTRDchdzMgWhALyi
dQloDJQVpb5EBzGPnF6I7Srjf2feijXwrpFJnBj7Z+/etrKsa8rq4CipzklHa9T1
iH/Ovnb4tXjNSUNdXNTp68YR/mYthPQ8VznAH9zKoPf83XJfVLEeyf5igVOw9Gt4
caJqyYajuzbD/41/59VKgVLr3wTjOjtTpgYGH5uGaI9prGvDCoUH5eObqzRtvygw
Y+pcCJNC5iLL02PTTLGo7QF1+FRVIHIXKWcguppoLgma580tNfuYB56W8iWY1zVj
2V5TkNtepsvBDohfaevIKPHl34dP+sfpTiyRv0Zr6zNfwEEgloD7vZND7MWB5IV0
erDRz3XnCwFDF7jDHxlwKDAmm+1kE+XQiJRVvzsbaSokkSAbVg/jaudVMdEfcDGW
7bhzAUrXnbQbq1qkm+mnTcYrk9OLc9BDVXseOXE3dW82XaZz94aUDmErEqAQesgk
/AcmKRXqA2WLPinZTVLGAIs38YGBKrqJ640cdCwF4djruBaTX+D+2XcrRpLTaj6L
hxwK6BEBUxH3HbDEwFFLs7d+fwzMshB3axIfbgBdvdWxZ5CZ/M817pdZZ8HKvnMw
rqZkGvrh7Tr+FJ5m6h35qpNKNc0Iphi5IJ7XyvFVfEGdQYnQKmKPHMvUs/ZOd62S
UDbnmVMaJvoLFWUgRUBszTi+u4VlLTObV5NtVJd7NLFPTVgQn9e7v/z5h71nl6R5
rWoxjj6cIMkSIi3odxzCwGHUuIfobC7zXWz7a06P2uV5N3dFmYxVoa7qononL+kD
lkC2uxfXM21H/dprpMm0yH0Ote6SnDcT1eU6Y6oAZxNOUxDcsKmP6b5w7osICEej
ZF36s3J6todWugPWxaaDWbyFGuIw5oKAVCV93mXRWO4TqGJU6k7DZ72WkCOoYn70
S8D1qquhLJPsPubTClalUnakprwhvYHCUDK4s2hVOs1DHWVV5EQpchcKVQs+yADw
aTSrRvJa3ahv6ABYWldaszWm8F1O+dT4Z/2xCvvpJO+v6UKhPwFAq0eVaj3n6AaC
vF2lz4mVaoYuCImpPpGSTJmboAX37yfEa38TbXO+ZaLnHlIExOweIDnshf0SpInG
faiB3YZndmVgaqfOzdtjMHuHo/L5FQjdWv0fbp/fbBvQkbtCK6dyJyL+gPnLJRrd
IEjrCQsCj3RIRzdIeKH+NUvlbzmmMspqcC4QMZboQ5MyGZa9JZhK+QVQeLcRiFcn
wlh/Aj4OQmxf5w285+YNozdxXsTXkA7g5qxkLeeorbTckmYup+B0MsW8UYtTD4By
aPPYA01l0bvPvhFqgHBbyKY2UPM2DvhbyvYJAt08CfBOk4bP963/Tv+oesLeihAa
MY/6zBBzW1/+E+NwtZ+LcCOsmsM2bZN0SXXT7RZNw5p6ZJLzTgKl6kz1DOzaJPah
MVSbo0Hr0BgFFn66EybXyqRD+pkitQkh3MXMCQ4ZEeVZUGcgS6bq01O7DvqgnaVP
78eu9YJRJnqzW8otV9SwxBxRWicIbYIQultm9Av2d9V5C4/zRQgKVWVeEGTQJ35U
fAefnR+8x7FTlLdVDQVxcdx0+sTsSJDE1odiBWaprFsEFCr03dq7FgG4wxTcRr79
S71Hywsexd3/90xleNFCmK8ybk1vCSikBrYAzc1fcKncekp3YsgjTvKLmhcBVdH6
A1FJmJyPaFCwyLWzLi/u9XAHwbpYV97D8tbNJrFW+RPoGmW9UeshI8ACRfQiizp5
7BvqaJx70iCPkwnsWHXNFApAfaLjBLPV392DFSPJyxMboSTMkeW9GQVP5PunNyjD
HvbwBlohrvp1TuWOx9jMZk7tuaNgvjQnFGTQZWHWEeY3IXgs/9bk96MPyDieVh0G
EWjLU9q7CeYra8vf5jvRQ1P634TaXrV9AHdH94nNFpV5vojXh5i9pGazEyju9Qk5
Y7lg/tvsCskbitnGtmDAewZpbpW4APe0UFxRxGfESER/k6TxnEP1AaynWYCvG5Dz
kfKNvBjpX+eWVUbEQgwMgrUc4QIEU8gDdvUSfjyJVY2pWHbJ678jYdlSlpv7xaeH
NGmulCPDSTFZYnl5z4JYOHyabQJwLg67hTANrQSSb559Z5DCcywSnCNrmPaSrU8S
EpTc7qF4G2e3I8FOCDiq/PfGjFLz/49RheDV0UbuTT1M3g0/DbiAKfoeB5FQ16rR
VdYS7SOonIKRajrKEaQA7PZXJEjRJIilF9QArpNzWMPEx+DqoPY0EjDk3I3eDe0E
ScZ16bwzvq8lurjYZUzK00WcBmZQGeeiNhWVD7mSOPgk3ONCppkAwBWalJyDNOuc
K7kPoviAkx3OLSLGS0twx5hrqXFxrNimT48vZanMoYgnHlTEsHQgCmrg/PjJ3sLC
`protect END_PROTECTED
