`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sua5JM84SLHwNhiWhorqwubjX5KObT7IRfCOtGW9J7PQc0Rpnks2BsWhhUekF6R2
smaT+83r97nUfkgObDd6bO/tIALHQeq/PUGn8rpzC9qKdlI4WrdIuONTQOwm5Qle
x5LL7nNhajADu9sHfrgEIiGNiUuFskMLBGrRZPyuc0+KpvT+uv7S6biPjPerroVr
9UUFCBKI/2Ogkq2ZK0m0usbPCzJWXcldGVGufIeqxBUb77ERkgGlEWm9jq5zBAaz
XAEWmvUpTQQ2kJImRc/2TG7dn2lGcWJBF5u7ilBx06VlAVGKhHOqWPrqtyYQEODf
+NcZeFM/qEr86S+VSIXMEnKapeAUGkuUwO3unOKKzVX6AV7THEuQ7Paz90g9EK5t
sXiz4XpEaWA8a6niwhs+h7Jymc2bMCYgv7FzLJE9shc9Z+euuWWUHngtWrE1g811
398klljKhSsu6HPws8yl9ciR10wtzXV579npvOVbJHcXZKkBwcrsmFuF6iDc4n7S
O6rK8osEAY31IrKbsjigdAXFSixcMcpHcQEQtGyq2s3WHqkmQNXxLyi+aybioWYI
SYIzYuViKwaONCuZ1LWr5FoPojUQj5cxC/M/FAkR4/Un1Um8HnGEIKVnjXkhOZFC
pGrrYgrXaeQwBAm4PIFr/k7GmGmxOSZWnMfvclRh3gLNeAGJPTnaV8K+zQo9AusT
OzCEghCvGk59zfvr430tMJBD7k3ljT/WiZpmxBN2yrjac5uhQIFaiJ/c/nZk5358
dz6YUeguhFesMlv9avUXgMzXIR50Bp8jWhptS1poBY3Pxl7KJ34N2aS84oNQ+A66
Y10aReAeg2zjn26t7derJIU/K3J+shJjHndeY0N7ppw5zT1OWp4pSrVw2g5R4bIf
ljY/c+b55jCBJYK06w+JcrHkzgg40ZcNekj8T+IjFw9N2DfkDdECyEDeqkzAAW2Q
tTmfv6GfwC67U3cTsMIjjPWQi05CW0MkYJh7RxwWXVInhkhs0D0IJqr9uAgt+GzE
1t9Rpl7BZHM2BShgO8pIXC0MlgXotYWqdQMx07LllEnSHJYqzxikODekLoTSkUvN
1XXIrqUSwaBTWv45KaFkwOAUwpjZCA4txi4/9MY6uOqrpm6aU59e3E8hucqeZhvc
IHttW1jxH40/u1/tswIq4pLorrFOJzJt57MYU9tXM30FXca5xlMuj/1HpUkMF4KH
vknmTm9qUp/zbY1RBYoKh5nJIiHVhYu7p9jX1pkuXp9coN/WWJ9X7TNqzJndFdIu
+Ox75A5HHLfLdLGtKSaNBM7g0lmMmLaQ16kxdS6LS45aaMAtgX/4oUstA6IqRNkD
295L/D2bxSLppf+7Z1kiUezpRuEctzNiZSRPyKgt2g6csdiPT466aMcjs/Cu3Ofn
Qkgq6B7CvxSEDe5yqjxuC5bh3sIO7Ys6u+gTYKSjQe8N4uKVH/qykk2NaLUsrZFP
i6Y/LQxdlUyS7SpY0Rq2lMNVGlJPttA3UYWiux31lplFZFriXuoPQaoSJdbOfP8L
FKtQwLtcaRskSyOgjiZkcD7m9JGZu9mIJuJN9aiao2/PRd68fSSv/3vtabrYfenu
dBPlUZXChEs1UXAGRbJ4CgerA9u1dQPzqrOqTteN9243VgJttCrkSb7xHqch3+g/
I44xDxXN9/8mIv1RdWFw9LAQi5eq+UeID4+YAJ0pWhp2O4FonkLXOoEJorLu+Z7+
TwI0+zRWw/PPVLhTkYSmmNUe+m87oSlHFAiXh/JFvI/aiswy2DVybKUiSzMFFDvV
BijxnVrSw0GQnF5epxvbmp//jBIn0wp9akzAo1kyMobP/c93lUst1Q7vy3iwN/qy
LCewOoQnRZELxuWjczln5FYL8UShKupFSh3EvKj8tft5IxvSuroXc3Ay0sW22TXi
CXsR5Ei4gZmQsclNfGj+TSJWrYi2MEXn8bwtojotVwV9XbPajT9V9ZtRB84VxOgk
qtS/tQx4EGT+/+NEwfvRWzitLZ0VHnwdo7iHydeEAsqF7IYwKxdpKB7zs72zMzDs
f1a4PBjo19K+FMlV9AeueHd5i1CjOe+JRLLvK00MsxZ1WXkFllYKvM5iMbmB4w7D
Pq4+5rKuN0bjfOsItpTFtZRkBBK+Vtp2vrgQMe5qkxTaJhe/I7AYOwxCpcR0EVe+
+txShqiqy4z+rskjThWSG4flQPtX4GAaO8OPF11Eu4yeYz7kmUEXtdqoyWPio+82
9B6D7ZD25m68aAU5arYhz8hrbCboI9gcO3/3KShHiO0=
`protect END_PROTECTED
