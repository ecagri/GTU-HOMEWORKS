`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zok7/aahryBouLVWW3GPH088PMFhE1EYsNNKqEFcS0dYkVn4ERP69oZX9j6pgsnO
ixxEOkSii4Jcg8hRnL5PVlijG6i5zJAg8bH2OhRVtB2cc4BjP9Ze53HdiNz2VY6J
SyYdbTyV8uCiPcXaRmAM9qA/120CCE78OBEFlJlNRIRi2N7zisJrQThil2cagcse
IgKSFcR4ZcquoPOX1AyvEMw/BRWhsphbL4fEmyagknF1X42kNYFe0CHklI5t2OY3
SFwlFENOHnj7jtQ2cZxLEEtvPxARHDuifdp/EkfY9w2GAnnvBSfCCIt6XuIcs994
6sQ+Fh1bpKPXtIW5Qwm43DiiAFklK2C2HZgmzoXPj83CAWXezS1838kO6CvVw3Qc
s+ubXWlUKvhXlSXInzDa+7fN4h/ZQabpEoQUaqqQmbRdKhYJ+y2Lzsvvm1IN6Y/j
4a3Va8vQSRERUUCARQb9CL2eRAf3n1bzWP0Bd4rGXTCuCzvqhJNm+3WM+dwsK0K1
nLM9bqSmlLw4Lb9lNGmxHMN/Sz3cQsELKV9/5tG5Hpg7KNoeMq+8+4otdVwDsQYK
d75MegPVsumChQlHu9uJEth6aqQB3POlD/5erLrFaFYeAoWo67gYDC4N8PWajuFG
0GlrFJu7FE6M7qde219hQiB34j4lfJNbI/aMiTfikR3D/CpHiENev8lAq7T2FZbX
f+Mh8N8kD+pdhPBGX2wGvezlNrD1frCVVVslHw58L9CYyF4jH//AHaIM5aeHpzoU
wo3vIJGn+nkRgvhy6Q3ztGYIPdJxozmLYaGtIkgs9QwS97ePYGPQj5KBHJJuuM8E
LJo++x61i+N9ig9MoAaPtZN8BUq3st1quKxUTXZpZpL/8WMLI1oZjnweatkw+Kzp
P8ahrOoaSG1zwiEHmB88vB+jzclLkhto0KlFI+z1nHM50krSvdQuuV4/bOkGfF7R
QUbCh47QLKmEOWnU+NTq39l/dOrrSuRQ8jL0YmoZaVOwerBHikWsViuz5SUmoAJR
xaUYDlKEeren0XNCewdXHMtSduvvDHdDLuCGszhbNSfhZadSD9YdCzO0l6FSTYP+
g1UUgWqcCZ45VCFiXCU8MUXCS0NCOxz/YtEheHVpea/bYgvgVNgMzcTaA7fN6UWi
EIIRUKdLz2nsGjnUFwi7v7/GzTcOrpNSfV4cG0SQ+d8bLolLd1S2iRv1t67hf/YG
aQ/KDyEkYY0uPIHYForZNIaE06/bzBIj2jqAUPRqIjur54msuM8UlVDGKpkV9fnv
KYmRGYknRyt/OU9xGieyy1LW/tSEfyzy0WxEjz/v6cBOJiVhagOINYPCRe4cI8dS
8pyXGhaXcjKRn7UHbIHlLkfDR9Kyy4bsHBppbqSsVhOsOB9CRtN3iY0pJHs0zcmc
QEr0nmpC3Er95hTebqete11pyD7VOufwVe1lKeXKbRp1qu+Ny2c95aHIZv7mqCPO
xT9ZTS8CKY7FjcdZo85WntYKOhLwfqfhbBdsbwqFogBjD6Wos2J6o80VWlnoG9lW
tqBmOa5xaB3CwizQnuX6IpNFnGTqpWDQIs+LHvPZ6MFAYy06Svn5qV9cThZhVXyG
jw2FOgv9AjEF5vj7faG1AFUFyWDiIkdf9LPWADVnCRhi8u1Zpv9SSxQB1gcDCDlL
UL8SwCv3vI99nr/E8ElfnJ10abHNZ3BFS5eI/qmbqnIqQ6IDoriJ++O7pLJYSrtc
sJehYeii+4jaRavbE+FRKjClXNNlXePs2wMv2QTInxpl11xU8Y5GrSVcg4xZxCE8
+zGOKf/dDNDX0q66lgSHpoweFOXsSPlbYPvYfo1wG7e+2zI9qXFWRh3hRnclg5Ey
hIjV4HL/5H9Vi838jqSJgNw6KlYPbvPFuWNcVzU4ev5Dpnjhe9K7Jq8wjMIl3vzQ
BpiUE+m3SJjZ+AXJmLPhrT3njiKrUMI6SRemE4Hn/zI3kRMpMgInAUbIgGbHLeUX
KoDGe2VreHiUKrGtPs5zd6wIs5VzL9BbCniCnWH6dEnR0s5XRFU+z3b7c9xiz8tX
DSBKtdLPCA+szo6svcSJgGGOeuUUhcUBdIDpd2toY3Mx6fQGFkB/YeJW6T+Npvln
5jMRW1QuDlvH/xyI3LpFVF30FN3cavE+UYp8r32SwT0oXRoY4wXrUcvZE2jCkA9d
vaxpwKJYgJS3NgP3nKlKuMNb+qEd3Fz+lCClzW6qEywNPH+Uy7BdWm+L3pC9CvZf
xOQEwF2HeUEYI3+F8Sx+Z386rNJmfLbBYh/8sBDuG2T5VNuuLgpsnlBQOONoi6fG
UKydltWcjcR07JJLFTpkm4WH1LS86Z4HCZtAkosncj+NrmpvTeVKN56jIArqsfQ4
qoNhyhz8r3ULNq4CBIHPfZj4wMC168vIjatqloCO4fb0its1ULTgj/tac8dpgPK5
dT9Wb2CkpxAUxXgUStlH9U/8QTyCNYSVWXZHj/JZr26mXJGidekaEIElkyPFmBBp
jE8o44E5flQ9D2eqmlZ/vbG8rkXZdqoa6+YI34kf3OXfHjGNweQKNMkiTos/4dPQ
WNnxcXHlEOxoYb5bnHgHfAQoKsL8IpAiUnLvGuxQRuPTyotL8dY4Z3SMtOCYSsxy
GMB/8EaF65s1Y9PfdLQE4N491kAm5Gen1s3F+Qe8oaSHfWSglQP6fXBe7kk8fA2A
BLJoaqFugFxnCVFTsayDmE2k63V9BqDVGJ3kfw5gQbDwlu/1TG3rWJ0Vq5OTja+0
KAIp86svsQ8gEeV7/rZ5QTgpzWUvDtn1ytVTfpAArusr2uc2ER8j4QD3KELDkcIK
5puoazJffkFOyFJcEcADjNuXT2CMl/yOsRqRv2aMXEDS4RhUonzWeR3K0lsK7uU+
xvlNisXdPjP6F+0J2LZhItTSZWHzprqwQa9OEj2dQs5G7E10QjEUw3i21DB0E4Od
Gc9JY8lLDpbf2MQcGUrp5LewxTiTDMs6Vxmit75pLDqdPq4NCZw/isSjtCFtLrq7
EQ25Iji+NM4aFdvadbZStSiQ+Ou+hW3ZtAf7odujpBeK1Kn3Zbv/bwh4p0JFhfvD
KksHQYFGI52jXTuDVurRPKXrdMniZxjVK6l+gCe/YfhNqC3bMkw3o/aV2WqKs05K
71YKdPlUjkEUFIrCLjlU4UeQDkKvp7F0v4Lb0XuBKot86bFm8IBZN4LjOL3x7cFp
zwym24Qzjt8AtP59Ctrzazfx17Xd3AoFlDfEuh1Vi6nGlhdJoghaeDnN4rXNUujI
Qmyqg97vy9oalayvB84mmaWElk1Bil/WNtkz1j6VQ2gkMQZAzaV3seyVMGi9E7qP
PHiClJ6WV/HuxdXLIJ8XnsbNH9jgR/ZgHLkN0gn4CDNDd1SCc4JuM9VzVQN7ezwp
NoF/gY4JyEpCz3tYxdHPGS5nfBcjSaDiJVt/DCtvDOLX1Xcmjjx5h3+geikzqRBO
7bb3LVYOvCf3vTNtOVPK6uOrVbjCe633AtEJf8ZtBQysaVkL5HLq+Hp5NoeSrFHx
3JdGU2WdATiL0Rkccsimpz8fEIZ4KjVcpvFFwSfDRak6Pm8tDJVEtIsLmKcPbTqp
v8a9u7j9DNgAe/22YKSphBwxRraPVQL3bc7MHEpywsttu5Tb3sUPO1+xQiYMhN8M
9OYtMCuEWemIa5OBkUWlXnR6El+3bPuCsptLam6H77Pmnccc5NAMIGp0aUL5sJeD
aZtYLsX/DJvovROJ6AVQeoF9N+tSd18U7BaKbS34OTLcQ7IYyYKpMH2UJQOk3tBT
Cj2znDAP06c6e2dzw7Zc2vF1yz4O2ceA+Jk7u1J9zEPJqjuR/eu5TrUM9ExYypt5
RIooF/qexa05S/zCYmXAUYiTODYGM6SSeZY2g77CmBbHLkuzErLwbBql5LVY3qvB
U3JVqKZ9ERLiMOaGfh3SoNuibN7Uz5BqeASxDRvpctQSZqcXo78xeyUVUzbv9DPL
kUF29vYqjQKr7MhRtdagKz5GBG/LkbviLEgvcizl38dFZLAl0NIcKtrTuhoDoEKZ
bgryjwU+cUisGXBQBHs32nstfJEpbf8LIIrAwvUk1aixbU+XgxXzv5bGhqT6F1R1
WZwWqhCVo3nz5kPODZyMcxS18aGRlwnQ9OjDh0ZV0eOIY+ZsgXT04RpBvZT1wQwx
LSQaysrSVttdoCmT9ri62KpsAb88x/QW8kk0b7d5M5JQlmd+RaoNLye/7ADDq89D
APgKOAyfDgE7CXHFp1pcpyeDKEM9ohhwmHVogLP7GycFE0YjaWwTm1AwkjEzHpmC
GIX3tnEON3cmcE7PUa14rU51uTO6wVElbNfDPkJydC/+5lnRvmyTnR2UcRYjpsmZ
kg15OoBtjhEsavwL5oBjukcZP/5JhJpil7/yqmr0ZJNzSKg6xGnGRfIS6/CQhZil
DM7i/UZ9R1VX7k+UeQBl6AF9ksnWSufH+oKitGgFvt9+Rxe8SXpJmBDWBcnhVftc
KTWYMXW7XAC1cPU6E+luwMThFwqLbsHShDxDNlLeDHIaI1D1Xk6dOh27MHGNtsEK
W1Q5TtKWY3k0Fyjw6nlPN6NNVppw1P7uBsUNHSDtNa/rcleRKWADXXA+gGB53z89
/eqqi1RvjDcY98CIl7gZcTm2+s+SXiOfpLvJYN7tLxx+byfmpOU6aPdVoum+EK2X
ZrBQetXuXAUKTz6M0Sfn0bmmBPECJBDJ9sR5SIoB/AffmE2TxDoEh3OMn+75phie
safp+mdC05h3vtHvhlOnGtkopcLDraDa00xhGbk8TvWa8xMxql5pngWUMIIzY+u0
aAIzRZcHpWxlpwmVDIfSPlT04Iw3jfW6kga3GmFlPg6dpYsQ7gCK9J308GSImFbb
XhNWfUFjAs5TSXRqDpkvIWdpBDvZXUeInfQ3fuuoSySrrgDY2KLzo8trsdb9o96H
c/OP69KUm5JdIlPaJRzEG/ZNpFA25h7epESqOgJbD1BtRFxHjMURq9+JVAcp8aoH
rja3G90rXdbnRerEJ/hDl6iUV9qIjPUUrZ8t0BHXCF0g8tn7L3wQDDEK7gUgz+Qp
P834LfLlEUaVsijoqQY+VYc/GQu5wBGsVaVb/GT2Lfd7unhxFimkGZ5S7eYbSyfK
DeDuEcH2bG1uN9PkBa2gQwxJi2RoSXC8/C2zjjOiSSLgcfPlcnl8F7x5m6jcD2yQ
PCxolqtM76/52IEozyAc1+AafA1vpvzU40EigT1IT0Ykcfzozdf6QWx04eYYMkzU
pkGeiO5tLsyrZPB9HQ9kL1RAkWR+fFFGwfsBq3xXx1NDZfUhmieo4fFurXtY7Dzo
wGa+xXfDyieopYn5U2mPqzjjDaRBcnzZwmVGghotvygtwq1SEdkyevgpb31t1GK7
6Gd+qmxgq+AyjOSdUr08nW7CmI87ueEwZi8faMq8BffTnTPq4Xuic7Ko+Nat1npn
gQrZApP4pcr8aZ5/6uYcRRNGDrIzvMO4JGKGhympnQlsAiy/qaEs4XKw2L0N/mxu
7L/aYuEidtcbb2BCTP3yhtRbszrxO9T1DAxOdtotIdyAgvmlzJkqQnbj0HyTetpF
YtQWoTW38avq0nTjXXySTCE4I9DKZS7w9BD5li9PxbAQdxfXE7fIHVAymD95+JLn
VH/kud2sZTUz12apz1WVBfkBeOhscYMOZ3TBjyeFGHkczHhr9tuYmPOZDB4ZbyYH
Gp6V4TGHTaE6Jt4z8C8antNOMz1hrcMWoSfDbHtIRLKb234rRqP+0bqdtlJXuw8A
qs1EufTtc8CcCSoQ260aro+pTGc1thfPK51amgInaRgx0F6EcAsPAGXSB5t0P7d0
7ds1O4IWoPA/biICcUBOpjSYjoCpJDtOGy5O10t6CkNeEt2aVa3g6wdVEm32A7sU
pZGKZRwOVmw929llm+x6G+jItewzIC6bx7L6jfJIAvAPRWd7ocjJMiznx8s0t68h
tE/DaGgs5DonI0TTbBwf+45OiBcMSaRvt/xNhEGWL0/bydhbxNafOj1olMBbU/e8
MJgM4ibGzTPYYFUZWgazwYdAZ5dW2i4ZMfNQUYZZ7askByEHx6nCA//icN/McSk8
LRO9gb71QhGzurfFKvGpsy4R7SmeYr16/vNNpufXsoDqF7hEsYn4XdoezF/S2u0E
HrfuX6Th7wOfeEV6fd9qvw67arPHrUI+p6UIFPqniZc6fzqzMwOqI2RcKKUoF+W5
caz+waY9wn2oFKPRjA0fmP5MvETiY7oSC4+o2bsA3BFiUA7jOl20FBF7opWC/Muy
qSxFMeAoK7wR1AWzOwGv+TKbkaPcBEz9Z3Z+QKiTq4ZF/9ncNcLFAZoYVsyoHS8v
V11rMLI0/W1LNCbVuq7kNZfKwTWdJNjSMiZuwFeQkaKxcbBiBAOHG9WOtHDRF6KD
rPOydHMUEZ3Yp5BU4OU5mYAaJujdHObj2VNQEZ8Dg813kdut5u7fMt6vxJexr7/z
K1ysQxxxCH1z7gVu32zN1ExDJ14Qw2pmowN+f8b+rYUi+6yqWfiDiAXxmCJTmxj8
+9/vQ/j0F3MHJ+bFLTz3Dx6bb0E6yN684a9FeyoIPwQdCq3U3mVg/R2ZTOvEQVQf
aR6xWC07s9tDRUzUTTBLZxcFrVFwP7RrDoFqeqNRVfd0gyQ44EKj52WzhbAgT0Ak
JNJr/1QKLMufkFOTHh2FH+bm4vsOqAndE5cTbQHqiX9dsPO3sdGIUY+wDsjFOfVh
ern/MudvS1+b0Y1gWvDipMpQOZUe3RvvTMDnesE6kOXuK2Ha6H5JciHVIX2Zt+Dk
pwJ12gj2NwcYB3RNZvIuDlvzVffutVWAI/+Uczq8DmAVTbHiP+zEnWyxm8QXU9Wm
9u491xu/7FzbbF5V1LvhdxwLKpl9/ojSX6dWEuQDDaBJHFrj/AopgDJXLySd+X+u
mhB/fETx3aoShq6YgYAc7aJhQBiwrYGphW2fHTvagNB8a22CTqMXdZ95ZZWts81I
p1ym9UP3xbS8nfald0O5iui/7MMYcvYZO2j9kh059hisn33V2M5BsCLu8+fgz/mM
rz5CTWQMk2tJw4+QhtWIOL1VEQPhYUo12VqAsUYS6ev16QmaSJrYfOn6uFMt/V6c
uML4Lo5/p6dgqljdmBbSWqhENZHDM2S0REnRQptwCsVqhWXi+X+duxdKJCnfKh/w
vrg1rT//RG99XH3/Z/66Q8tttuNGljFwaPI+hp2TK+gjAkG7nxpRmWGEuUjQ4dVx
YWeJWul7Cp4nowvg+kyjltmclQ6P2TXi7Habw5COBZ2wLCGYTzCyRh+hY2vtuacy
kS5vwF7cSeWQVfxYxys7w3Bf4vn26O4bgAbgNX4Xl6lM4XOLEnuXVnXALiAND13e
WebqQGUgYQp9dRlDor9oa14t0hFoy54yazttFlEUcMjiz0S1sYngdXzbeDY1oPkA
Fh7yHCtID/zgV2OjEVg6vmbyo55rdUluoFKSB1oJuLuuNGZMR/YMDHVuR8pU/8WJ
FW7HPyAZtp/spV5G1gXAFFfZMtZ/TqXpc7Gqm07HZpkJWdSRzJ4vxTC9j+k6pd5F
lobmy+9ZHsvTSwRqVda6OTx0RJwMTQmE/ry4BKWPQZn/JgXwuTPDY77PRXv6sspw
+J3fhsCbGn72B1v+GVBFpHu6DRIEIvkmN/HIKK3AiyXHVlgsxnQbGXN4vfxnJM1C
FCtk/+LU9RXuI7vMHg31MU00jCtKY7We59gh3A5ERF936YByJvnA6C7ReBe7MArI
3LQhG5djKA2lK3FYMz1NdVP10xbhao0JDsqHUlJwofmrRbw+CY7cYGpR8BWu2kSq
Kp1rTVIWGS/rXWLojHO8TrvmH4NI9lLWgWECAdSmhIBVdfOeK/gSglvsXdv+g2Vo
IC6pJcE7hXiULU1kKPSj3LObA/ha0/Xprui+GdriZxh8HNyqHcepO/a+j8vg3dm4
tZ8YSVhsEUlMNvhsm9WKV3yP1WvBUCYYdmJsrRwdIKS8u6sDdj3HmKy2M5ftACd0
AZgoerVHsGfMbz+gwoeRDl9HF3oQf+XS08Xl/noG1SZnK7OW0ZE+eeJuWPGfcQo+
/wwwaJD2Ytx8JXAJJQyt9ONd9Qhoh2//m3OyJ5nuF/8Mt6cbqf3vYYifpOCkBhM1
egutFKHmJgtJ+Mqho/rMjZFy97OJX0WbuRyTvMjHXM3IG5I2VVBddekuwy3ZLQWw
o/F2LDhK31PkmgIroOx/awAKpaUS5E2g9QcQAtC/nMmuyLLaSirNcTyzWcFPXH3X
ymzkNh9eGMmxMMX1Wmk4VuB6Mzc/rwbEZziO11nlDb7+AmRnGo2FG2WBekLskfYP
Am4HsSlYsNQo6hJ2re0rWIFGnvcrLvaitoUu1AHSBaJ5laI8F5qENYfGur9W49HE
tFvU8zpi/imv92TASDlKvi6L64CGji22BG/A2FzXJNvNt7GjQCh96ZyWiQZkMVWP
VCRrge7imbNx/BkYitFwoWLL9g2Itgby58d6pUkas9MTauyVxlzOzKa5IrL0acOu
w7yALmkY6SKoCzCKejaPp9Sn38OovtejnOTWrYKQNQudCvFlE5a7oLGE2fAdmYjb
lHjJhbl1Yf24MqnHH/fPTXF8/kTiw+7AgG5uuGzoeyDM2kxBq6mFViXdPjRFxaIU
6cEO3UgQJ8WVoPfpLN0QwibGs8Kw7chGfQFm4JQnaiIGSKbsjT7a8ejC4ylz4X4e
Ql7c0sGgrFFWAT28gRBsfjY3Oe0OmZcQ3HbEeyPA3in9bD+Oo4yFuCpeu4yaY3ki
6PWwKV2L2cDxRqAiRtSf6SlVdrlh2pAUsGDr+CwegCkOIjcmb4/T/mWQTrqvzDaI
S4FED1R7ib6/YWhL7Y7SfTSQyynB8/s7kshgdJA2iMi6oyG534pZcLPYVAgtOGam
BDYeuGvr92BzrzPO/snCBNFlAhtwIlxOdfIo6VUQTx8b2qVjGtA5aeVxtKSS3w2f
UuEqNfVqCtMnUQ0vTQJqet0mxn4UtBt5/rNl/YxLVY/5Lm/Ma8vBFF36xJauQQTl
fTPq2qnKxXwnnLuh26vEtWNgJqG0XEIU65VW1Q3aI0WWfYkqIRKF0bB0hCLqL2En
rreULbDyjNK6oX8yaBAHhuGm+Pu/WHH/0XxvGIYS9tL9qIZMc2Kt7WEzkUeMdi6c
nM0ZEcEbzLTPzHV36PwRcnK9YrgglsdF+VUn+a8wIhh9Lx2pdIUs9WsSSx7vTkuD
AcpFEFtwQ7HEGEmxjp+FKOA6+Efl1XkDaYCK1TwpH0nUnzbFxkGRXrMj070CFn5i
t26ntZv7/pLiOFQexzYlXWSIvFeJa0ez7p+CrejwwnjAt12dEOrdj2tkD6+NgJQ5
46pxusHGKzMTpFW9auvD94xP+zibALQpaR+X8AhPvQheFmP5tW3O+qmUt6sYbj6w
oJcB3vh0pMQGQ81lQMJjFuRZHM9Hs+bbnJd1YEogZb+SxgpKyOk5+H+6/qRu82cJ
3rd7o/5ejc+k6VPXpKrK4iDc5lmMxMNu21JPkGzv6c4oIjp7QsTTJN+PKATnKvRs
SruCtgzr7Elsyq+CcDi5LVOx2voS4+gQDquaZoQSqBHmP8DP4QmsFsq6D6DuGiZj
aJAnHVPXltzk5VFlG4LoDUwSVDEewoxBZ3ocRsIFjMdlMAdOXFeigAQYZE0g1Ann
Xbo671Bbnn+fP9ohT375uYKM2rMgNAvwP30x1NWu+WsCrbe45ND9LJphKC6rUU2c
Tiji8HLL6CCbdSolATvwDlo+JjZlmfJP2lPYYuMEkrXE6axSG508O7zS/TwSxfZ5
e/OdLUZk3Qo07lvQb9UnHDbmriLdXjj8L5iAG+5Bgn8Jkm8nF9gUeBL3wSXqlTff
yhHdybhdzX4GH+LHmHwf8n8cI/zuHe4HA+2wj0wiQuDNUszZyi5iTGrY2uagA3hO
bm4cq60nC4Gb/PbVYSu1x//kL3hoz6NPuKlFWIOLp6UhIYV6RDTyJwDF+ijUAlu+
NtNa7ZbzvvQNNdfFasMeL+F+que0OgvaU+dHhKNk3ML8ZFLVv1lSAmoit0unX9KY
MncqAYB/sXQHjAA6+mfO1CUl10v1FnmM+yan/ASHlMdRz7rBU3fHdp+IkUEXvxRB
FWxrT7na9OCbID3ryEO2EIJP8kHkCPqUpub8Di3MW6N1wzkllA5fi6zM4Y0nkCIs
FSvkGkSTUXZ1NNc/fI4oCGWoipf+XDdSk/kF0bE0RprecWckt+9sPKxE1r3yIpNf
Jahdk0qTLkY6qcZ2eA2HDD6OewYg0pC0Mobw3q6qvkbIB371K4vT3/kWyjFwLLfP
JHVGvtH+X/oMcWdvnAr+y993CAlWqRWoMWHliRjN1ibivz24gubfxumn4+25SpaX
y6TGsY98hD6339JRLTvFm4ImVnGIjIdJxR9w3h++71gQPottjBxEluv4cUOvaDCv
xbHzPnf/jRLy+6c3wZ5di02iSFziv6tWJiXypSkd5VlDlV7ajAXt0zNsjZqDtYe2
yGe/20w1j/eML/VbXqkIL9flcKpatVUtFAoWnvH9T6HK09wfjKeoaLwAKwgWuOME
HyZqDGvxRXvuUFw1ZZEN6PEPYQbBCj4/svy3eBj1CVApW+9MJlneNQPnGaMlURkg
uk8Jaeu1Pa+7wkRfRnFDMOATIGszycXya60yC4K9xZq+slvDSMI0wIBeWPjvHPhQ
xb6k+ddRvTLmsmlpvplOiY7qNCdxITQV3qCgYRmDfA0G7ZcnGwIFB2TJDgYg3Dyk
NP5UWgaK6zRd+wOaZO9z+sRmhlvK5CYIgz1IQQlEK1fgMa21AFCtS1mWj4g+i1QD
mAY3tzUodlMIf91SKvqNfu9lygKTIqJJna2fdmkD1lB8roS3uRVeraTtnBU/Lr8U
SLOUDTzWeeZV9mumLpQLK7R8zAXjsZDkmQFE7HIh9rOCSUvb+tHjY3AZcmEcV4Op
2ZROOsD7CpJe0USp3R0R8//GXzUpWl0Jh8q9TbxM0qXW8pGblI2jAMfY8TmM5VJ3
plfxZRzhB00ohZIXv5+6SyeCh3yaDf9RRbh/dwFbAXnrP+1pBXXgL8/xVYSxKlS2
BtvX8Sfy4FkmPyG3q51aT1VRBc5YeX0xOT+OmyJD1UwMcxo4/cKZhHOftbDKqgCm
slSgmXBlDGW//r5N0RaVjwZRWHYx6HC9wbbZO+dULA8YHw1241HQK2qz3jY66o58
mzdXlXSsnodJTWB2L2jHaJVFdv8qutiaBrMfFSgWSDKGNOs2f92L4ouQYsARFCo0
GFtAJ5fBJR0pml9s+ShVYhzfHZLTxBpk2XMFtAsgWzK3JtvnEoGUDlTQ8t2kugYD
oCcm7ty/3ky1jXdBJWVqS1rNwt0aOmXgBcYM7yeSqMAdb8YwlKaCYNif9UEN1sO8
AYkxJq3bbJk66H/Qf7oGcDyXi+mxrDcGhDkcknYsRXLMqeRhjuj+c33nIE2sPwPM
mpDgD75sLBbveXI++kUBdz5zne2OKwD9JXDv12SwQdmAv95eVplsA6HSPSogZNsj
gUgxq+KsWGHGY35Ofl365QFz9j574xz/ezRyhybjRb+FAjerTym0jL1sT9DokqqV
SmkPgn4qme18dG9aNP4Yheu/nMgJWtRtQpXQPmGnN9o1Ow7Z6Drrrdg1UZ2MJ7kg
Lq4pp1ko1arXgxQMbuyF1IU2bSQqSP5m7+ZrfNcS5BpBDOiw2VyCUe+osgZNFa0d
JpdMZUngBYOreWu6ybcGM8se9Kb494GXUzEutGt8yb5/5azD7NWcrYo5CA3XdeSp
xiJWr+UAzseFBJ3FqHvXH7m1LxJvurlFiKtQ/oQyYLKFqtmuPnubNGFlrxIuMOS0
KhUKrNOcyWtN+Sip28udVRQ8zLFfjjDKZkhIFAEsQQfVvOZQpaxQC8LyjTeEswbF
LTxVH7yCDElBQxJGvz9CQH+NGNoAvr7FUthTnjXn2XSVHiRqa0r1VVTQzFZrfYZh
lS/OgPh000qr7Mk+a4SVzWkqBoO2uD/GRHYXssbbPx8fBOi1CzpEVi4hHAeECsHs
jS0Fkdwi4pIeBfXCqc9xyUqpXvDUb9iEqWi1aNkYxlWLK8FiTfHoLXqSBL6BHJyb
yspWtC8l9CqohYaTgKV5yV1vjuqVtyO85VkU+lmF1JNhe+iRb2NWDYUDCnAlUyuU
Oxv1QQr7yYR7RPTC3uS9Y6+L6HqDT0teegv86JuO59LxrkvI62q/gNbGgm3/NvjY
gi09bVjR79vgftCKYpPy5dmq9q6O/h594CxLDTW9aS8Q+Pth92g4zEbzFNoGllMh
OxhYg82BuUaDyV6nEiC/ySD8UnAdWgc37gD3MC4czl9ARRPbfqXNYzi71E6E3UG5
exAC4u0QPnYfduuQKN9BEcSj+pyfFgcIdv7410IWCdD/fTPa1Ys/MyyuwHfU/pYe
YYtWfEo2fsNk1yaMgS1c0m4rWKorDR0KRDdppYccvoUyc7QbfBZdEZIcU5BXXk8A
q3lGllMjunrgmyzwDU5Fcr9NvNCFCR5NbO6Vp/U8Lq0nwPhRuWmas6AvMgK2FVQX
vHoaBA/A2/OYnq0gMYQOLclYpu4FKBkUou/YB9SpN28ihDpsZHMzDhc56jW/x+k/
B6TiDHu7TN4jq2dkVUsaMxU95uEo6kTtwzsCZGJzn5Lcm96B0yJzStdln/rrcqGi
JCTTCtnaee97ENosxmh0rXQh8bOr/BW/9LRUmGOdXsElV7ydPMf1E0FaotVCR1WC
7zAStN8TvwY7aewxlmpWSz0vF0sj6f8n7CsXe0S9uBWb7y9dIPalxuYm21jU6Lxg
w/F1MHQxQFuFK7npapwQKkTVY6CGRbtwqiLDrP41h9dGP8FDSAvqSfn/6kQRbOIO
vrUCcSnD1Lmpfk6JeFdLY+2Ws7ePUSsrtWQpqeU/jQTjeNX338RSbsJ4v4FjOpAH
KMIAYjmImJyPSsPu7WSJM3eukSJx2hT1Hv2kSV/7sIweOqRszJO1LT4Hif8QHq84
7QT5Hvt7qkgKvUZC4WHOx8W87kGw5XRfwaPP+PLd/YDa+Qa485M0sodFUEtAOLi3
Ul4EKfzkaXf98ftS+wNDLqijYIFEPulkrBoTY70tdnFANxyQccuUj4ofZnNSKFzQ
yzoN0xojZcjU19Y6Gz33Ygdbn9Ngk3PeiwxS3Mo0RAHBZ2pBC4tn061O9tGIWO1o
HL2NKkmCZHUb6m/FJcY58H2b5qB/MdjK2hm3Rf8ljo4YsfBzo/2vAqnAs33+9Z8w
JvnBjCKJV/GELd7NdwFa1tOjalrgz48VGihEPXUNj4Lo220XwysLeaUlgs5NM0nL
tDfyL7G+OAHkFGxf0nN7wM9C8g3gXlRsUCNma3Lr5nSRwwmaZ6H0KA9qBkLeMp4M
TcpmMfEGopqzY2pbt762gB9/BO0ouj7ihuEnTDomXPNOTW5FWqV6ISHA80qxmNfB
PaIGOTfvaHLRPcemyHAeXQ16YJZ4p0XTDNuUSg6H30+jhoeOgSj2w822bhKCYnRx
IBPWL1U7Fgt75ZFnWGBMkkKq+n3j08Ie8gUmAf+TMCX+N0u/ii3YMUUc0u91C5PO
ElxE25YbGCLc+zh8yZLG1PALDq/wQhpCCdnxOsnOCvv1AJVwJ4Wxfnnzb5O2Xkk1
zf5M5VjExdJm0wG0qk5frQrr4nah9kvTLsimSPSDQRPaLEf96azjQYieOcs74zGL
cM5Ra+6TCVSE5nE1C3xUriUvlLj8ULxFLQ6eGlkt15Rpvw2q0ySMIpijVFnewTkP
AS1fOFixSXXT5w9ly4Z/Ge6C6eck8QXFEFGAOz3RQDZ4EAmRvHa3us5pg3U/7YHm
F2MqzhmaTw9ylqxSOQt0xsNVzW2xhTgGfi+laK51lGaqJt4XodXwDO6kpN7qf+Dk
3J/7Ku/xDd+ePj8zY8VFJnTNVY65ocZv4XsAEg9YwfGkmiOl+RMw1RM8WdTArvkD
ssTb1FSHMJ3WylnT7os2i1TuY7zpjoysUPJs7ThRCM+ejrdDkv4EN9SSRf1ety/c
Dku81i2nNA0mKihXfwMkhSFgl3fR0TYCET4wL7xc1hjqwstmwac5FfcQotpBVaI9
vV3zOU3MQen0YRwBsWRRJNUbJhiH74G4wjTljriUkPe5EB7DOvgyvfei1ClVePKp
LHSt2WJBpgVGvQT7FBNqofiXKyuLE5aKQgeqBvuFslPcbtJScog2VK4zmixD5X5T
9BKs/Q6EjQB/qFC8cRDZNE1RzgKY+QEPuRY//GKYnF113CsPpU9iqx8A4Z2J15tB
W3mNMv4XxA/+pTqQM1YEG5DQmtBdU0fHyYptLeGGDyST77O/ygyBBGbQOCtabDAb
HZrDVgQTCDFivJZn89ymEu83mZmE6QRVaWs9VAS4z0EymERr4sgcjKM3ezQMZvJz
zvSJh1xZh8C+Gs7fkWwREJa3rq6w1Ud8flKfyHHCPo6iO81Rpbxx54HXRQ0Hg0wc
R57pyJ99I38AA2nb2O98LLY9PIBf7OztRbwpCFpaVA9KX5JYUvGWvdHUlgwW1AKk
Uo91tba95as3UhxaJZYxINoYgIPzxhjL1voJzE0BZrUl0YK0UQfHpFIedaY+2SJX
pDxKyuFJLhP/p6wn3YUtTe3TknmQWy0grrC/BlvZWqDN/yyziGjExqUso0WFDqlU
3QiKEZAXLp/Asy5dviaajm6Lgb5/Z5reCp9oRzJzvqr71N+2Rvje/dRUI7TrlD9M
ZD7bokKdztXho7L8csvDx8ivSAx8ZgUNq6mivZx29vkC0WtVt00aGUsdGqWP8uYZ
w2o2nz8JthXZvJLaHEYv7/pT/+SNtdHKs76hy8v4VvbR2ndSfb06vMLBGG4CjVJz
zD6JmZyWX2oKpBBdAUYYTvtXNQN6yrstWu38JfRRZ4MGmV1y4B8717LIwVWzuOyR
Aj4BcmiGXqEswmGMJ/Ovh2TnbmvUZg3Ezz4JR5/J8hOd5deZ0fhcN+JImRY+KxG9
g3zlUgVpoafXBhZDYceazS0/oKEB94xRlR2bgAsIaZx3JDbJyV+9p8cL67uXQQdd
TJYta04wYMy126ukszxtdMuKVfEGG7djxA9aLpOepZh6n6CXxnberA5UmpTwP0WQ
fwE6/8HL+5iiVdnr73/7WPVGq4ExIYXi1YLBqTEg4SMH09jGIDULBeEEJoVxTSlo
iLspUySzwRqxGggPzxsMe2y8TbXfUPV1xS9Ki1cFRMu4VYBTO/hYT+/zl67f5OIn
RO5IXGYUqZrsVwntK8FsK+oHvUgyazEEd3UqOirdKVPDmqh0Lp0Tf+SyIBwrsZlo
fpTTEymJvZP8Pm/u37I0x/RHEkvRG6vVGgaE+hKEttnYwzs0yBa0fTlZ21xH7UiN
0iDmZ6nntTaIV9bYRMxtKCJMW+dB3xaE/Tk3IRJmtmfmNprxlFTtLWfMBYqX2hzU
A36EkALxkYStPaaStUD0X8JzJwUXU3TwA2Fho2tASQRtpvB7MYVJ+KeK5mgbi3G+
cfuL2vsdjQwvnt59dBS4CprIUv5dkOUsqNzLECu4jmI=
`protect END_PROTECTED
