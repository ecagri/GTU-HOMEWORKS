`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4JdZNayONx9Heis4dBAfVKHqPd85hXoGipZt2cejEatJoIHSp97cKohpL6V1YKJ2
amsnbiH93Cw8X+/dVeWKYYfBsM5aTwruvXCRDX/42oPIzHqMGNqmKORnYMh9VBnV
sg0s+THYeF8/PbTCiBycwnEBHkTgy54kyxC4GQV8UI6f+JrZ00b3ZMC3eeXRimSV
+oBo3wOH17uDJbzq6Z2+IvBe2evsHRbg+qFdjbTdSC4oQc953KRQQAGnzH8fyxWe
YfMuA7FRLq4E9Cvr+kYA+XO1L87RA7VOvUJ9SPH9SNVM2p8iCBTDo0z4gS+9HePZ
m7ImKs6ikYBS0XgOGRDZomeYMkST/fpaGmih0eVkksLB+j9MTau30w9vNTK2T5gz
DFCVz52snR9txOvad//EMq1ukPpR/NWOK6MDZqXW0IUMqxJC3xXtngLZeUtzAYff
meEGk9sK5bunui8+YNScbV+VaovNBXzqGz4Ne37lSL9elc76GDi/KsUTIc79zdJu
qFF5d/NsD28ygDnZd12Smg==
`protect END_PROTECTED
