`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ql6leKjML37JD0sKZp+hCD1+AEcOirBIaYNVd8Wz8ty55y1VK7GOsHf0ImdGSGjP
gcljlhlgooxGm5sMVbUWZOiAty4cBK+Zx1GO2df3JhMk27gjl8kjRyvubnB5K8rs
6x+cTPnayktHGkDV5ZVTMzeH2KJkE+yPTGuBITQx8tijHPFDUHWBqa47TQl0xZJ9
/xDYCsMkSjn/xTjfYGdxZ+a7N/jw8ZgrdDjS4Wlo9e+FScjw0RAqAcXgoILEw2p/
bJErE6ECQY5UYYYYFoO2IAnCRNBK3w6A7eSL7h7FrbD1OertUKLn1ahN0/lrLWiO
95u/ubVButuGnCO3EvRuy5bc4XzI9v6HhrAPWpfioIDfsVDHan72Vpa87Lcugk48
LmJW/Qr/cf3HuTTVXcvP1NWNuSKcrQl5vPgjid6qyaPT2ydW5gRhwc1YOX7UwoSI
mthmeqDSIBKWbeKcLR2bNNjU1JNR3JNShO2fzyJBhl8L3OOi9RXynmgx7HIPucyf
8KwX9I9PAhg9ww+eOZZewHXnJSm/W1OBs6h9kYMTj4jmQG3RelQw4aHyYIP6oNSx
LEFWg9z0ocD0KcKiyqgJ97g9NkG6aP8KUdQgAhzQGkJ9KuTCnw2M7Q4bF/pduant
IvwhIFrOJzPVBVGs70EoqZrNy0h1ijRAeb6PXY4gn2+o9/0PuVhSa80i6dPYAIk0
C9ZpLWmOwf9AaEt/lcj1HidJNjlQ8zgNVX8czhLh/GlL0HRnOe/+TJjeylWd7YWA
xawBVOfIJ6fIyJJjcW+5y4mzG8iyj7sreYcLdBrwlQWlP05ERtGgUwKx8YEgTcFd
+p85twehWzFqRxBlIW6v1xluxEVqZZ28siWditz1cHzG6LYE4VD409pA8BOe7GLo
5HR6W411RS+yF82JJ+Ni/z2OjKjizq2EJqe1Ce6tdeVjkBZCurvdqqBm4fvOkEyu
3Q4c0NMXAg7wmtnnfRy4rZ/aCYnZZ/9QDaegx7rNskszqz66HaxK5LCIyo5bNkov
ACEzoL9AM44/Oni5mKjAGljoLIwonoZ7iMNWynjIXSHShCFqBSIhaZuGZJn33W70
b2sY5H7cvk+BFQNapdoWsukBf36F0d6IzU9EG07aEDUKxrVus0U+FKOGYek4FwQB
tDA5qGIL3Lp6FdVqQI2CFnrGJSIivP7q55/+EKrOa3YkLa5XSpTa13HNJfE2qOZS
KPl8IdJgVwBNz9jpQ7NhUNXoqWRK3Hihd5XIeWQ5PwvhK6rHjgLwzbz3rP4ei94o
ZAGJ/0gGt35EAwjANsuw5tlFSn/DKXViDWbmvHrspxFpyBZ5Q6fdKK7oxV6RvYw/
7qhDn9OjqlXcbpm4rM/3qdBLFHQUfwQOic5SpWRd9BZpPeFymgJOd0PYKM1hq+J7
hFIK5kS/Rqxr/+ubsE7v6rA3l/pAi2tXipK1uGgo4jiIk2D/rWtbnhak/WDeDdk3
a/DXlMKrOXnAtDkxQhbDhSeYFs+4oo+qHsctkRkoT+u16AMFxuJbNAi4dEfCeAAf
FT3j3atEazo+YFb0p+JYD37d18ZfIW69R9RIW/ryOKk1AQXzGjuzI/yek2bLJXx2
ApEqxIHw9IUHJ8bm8so5G4HclxcXo2eca5y0oSGY8NLAFe/0VaenjJMw/ZXPa3Yo
KqJKfqbmItYcJ8vdZvWoOV22bBA0DAVyR1idJVz2EMFB+ui4ykSE8xt2cn9Zca3O
80XyO9DUW8Enq+BqWlcimtk/Ku/iG0fdhHpptAgk4i+nbyHbJ2VCAr04CYtQtXsM
q8cy0nFW+rpBUPLct8gQKDKCsYq8PhNsz9alqdILGWPbHaveJET/sWgQqbeyHMAS
V3TnP5u5AH5JYT89Vtu04rKThjIIQlDZ2tlB7gITyogl8H5O5nGGUFQTKxq0EYHM
F0vSrbaOJUZiOX7RjAjmaJSZ9vAZ3udTwNY8/oo4q5ekqVtmtDEJrgJgLlOoSJ9f
gefdsxy40K6OhT7z5oPjzbmc/yXtPhNPvrn79zye11RyNcFbrRU9wZIV9bWZCg8a
MxichkIyEKmBDIOiBRBqa9pC9/TyJJ7c1LfbVt3M12hBZfMEUrWMXLVTluirhaO8
SstMAKQmFdurcxLrCo03ZBm7GcWeYeE4P4HNEIn1so1V9GgQbBapmLuP4Z/SBe0A
wXp2dUkBVrgFJXHNDIAZtjOYrclNI/BAS6WQr9sEL2iUssAs/jQGxj8waw1xFdsX
YA2gGo3Xg3lGtPHcJ3UhkCB3WsFuLDn09fayZvwXBcipl1lsUDOd3ixl5cYTYkWa
KPz2ggJE3lT/z1UTAPtCZXYg0Cd+AHF4y657/vEHlvXFyg15PXdTJcBYBw2wkHmV
R8Y5POsfhBWzdPqpwPwTcP5YqW6FGxvR89j7vejB+IYORqdkt7PZJ2ViLujcYfct
RO1HnOkH4BEFr2+vJ1ObhfDP0LNblLyIMKSIY5PTSJ3REpyX62Qh2WHGZDZbKyR6
093vuQMLAXtDnQCQDE0CWKzUFlFPNRT0cP4UbkKTe5ChwT22y4gMOJUIgkizumYM
eUBKlNXbHbUriGQzSEom4hwIL/5dLdgSZb03DoNZrnNwBXBrtIeQpS8TdrwLNVfq
rp2LbdpyopMqGgupq1Ma7t5bWuENAwuIL4FGftGnaOsCItIKc81rvHvVUMTzZF8O
t6e34BjyJmHgIAqtdx5o9W9enCPe8thAuGh+R6zPuDNidzhWW3BCfM5i8k04qek6
Io3X3Zikxi3eWEj9zPoLAIjC+AwctHGWayPyUz4QOGh0ZmFqdFyqC15hP21KnM0p
u4MrzmWOgBaWd4iLS+zTSt2TrSOLAsKNFsDr5B+L1B27EjriYy17f/q0UpvTx/qu
9Z1pJeZYB/oo2MWgT8MPF408vO3Ve6lPjbFd0QCTcPoeK8NICq/FU7XBohNrSgUJ
t/l73WJVkXaEAFj2QJMdnVORLRW2KP+blYSXfVn8Pqs8GV3Yzb+flqcZg4N54/Kz
uzJSyhL3XYIAgw7UKckiPinAB810TTFMT0nFxCgbxV4mG/bBmSCvFmRgxVJV6VA0
egSDodoVL7Ab1wrtqyfRe9tuNZgrZWkCvuAcNOJHu+2BZ8QJyzF4D6SiIXt/xrLF
t+Fvqr73gjCp+k1AIQ1Cf6ffjRvjI5fHA48ra/bB82HtshLeL+4WbUr5LENIUb/v
XicS8kmkNSOqgGijcNMStNxUOeszHu6g50kZYa+TOk1zptDpnjtMmubTAty272jv
v/hB4gLIH/LAkZ2eQfwSX5tEGhaXNqslhMsLrf2wmDB2VSE/IBhfHrSwc0eUV0XC
OuQyslwxzHfqXzz86tNoDCVJwJat1yk+AFc9IqQ4jBOOZnnfi0mw76/dQxpnNTPJ
gNMZmIHk5yxb1H/4mp9ljyVz87BsjlppWFItZN4/wpkna+l/jMikgu4ifh51+rSN
OTnf5DCY/zpQyonziU3RU3oUBje0NuSQ+DT3Ng3CdI9LouBND7jkBntN5EFJCQIx
6OUPJjE5AveuscfXoRw7RNHuYXbr6d69fVj/qv3QhYznWX6yogvAIlU/Fbisaxt3
d/N3a4RMFKJPDVk8NpAqZ8IlJYNWXnFxXbrziogP9zYLj6oDmHiy5qBIlCNiWwdc
zMtvsR/aekXoFDlhnYCskYDgwnrLLD7z9TD1P//wW9LkwpCnBf5o+5zNdxR5fJaU
3gFDs/ug98hDm7D5gKtYIOlJiO9YfU0UsrAFfr7moK3VHsRAOepzbu0z/JKhxflS
bVItT1yRiBNAo/2bwVUiBW69dHTkDb9jyR8rUi8Uu2Vr7K1cvE9vJtisOSfrLkdW
mLShbUzqygfKPn4v3AoZ0rcx9/kycFWV+5FjxJYo/ArKzRweZHhNj1W2rRL56cKo
j532swOWOiIRcDiCkY8Lf4NJLvuMj2klndfsXT4DXQqSFzYqCEF1E1bfgb4dqPtw
88SB4HuAqAZP39j37N2b5Wed5DMTpxemBCAPcfrplWRNCt0+NARQpWp+Z9SlrmHR
8en08kV4zHn4yrSXWDjI0ax+gZ0i6iGXzuTIbFlLjgCm2BxIqopBzAhO5WAkb3DB
EEEKRt69GvPT3cHNAL/RH+YO3qIELQkDXlqbX/CiXaeQS0EQUSPz1dtscLhfcziY
B2U5snRdJxOIefw3hItO+l72ntMEGtCiO+fpYevWMde08NDYNVMFjKTQJpKNc8V1
B4fGTSZ83OJQmweau9W1rO/YALz31q1t6dZen/oNcK7lZW6gRuAJfd3NvK4Ndbcn
6j/0S/3JHCixjEFimGyAmQs4V11sAYb+tXrxiY7t820HZBu1LRYuN5RmnXZkFoUz
PPUnfVVdMpEh9oiwImnv/i+PBdNZjFH5VyH5VjrAjfkOx9riWDusDZZkV7vbCr/T
Ny0c7MK8QIFMZZLBBdhuKT12GcRPf20t+qAfjVe2K6+SiWbweaHeIW4Bb+9ZdYKM
ZYSgKcQDVQP6VLhsQzB+hBcCLS2JKG131JKVIdE0LIXfQtsT7ozNc7z7q6es/XmM
8v7JxXYZdqpGok4dK5VVU9q6EHNz2nPySC1vRahKmAL9EhslP4GT+WrfVYP/4eHz
bmod7Yj4202ZtbJTuGMAMcV+PmbgXcKtIWAd5mkx08PVoS/7X/8kOSzEgQBaN5ZE
+ubrzBRTfVMWZ6WtuWVKESjUAC0iWz0GGghbXVStHvJYsDA5APyT8fZ+KOUwaMlr
4xDJHDrNYUnTIUWgmYNvpkTwlpUTa2wgUqoe/nYrnIHJUqoVFCY5M7fTZPOCX4gA
WiiDAK1mPuCijsSOk3nu2zHhdbged91POHX2TcpCrycPLxMPsY2XIf+LE6lZWV5D
a8Wbi3tKFW3bZj0Sqf6c88LllTBss/+Wxd1MaiE2XFYnA4+m1H7ofk+6tcs+Upp3
aHRUCJGWkrWK4lgjLAO3KFZ3P711IM2H+QrZWJPcljgKJb3RSH+RB59AWuRFr7aM
YfoMXDN5Vn3CioDmB+G2zvahp7wHFkrXHMPnNxqISkcINTTFdz323UDlbk0UcYu1
LxNyV6hRvxK+AWJRFXXrd8icPyEZoVbjfpgHQ482VEWio3STmTol4unckZSCXWuO
uVykP4oJ06tw1dfFwBfCPLqCPO8B5T3twjAeR6NHZFKQkrZq9dHK0sKtFL//emvy
h0v/NjbU9GzdAHdXQaTnXV+haUaemcPlAgaZxHRoXXuxZJ7h47Y4U39ve03aLSWa
+egNM1hcXL6hS3zR3ze0koYyXacK/0qdjOQN1wnw6Dk2bNQvLf4fT9/r+LCGuwxb
LpoGq/8iRqybCjHKHGFrnIV71oGNbgR0wzxORTREwzbxC3nmTIadISN/GQ9AFWdb
lx5N4FbB798W2PgI4v6IX5wFkc2wKHdTMEJPF1GTNS0tyMPGb2DtiEOQmLPOJBDJ
2cfLfxtpBnILd+EUIxTLR3yrA4v7y/6Fmrana4TJPON+uyjZcj6ry4pdkGv/s0dV
3vgs581QMaUV/U+GFW+qw8SAKQDMnXhSKXyt5ftUhVaweB8JBO7KGHuk5tJT8Df5
d/rvR+DSdALGPePWE8AX/Os8QTPOFhhVxEulWi/OK6mUJnoQDrTIauBvLDrjkqCW
UQnkdhFbG0pmv4wjy5TEb9HSADR+Ov7a4jgxfD7yE3FqJI/uoT3fE2X2YSbi7WUk
iLdkTnai+/eVMm2WD4FfrSiFFFiwc8+nlTeAgtEEzvbeosm7rsSN0Qi6qg4UdvlN
R6nYIGsC1irWi1R2As58WCRq9T6Uu72xirJrbcf3D5kn0kAi0RcF2XF5n4EL0YH3
qOp0BwC7fqVbcmFl076uE996LvtXJfoHbJ/g2/yeSvA2hgwbY1+BDDwkeZf+wbyn
WvndTtyLynUu9eft2MlNDiNv76sWV04B6CbmBP+a8hsmz2D6mAA/ELJOXRmEDm6O
vva+hO6MyJzaVc58NdTzNijcS2KXDij0yWYSps4FDQvgTlcg7llJwk840nsIOPpk
FifrqT7iGqSF+TLjGgjSoFkOPBUvIoXJ+VxDYCptLu9CJAbtRfibJZqNXjn99AZ6
Zqk7RvHPiIpvm1ofUW+ktrGk+JqPd2iALu+qLsD8s37kKQHmtkzC5Kz2gJQWUi9n
Lht/JeTLSVj4w/gR2WjQx0/okcwaYlP+P3k2O9RVQYfdLQF9r6qRvBMCaqSjyTiT
flmrD1YmowUNfP20ZPtpXHGymWTBWnWOf24yqZ2HQ98Z2D3xNCVqV2/leVDV2Cb5
0OGdtJ9c1THflMGEicglX1tFbu/5GgQSxicIkUBOa4GIdTTA7TZFWGmerpLhcZq8
henbUnDvCRbpGrhfsThku1mE6WGnx/DUpHBKHnHgGklHDM1bA+389iTuQaZKoqzy
pj5ZU+3kvqDZpDqXGytKWkeWPbJ7QomvJ6lziNh75QcLTWceiJvGjULFo2t3FbRr
NUo8OA2HUYDvXaHDhxZ8ZZdMvgXQCDjP/pFqdb+4FoeOnkgwte5mQLuB1r0e5lsO
yOygolg4cUFKRATTIuo78xG7VVK2MMy/7K2EyFCQVbbyWgaCqiN8q8EPbF4ONhyb
HWT0vmYUXGecWOTcr2HvTZ6B3JlEEj1eEBesrTleA+3f+AEEilfY7UcQhfOrdpkq
fOO6EyOEo3JChfJ9HCEf0YYoa2cqkXY7DAfNla/Zfq17hlFzWNdWr63QfNmn+IFh
PYxlxyjw0EI0wxyGkJB0vjI7ZV3QejeSMsB1cELXetJQVHbH1fJTX1yP4nPvVK2N
L7a98gLGm0cQh7l1/2xAvQDdOFQTyuDN4tU7v9u1MpFNW/Yj4kKTQlWY5YZyt/Rd
0xKgu4MOfOet6dg1JJv9FQ97Pk6fr7Xp2SyFh/d5YNhFJ9Kv0GjH8015tI0d4PB/
f59z82G18aQ2Iqm4gSIZE0aqbgqzLBaptbBw5oiv8VlXvfF7/SNWFb4A3BU+1lei
BNJJoU+4nSKJV6jm5ikH3n93l3cjTZ+DNXttbI4QUjX2CrFw5NAIcHzHoCAfNVoM
foFCWWetV4mnNwN5OkFzaxvAU8mDyz1rZi1fG+iwXK8d5M6KXsF/I5AB2gHKhCMh
K4rOIG7iU91pwqk/ym5yDQ/KntIc5Pz+WTRGmR8cI+EhnktIfxJNMKosv8D/i0zJ
Xx13WlRWeY0Muc95ESUY/eMmoUxGLTEQkeqA5b4vYC8RGhMcb4WQAoMupa0hnsSy
POpv+aj4NClj9Z6/4OmbWcjq0i3axnLrRllCD3DilDW3QKs/OjokREZ0Vd6fgbfs
wIAixdEaZ2JRh+Qz+FLnGJv7g6uh5oH090zh9Rz0BoKopDmxYys/A5Ka+PwYvyGk
syz3d6pYYjjVmkQLRayorGpkovoNFjs4hBGK9+BEF2TqgnIC1wAAY8n5rmsZS7qp
v9FJSIMRbU3rLObF0Vu7+lOw/Jl2qC7HXLMNFcsPa9u26GBDpZw8imveUmb91H4e
K2T4w0brl2k3JjAoVMjOxKnRSDWozPEOiuF4fhl/qS5HOdCvqhCxjs6oevEQ8ri5
h0tAVBGSb6Gy6IlZ0ZVwGp+r2516D2K5/zMDBEJAbt3TpziFOCbQpshXcoqU2ndo
B8zojoHV5jTR8Eqona8QLtf8VkVWbQ57aaYRVwMqDKewH7oXl7hIbTigoqKz1XfG
gwijh+QwDooX2jq2U5tpZ/GsY9yG+6Rj8QGw+XyA+sCXBiUKZAtbvmx2ZYjoN0/d
3lFaRUnZOGYKWh6FHIXnHviOs91ipidUYJ8dyQbAJzdKDU0cjKxPJQM6tFsAydui
kDf3o/rSbPIJd818Q7c31BQjxqpeD2ExgfS8nxqN9ejN5Rfbcg1DPAWQhFiZ3BVg
4MnTFCKXimSn0vvWgP7KHfKKMqRvfo6LxrX2yKJVBdVcEx0NXUrFROFzBpZhvsG7
QQTjGuzLu4nUHDxgJG5Zpg667sp08ynbDdLbHHSIzXZfh1cXX2CUK2g921erZiQW
cfMKoHx0hcdHcsky65zEWjKElA8jcBFMdxCRj8CBn3o49nOMDZBGQDI2hS4MFNoV
16B0X66nCQLzbkH/VkQMBepM5kBTzcZDkXzSBzWS0Y40LQ92OFHoAV4fKC2HOmqK
rf5IFdeDEJqMlysw8sOn8zaWLr/pDwAQD32+fIumh1PQf2aTuKBWxK8vMsL+LwGL
Ir4mjmj1zUNC7oi02qzdx4wOllmNJDUmnOSv9PxyD1dVfZN2u4EUUS1e89f17eKT
jVn4Jp61jL5zVLcKFtYtYSpZqIHoVjOogKhZyIvKd/jdRzbSuNHLyAEGBT45lcUZ
Mzmbk9azLNUPieC6MloOQjMjBrFQ8/uJ7x+yNeEFcM/TrGdgybucasKhMNvPYPLr
RGPGWi06c5l9nkQG3HYTG0KqHx4uIw+08KieROzckNOux911RwN0KCODZbg9aELt
kfEz8uybTRHdNPn0rEZ7KlfFYu9Fei2aN23n8hdEAslKyH1HvAsUBsJQy3KHkONP
itxRhX7UFwnkNa3dmZfepIaSwK3sJtDaoyvaet8pn1TGkohTKVmz4feAwKOcHsgX
IpnPoWl/S2dPMGKmZg5RAvkApuVi3oN+YgOEqdc+xFndh9iEUqNd4vuExc6CgC2S
w6ibpfzL6dYb/XY7lXYz32hqJ8O5b/EUDC5SOX1xBIirzKHoRs7fWX/fYEdQVPf7
IBD0HGRbtL8f6b3druX7xB5A13GkLSLdSuVJFCVQCucXrssWofd14DWFkD90FYo0
o0gCDIuGeW+B701pjMxZarN3E3aC3F42/04YVN5pjylqnxG1jZcmS4sxTU/L2i2d
uHm6Mfo5FbGlncMRWXKpSTj6jzAdPGrrfJURndP5OozRa/rCVOuSX3a7D2zhz0lD
VnCTcemAMxA//6hiSOP2lFY6O99lPFgWRgg1cOgb10zVsQ0p6t/mWYD7Q88YfRG+
244QedQtcw1T6qJX+zgrSzr5z7Zrzs71lFLaVoFVxYfBU1KuspqanQAseA6XiG9D
lPwt5Js+lkjZA0ESWVYRJOq4hs6EK7qp9D9H49df/UQy3/09z1x2ByA8ILpLmtCh
xrowgtsJqIvO/iALviFFrcjLwrmicaAPl7KRWkacUALdvu+6aEys/eXkyZ30l0kt
WlX5YEi37xfLQNDkn4gvfLP2iudRcbOQEIEjEzPk6qfIvwpcIpjRvzwj/sVKB5Ge
+Ej+NslBJb8PXFVFsSpZ3tojT8uJFczIuYyHOV8HNYIflykeLJOqMEekX9I4lz8s
RZGiejSo5worHlVOQ9zqQ+kkOpgq2AU50tqS5RF4hH+nrlq4KVDQ7OjSKtY5Ewcz
kDOnIYu87G7QYERbG89nJ5v84tnB8IzadMH3ZwXkvH8uVqOZVZOF6Zpu+msD1eHc
qKKdjCFtpHt4KozXYri37WBuuf+jyagxXDrgGMQb+Il+mx0JN78Y4y6ElIZewz54
6Yz7asVC+q4V9adD70npZ60keTeqDAKTS/bM8Snc54XzT0Tnzcc2fvgPk0iArw9z
t+VgdvOnzP0x3qHiwzqMwoRegkZULNfqyMhOJyybGNx/Q1hweNfC31v/noLA0s/+
oIehbdKbHUpiJthQCAXT7MnlbRONioajc14uj+78xbJD+A7tVABB/DKXdgGAupK+
hQAJf2ouY+eGtvD0hvepTc4w5YBiDBwXD5ICEdN7/e6LlBcf89/gD0wsz2wS+adu
P/VyM1Lz0qyZnzD7b7B77Ft1heNAZOF/UEWDoj05Oe0U4BgSuoEGRv3TSz8Miyra
q+v0tR8jH60iy/7X6ChEiVPb8RjAARmK3kAuPdrWEHEV5f+6wH+VqeVkBhq9UXHY
LgJl4rM+vX/6JvdBZLW1/qvvwYMLMSWEvVorywumd9SiMlUs1pnvhHR7JO+yI/XS
7cVS2VcbshN7yB5mjQ/OlR318nwJa18POzHcVssqhO/9S9YFWM7jaHY00PaOW1y0
/FHTbDQOFLWoG84pfPK7kCtcmO/TpXXusvWljiMpP2XsFpJ4Ja3208YxMUk9UYKV
qR80HLMN4Fsystwer+notziyYYMinYwhQMkAPIpAJK/OVFjBELosbQLDhPTDvyTX
8u/JDs2X8n1Zl0h9QUyPkzMdza7CoGCRm103SHxrtGitFdKvpUQly9VNOP+1J2F4
y1Qq59kPm3duRyza6cUpQdo0wtYyLVap3Q4twVguYoYPdToZKFJ2SAHkje86BiFz
JbxNouYEXxrumTGhDfVlxi3llD5BTDb9w9BHDDt3K8wnLt7Cj8lV21Vl+FgOHYHA
4IIp5eSY3OGFmOwZbAiDJLjlAzBwIhpVgnRdW3XX+LOj04y9pzwp3wp3gqdYXOfF
n2FJetZzzu9g5xCkXiyovlBhFKm/e/jrREBizCkM3Xd7AQdC7O+ArFa2gpB2gqQG
ArmhuSQaWhu7GGdxBuod5mQPqcoKRrDBRg00ZJP1PkhRl7STz5LKvIN4gYfTrvvN
gQadAkT0s18xuP/BcVrNCQ==
`protect END_PROTECTED
