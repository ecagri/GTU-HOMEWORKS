`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LWQ+CLlL320g5FTzIajPp0yVFt2thSNHa/L4sYHgRwUpTOP1WLl8VFwJzZCnNf0k
kvusAW8Smxuj1PwUkZj1Bn/HiqROEBUBlO9Rp30KHv4uwG+Rr/YnW5NFeT3mxagu
sxV8MQgnStqeemM+7ldJkgOTZ5h51w5M+CF3oYplHNc+X0sFnKP6FCpKi2W3ojST
122fF86XagiAg1yPc5fuPeswRRyX4zUBLsgxIkdVnzZ198RAlLw5ZOpWfcXo8fsJ
JQOwKAhaf3tT78Utn/4J1vqQ1HwyTmpRJBqcrEyaDkI4RhyK5y1GBNyukmvBddxs
l10yl0L3ynYH5Gro+2vum/Q+G/qaMtFNEu+kOd5wM/b8Z/Idm/xUGnnkHRbkhjxu
Qrlesrfv8PEztSUPzFrR7NIYq2Ff4QE+IOTKILf3ciSHTrVHY4iderpzGXNqjUEf
dU2AaUEnYbAVevupbxoQTQXIywV2cU/5mtl8eAb+XVqMdyUIgQkeC+Yr6ipsBjTu
IF4INR+e9FfTvRoJAbNEc7IfcqoSdH/vh2eeTrqCRohA78fYzVhiaXSJITeXKaLM
/IXzY+LA8jUjVTYIAktB7b/ZJnjPEvG9amFyfMq2EEuskBLiMJHdB2QlWmQk3hBx
PLOzluiZITjDNIMDbj8ya/kdxB1GddqmReCMXpDCX2qXBY9Mf5MVjmUswUooN1gZ
4RjC8nKFT+T+XDFhMAL0mg7gk5d3Pp0wjz+flhelqp7mM1wD+SLwEeLf+fv9n7vN
B8VFj3pEcjFPBvcv9Eglf6DTXOgO/0ayXolgdZDQCcaPIgJoh5uP0B6TNEGZ68CT
9SVH2FwzW83BiRAz/puBdB5ZwFfPySxHXznhTr9uI0aUi1Iv7/obW/ue+9OwSx+m
SUZU6SXvASbom2C2ckhciwmyraKNxF/o7vmbfrgLftRPigptfb8pGT5wi/BMK30y
9xITKdJCR33n8Ou3agwh4W0byf41V4QOlptYjA3BRpnzTS1fkw+oXQMxGev6cegk
MLuRxjDovlGBUWF9G6gEeSTFaZysHCRjobHEUQsrlPpXUJY1C/Oe6rwNN4wx4rt3
HK633WlbOPjEJLy+PJsn9KAGxmI5St1+yzekF8XTjK1Xcd4t+46tlzFCWHTVzNtg
yWXg0CDyUmMdHM9tQTfQ6vgs7bhGG2B34O88wJ+xWE0Z6OOz3rmdRtRbHmXBnA/i
TMbJIKKGIKH9HI3dfXzZzl5+1IBwLfxjnQyx14qsg1DbAzHdTRdMEEt8I7+rXrgd
e6v1vj077e62LFcCwtSWp816FSfOb6fsgg6gDRgb84CNu3jh7cjaqyYr5kFZnkb5
nYHpormHWuGPSmzRQoZOvH7UnI4fUmfVHG9Oo//WrD+ro6ymMl3SBZYIw63hwuJd
hcFf6x2auI/ZDS+3Yp6GyF3ogmwYLjRRVGazrhrj72Wa0/BubS3Tn0nzQq6cS3Uc
t+ToQ1TuV/xVdFQ/OnQrKwhdvYulBQVPvLoRqQ96W+f1xedvZ18MGck16+bbNN0l
7QlX7L3lM5bSQYi7AcmMxQ==
`protect END_PROTECTED
