`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yjAixkGp271coPm003UI/lh3kNndBiY1R8412k/JdDTOoI24uS/p/WAyyjQGTbX4
8o2HaOAZRLl9M8S+vsKxH4BgD8VkJAvA3ghwViUlVAvZnwr1C8dVA2d6txgOQv9c
f5JX++Gq1zM0MktWNM7lJDAg2VQh2RXG/+C7zxLHW8Ld2Vi0NtGmddhbTV6pQ0Ex
BtBnTcteUcJmgBRZ/FJNSh2ZyDKT6WPnsikszgqFUnf6UznJ5YaSgXGOvek2Ad7w
9rMXdSgsvYUKq+uZxkhFt2V/fy7VtUGfOrbb4w8qzkyPwnj/Uaccyp/ddvmx6Im0
BREyeBOAT/bCEIjlzJFzGKzDhM1b2Wakv7R7aOi/OgmPtL642uKl/c3C1Km5N4K+
8e5Wa9RaNpICftPvZjnL3KPdxHbrLSqtq+3l+gJDhzGqijLk0eOapmA6DH54QUnL
llXYe0T2jwYM8JJvTMXMPgJ7wes6tZjfBFTXb3rVdj1vOdaDACwXhgBeiXlUEAt+
/GFOTiNQF0Sp/leK3K7KO427ukmZ5lXDl+FeHAlsWlHC8CSoRvYHv+p32MTvNr8B
foVzkkVZ2Iy+Kj9/yuOzoip+pCcB2WR6+lpw9uTqXrgoG1iwWQf6HcCKKBdb1jTy
LR6aJ8AF+OUSkk43zcuywqnO660nYrUDDPjMENPZnlalvWE06GGT4aFxzWlsUZf4
gZuZWe9EsPfJZMk3NoXCENHhGzOF2MFJjYGJEfH1r2oBjCZSVxh/OUcqDq69VbPs
YaqdJyA2yqAPxMv8aEasESBcO92Zfk/d89UshQr5MohI+BrfL+aGMswpiYzpqR80
Tvh+M285TszUGTUAaxdUsrN0myIp/hq6MZUfLiswwg/EMoY3v/ce3D/htnhTy8Wx
x+RwBVZN1nAQIEnu7IK148pCFlmE6zHi+gqnNdqa5NV8aBk1Q5D/4CBzueB2tRIG
Sc9FsRDWL3Rgb5pfiLv75rpSnkTOulqzqwfIiqZ7uOPEdfNYhsY4A8ZTc7z0oAyo
kpsuiqqe5j4UjCUJrZLHxDHF0PDYi/8DeQnPpVeIzTfnt9Dt6NGPzRpoXBnmxLjk
KuqrQBafPwKJHPTlPKE3+g==
`protect END_PROTECTED
