`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
asElcmY0I1G31r7h0X/KXl1IXTCRRFuYJLkW8S2TjkGKIKfmbZNyyE7vNAHRkz/Z
G5eGJIsQ3EBBbh0a3h/AQJ3cI2IFBlf+XsgCZ419dGx5Shfb5PWurZKZ9nD8jvoT
Kninuif3G8KmJGcsrSgynUtKqVj/H7ErTTrUk7sUsfeGBnkWTUAuoxSVTxrTIYdG
Wn03q1lGTfSSqIhfL3F424Xoo15PfX3uaxgDMwk4RTvAiyRL44sL9DiACFSfTU3A
OhEAdxU87pUorMSDA37IV/gZeC8poWZSit4c61tL59FZ/ZL5gEvplzHFpQhqx6jW
hG6s5iD6USfkCc5ms8dH/o1A+x0s2l1dZALRJMQYolDPRNKSSHPwweMmYoChVR4Y
SkCoSZq80TAaM/AQqYf7z45cSmsQmmBs5/ulgs4dpHyKg7pz0D4RF4Qc30et/Rk4
nH0FEArxCKM0oVYWKIgcyrawY+vr+SunOnd1Zh/n0IZY/jylVn3esO8GmVsReCPc
8v90QejMBtpnSwULf59f+ct4zp8w4hRKe52HCR+VNZDMo9jGJ3WPDvCIDNse403I
pL3R7h5wi8TgfDZt7vmdOS6YiREGVW4n+JOCI9EG3j9HWKyFHH+HIfQENO8Dv0y0
AKtHr6fhzlZNS/3FY4wu/IvDrppSGyhSIpx8SK+FSF/6uEP0IaKMEzBipxbEZYHd
Q9T2yRSZzyfJYbYwxaLtD7igPgzZXgyW5M/bm0fNiLurcggsqY3xG2u+rHp2LkUj
POfXN8umYDk+RsfuqS0R0i4bE0bUa+NmiouzH0hQgpXayQcrUY2NgBRpBdDdItmv
F3BJzfxzfOyRkuaqMSKtYUp5UJPStGeU9xq9ZrsA/tPFJggDzGHmofnAd1nRHElq
bmGWX7iArySWUWG/F9xntMKz/UlLlummdA0egNENPNLOaPXEQh8RroMzrYScgspz
5ULc+RbGz1hgq5kIDcTyU0t9hIGgYq9CvJAiJSKOe/TI90+elgbpDPquBA3b+FpF
cXNTHDmoYbMbF/BgL7r4/BMPA3PLCKkZt/58I4fxu0xWIgGzv8VhM/R8qJxCkWgZ
dn5GJ0L7tABAf6J04pm1JtEd1Lii3uPUbfw1g0azQtXJo+YZ78sEz6v0tUAAnaBv
NgLT/McosaD9uiWjVcsdnEDKieJqlCIE/5RpnKA2v0y7Is+Ak27P859UqOYOZxdZ
gjKE/8VhDqjJmllfqhnjRntdMBeXYaHhT84nk50ERU1rdLKBxV1PBO3z9u+pKzSm
qKYyjoZ1l+wtFNM2yODC5aJTU6ZFyLkkBYVTIPizVUOIbfQDFXcFiXrMoX4Ro65y
ird9qEnvesJ6cSjjHHZgyn6U1xKELzy0HsHf37HZYo8mPhGtZAzlFo2tuMqW4p2y
mnw3lhQGZ3GwuD5FnuirWhKVBaqFCspJd64sm20TvmT27yC/diz1n150Fvd/f0QH
vtgRRbZgQz9luv71psFg7RuFYF/8IsWqTuu4uakhE6BiZpYl74CeZvl/dPnSdeWp
BRwLcp08gyq3QJyMKng024jcfXmooCG1U3sV/DxetHWAzjXwl9Rdv81QP5M8PCBS
efjh5IpCPU4I2JE3b/CyqgtlqAzssTF4EJe7+tcXwwXDHCEQ6hPM/Pn/ypfB/GyZ
mFDu3K5OJVJTDM0p/1D34Hgl114tyTVJ9AGJLeVIvZKmvqrqhK9FvIRxhT1I5gvp
lPBp7oVOtF7qlHJ3KMVLEZgKTUIhNRx7jqlWRiIX8Q2axATdR2Op0SH9m6OBPp5w
fsRaTuVwYsksfVG8smhA7roU9vnXcyeD/lBNZyNgjlvrItaC7G5QO+o9D8xupCXn
szXnuan6j5dA+4JVcKRTKF1uMaovPc9OkIw8prd9LJwGtFhE8/p2TA1CLfmQp5sL
X1BGLlICqo9QIlJnrYW6S6Fl8wEPcs3dEFDjcX7DhxJtB8DhnuFClOtc5cxdyo5D
x+CdKmuNH5ax+QrtzdFX7A==
`protect END_PROTECTED
