`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/gNkIEo5p9W6dQsmbqIxzsgp/eQZOpwHSNsnRZuG5r7VsXhJ8Hz/C7xEM2OPJYrd
smSTQcn79cBHnBCoi1NKl2iCcRos8a5THH4d+2HChgmblgex+wyd+aHUGxtb7kGK
gOAsZgHal1axdwR35Jadfm+URiClgrM+CUtJeFGk0xTmLhh9An+Jtg731KE9t2oK
55pz3C4e8R2Rx8GO/jt6vuX2XofrTDmOb7WOQiivJlOo55cr0XLVUPXCjAom6kOT
i8zJiOBAaZoR+Bp4yBZu6IBm5D2PnnzZjK2l3As1Ej2hDUFOKpmEPNHid5+lo3az
Kcn2CkWC25O8fEP4spZRTlzuY9gwhBQPQQ6wRUD6JqMjBQ/BtXBRgEKsh8cALFTI
V0/dS3G3LlHUb6yi4lZVrrM+NYBzS9L/Ozo60xIh3Q7bsMAjMqqe8LJpzbxxX6ao
Zclega972r2ibJUal5pFGeOxH2OTCXIjucV0adMV6bMKTexT30LxmBeUbq+B5unY
Ng4OABNi/CLEoxfCOqK2qmiV69j3DyZQNHkbzubKiXHI2jN9P3L7m0pWX+jmCSmB
0Qx089GQEupHJx8x9VKfpuPq+sAWUSk2j8nMG0Sjp+MInAjRjWzn3DstqeC+c2Fm
SIGGDK1CNQaMMy/suM5odD/iONn1jYj8Jgtyo7m+WsJUveKN2FK3O8Qq0GqltY+z
mVNGf72SImLNVbirbKlYprnf9aMu9iadgowfQMFLBSlgiWc4uJqjqQ8n8XWJLWNG
admI6jZkfGjyW6M+Sllo02L4c59beSwHrWTfwhL0UmbGyo+Yt1Wh2SyaJLiVyD7z
nbTSQT6sO+sHuCpHBxybKa9qEhlM6FxTf4r28gNj91HvBoQi5a/xF6sKR0ZpYqYc
svKl75mxfgKhRndlaUDw5fPQxYpDlVIv07CYAblb6UiATAcegAsGVc/USGkUm49u
2v05r9i5Ln4UmIRCwFFlmYvgQ9OM5neAf03MgYZ7xKPODHHhmHDAsgMzdtuQMFHS
GtcHKIo1jzfiepqYif1Dnpi7x0UzKdvWSYtDPH1PA1X7zMbtqpyFJH6E5MbxHRVm
V7zkRTWuANypger9vdm8UsQGMqUcHAaTHn0b4/XrQFhm0XmjycfbioozYGkPTD0y
Ic2sYX2fefhDWlJtCd7QZ/V4hIg3Z0KA+q3oazL//FHr8/Epc2JKGRSXcAOyMu/P
/ANnU4KgSy4Z4SwBCkDGmhs37gU4xOtlrc9DQJwhWYRjfMw5740SiKp1WP2lLvV3
DstgXs9Ks74SWfDi6/wj3kDViMQKU/bQzogeGhUGk6s=
`protect END_PROTECTED
