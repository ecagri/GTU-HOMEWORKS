`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QQLil60/Ghp35AdzqVL5Abm1wJ2LSjRUaii+qEHIFW+sHp73ymedQxaqHpsL2qwm
1h8KLxelfMHfQr2bU4/I1PBmePsrmmGfnkqZ0pYb1F75JTq8+U1UBVnHkIgUrXQM
m8he6cjXF/dU9EYdRYyQV9Xiil42WbwZ/QqhpJ6GbKXniuCZ4bAEkPLqOBJoXzpW
XbFvKZO4yA9sD0RjOh4RarHzgU6RtmoUr3T6qne532DCEzmJtcM0Hhivnig8RAHD
CAjwb1PA1vBXy3ZopbuwtW1jQOI2k0tWFAx3iYIBef0grdYCF3IiGxG/5zEf6SEk
3cR4ynG5vJ5NcqZEt7BYntYSM2hVL0SpSJ2LS30oTXjngqFxJDCBQt63V7yjfy0N
MbHuHFbqQj4v04Do182phQ==
`protect END_PROTECTED
