`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HniNRcy89EBrr6x2z2Fhr6xVneYGgUK4KRG6Paub7zIGfdduUYG7SD7R+xbsUY+d
3NBG3r38q1BaALgmdv4lDJ5qNlkbVUJUwByvwIpqtsdau0IdwSRJ41r+VudmatZz
ndWO1De2JbmDuMb2HaLsaTiVVnwT9DHN7YnRg5TAhFUIOTBUJoVheXhWlYR8/hNn
TixfEdHXbiAz+zQ3rQjoIKSzEfUfg9tgnEMj7aYD9019Gvdi6wKQm26HyBagJmj7
yllXmx19UdF3+8iKH5cbC5iT7xWfrjnn4CksSicUUXzkz4Du0cIFDg0182L7VJYE
EjGAt8s2bzu7uekbRy69awJHU/aatxhgbbAUe15ZArbVdxOPeJv2XSBm2WUY3NBC
9aO2ouRSgRTge9EJZSDroBvGLTT53zjlza3CGGcJ27aink4Z9sEw6nFFkqrkISeq
S+9QGBC+AzQZ0JGzFbjHXcbz/AQ7MXHWghfcKx6/32Iz1MHbkrmRTacYOMiPSRkt
m7L0A1QTaDHcGb4rYKNKAaxTm0Ef778mXR4hVizf0JXvB+1fXiw+X0kw46s/rCoh
ZUEoiZela3B9cixsBIt0kCbXOvPbKfKj3xIsnZh3BqmjI3pXpUJxejOb4CkAXSWl
qrUbApoVLQX++dvc21M1qNhqqLLGmzI5aLNKu0oEQesp0JsRjWYuwKzNn+HS2IQL
XCVsSpOG5WXPNpA+gy0M7MYvGmujtI2rOC2bRmwYifUMmnjv50LPu2JhcicxQbtm
kktBcy/rcfkyWueoOv69mbc3bxnlq5L7DHcxW1ggTi4yRnn1cOQScDpzA3Cw+Y8R
Y966rlwipBcw3yqltA6UEHT0tp7NY/m3h5oqI4CY+yxQSC/Q72Zh3j8ROIaqIcdc
QuD7k9GSPqJOTByjjpqlmoWVoUQfJni14wzrSx2puMc=
`protect END_PROTECTED
