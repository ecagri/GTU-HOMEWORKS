`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v1UCPSd6ZuFu6sEPdp4U4RUqu+pmMSxXVmtb2ORSLotwzD3eazs1w2p8CsmH/j1T
AQJB8JaZCnWDbxHOP+iaPoVSC6lHoWRjvJNpr+nJypflVGvS5uZ413bv5DxR4s5P
EUxxeoSrxX80AcAJt9UwhId0rShbGzPsKl2wszysGvR9wR1Cby0cS9kNb7ikTay/
r+ZomDdG1up5etqvXPgn+e5EZDj/mUG7FMmx24eMCJGEyrfzt13B8dHbwYSJqLjj
uTjdH06AR3nnnFDRz0+A/9pF2m/RI1eN3Wvwe1h3LSYz/oimY0sseJoSEhEAjjMA
GhHGo9RDWvinlvY7vWCnTwzvSYs6ge9sDRDTmsLg8qOl4/VSTZYf5wPUjYfv28i8
iS9VRxSDT6f7PJjGqIueBFbe9ls5ErqA4Rc3Sk7dduQonUuodeg/nFK8erUWaReK
QxUrdq+Mzb4WJInq0ugMBbf8PxjGUmYlNVFCOuWSUNeq+z2sVOEU3WFdV2n9jEmX
yp+RqqBZK2cRZry0oa4EHOpMCnpMSsWHEZYc+4ry7ruB139nm5fY2XX6CG0Rb6jm
afpPXa4EpMZv7u0+CSzK/WpSMUN3shOdF0/YHI5h93kknDdDxSjxcXqQA4pURnHw
sRF3GcEoflKzX3MuG85DQ4e5gwuXk2RJMyeaUhXkrA6uLmTFeimC8qYzQIllgPv8
yA159HzC0/nk1Xis90cHfPaWhHBX2WAOvtc54+MOCtWElS0xlB+7f86tCWCsSDB4
ys0YNi6VKgI83GEuIfrFD3PemYL8OF1G9bSfIOjChFmCXWUrjaOyNkzFZXyoOtKl
1+UKspqu1yCPDTg9+fn3ZQ==
`protect END_PROTECTED
