`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sctEg6EFgnzapgQDziRjbSSv/EiDxDnvvjRNUe5lgdVFvbRs1nJ/5goJggZ2162b
mz9LcnXfdhtr8u41xJv1TNwpOmkRJokxcwyHWlXMwKZ//8+V8P0d6aTLdSSq+xQ2
P6CwQBx+MQ0u2+vevPv2y0Z47sVVjZMKgqgcCvC28qMfP7ZEGndH1o3vNBxLGZae
gy2aoSjhEs+eGj7Q8geBopTyUT2Vp5pRRzDfVvq4xmmjjkR/hSGgXUgvO06+vb/v
eu3brMKZs8e44s8OZRunR8EXrTmZXcEFLgPk0FIkUFAO1acfXDmrklTz8PY+hiLt
LOF4dPNK6DTpgLLzZRAw8Z+wnKlis4IBuesXb+xV0pC3k6o2dEhuN7oI5nMRBqaZ
t75RD8T7TwwJSboM8WMWtCLTxP+emQkMKDdQxPq+EXnBbnQ45/H/Pjedu34S92u5
DcYxLRPYtZjI6HM0g91Rkh2qIlgUsxGSol4suAI4zGepXLBytVHGm2cxUw+RosNG
P35CxlpT4KCwzZf0VCesDIVXsuumfPThcXIugEdJwGDvAoMfUSJDh3sotCWmkBZB
jLc3UwXkoVf3GT74fjCIACi12eqaeBn6uG7D4DFJSUtudLOgaXM9+nGBULYb8ThG
j7kNmQWdRVwfsNmZR09WhJuxT+tYY3g7Bc5BwChplKzPYmDjQrlERnlZcdXsrkIh
Jfx+GVRSiSDKZfyrOh1S3exLwi+MrqBpi83q3CHhbmiiHg6osdfG87iQfXaJXJkl
nJD/siNkepXS+ibh4d8hXj5wKHrPxIFkyIDFw6FaQHUQCfHAdIS4x4TlUYfCcNkm
AKrto5h3f7JetxSx5jsF4nB5JDXb+qfD0wH4cYKWyV31QsrCbgzgowBBJIc4wjyF
z9fmh7lTsoWrs6CaxY96+joxbmAXfMhbs0THTJ7pu/+bxjWv/dooDePal2cyv/G0
6A5Ak87vGXdXYw3JUIu1g+k21fSZ4GnRN6GUzYm4K2Ju5Ln1IdYZJQKMrl6loFgg
F9rxWFTpufzgELZ7k00jMYvwUpalEe4qsAUFlJnItwXu7w7bo2flq6t5HqrOh/U9
PBS7AP//5D1zQ0KcPucBOfG4IXA3NdfZgRA46sB1LTivTLqtuDuiXmTGpM3/Rvk6
qtc8nV2U88GvQsV9vaQk10x1KqJTyjkNRNCfA/TIIZTaVQEBRd1W0qAc5DfGRg4b
ZO2+3YClShJVpQ3nJ4Vc5bUO979SL2BExrSi1ZcbrS1OL9RwQi7RrPzeJ8C1KGHw
mkthhpvQtiZYtklEAg+hsjhTfopgCFWHkZsDIsB51HqegUlOzoI06JzaPq6FnzcW
ABtq/5wYAhzXXeXe3qiQ06pGGybf4hDIDe60ugbYmcQOpzQxo14jI4THF5/aJMGm
9yoNRNosjgCHZtaQh6chRz7oLi0BRMREaHPYk2IKxntZFvx+Oskk/JMKqsu6EbY8
ZOVkHPb3s9TaOCCAe3G2hKq7+kyG+O09Hww2b4g856W5LJ5e0bmWPY1+KNWVXojL
iDuxnmIeL0n/mHop6eQYwIQG8MQmO4bC660MG3FVp0tqRbM4mfr/TVuvCr3aDDVP
eaCFDXInStCGvDX0iP/jv3aEiWH5dJbthHKE66PnNIoypU9D4S7q/dciRYHB1DvF
9gLWegmc6nvVS/32hdp8Z1WSvLE3XSgf9eVDOOnx6sZP+RMieqF2Kk7vxCchCW91
iH4P+J++RLXgJq9Gsug+YeCI+AueFdfUR7hEG4ST2gvShXN1Jwa2LORRSlpiYQeE
nn/j/n09y7XZHX0FcUTojS6g8kQnOTZZmvKwWZdkqVbIjcZkqs+46YnqfhIq5lSZ
UMYa13s+N2pTr/tsCVY3ovCTqd5fyhYOY3aHl0D3EFwnGfMWjrJH8LyOu6epEkv6
LxpSTNaPK+9wg7eMCKQ0q0oj2FJhCYdOlxMX1tS1e9vQdJv0OfXMbonel5/zTu8G
+2cvEBU2Zr2W6x2iNag+RZGIF7C3r4SlX2C6+bQuoWk93YDKbX8ERBVoM/W6saR7
E4RUJc40cuvOKhhR/zmG3VIxphNDL8pH+4MPz58OakJlICe/adn6loxNxyhP3gLZ
qMvp5TMbtCCVzSU3zy1j/LSbjWXHIu2Lg/luqeBO/DwQGZ5RHuW4dxcMU8d375uq
q8ISyjECUKkGGFWJlYqUriTxH9a/iPYcqPBwWkibmBmRj/8e7C8lckyIKzABkiFN
utIgpPDpcytiwCqnAaWw0VQtWwduKVR6kH1VXPGohwNM6nIDN586WMPDFuqMsxOj
YaG+fKLgWtTye4bPb62F+xduV0v4wXk/rOCeHyfi5Yui9gYCIGlptdwopZx8E7bL
VRKWVIpZUjgD0oqwjHsZZwHbK+rF6LPWRQzcRhgEiOfVHmz40esGqKJk2g7OLRbs
yw/QjDcskksVHyK4dDYT9P3ayERohLGPD2Q/K5/3AZiBppPd632W30OnFf6LeihX
Ov6ti4vyjqK4zAuX7Nv20EOMORikRE/tONQX5sVD1cKe4s+MO7RuMaNg7QefCm02
vpnroYLguB2mWNKFyigUPcEivzpSjeQbTE8BlpV7y2zasG7ZE8GsOeU198eHvu4l
SblsZBULm3r/fBK3WTGuusW0m7/avlzlBr4nnrskxZ8+Z04IbfNc6RP2EAknoHLY
qI+E2QZPxmAcn++dDgBTVaAo2VvCOxHI8BXGXQjnCA0/qRHUrd0T35dY9M5aKrm2
l+FXc07Dd7ueQBr4JUahMW//x0WkS9skF5vNpkjACDZEHWYhn8Xy/FyyBVisYgBL
a4JLC19KtZu98pAuAhRydRwn/XaVnQ3QGnxTf3TNtPy+eSoEhztPJoDiMQAK0Tr1
C23bsTicoQwXnJBLUHPDb0IdTTQwvKxeCBf3O6/DHtvN8mZTfY/RMGnBmShIbFmP
LUCEegX5K1gWAmL3yZr3D7ka7lmr7mJbI+3glPR35NrdJ1QOEthTRUng9SzoVnqj
v62g7aPDUa4k70wbTkqwjbKUYspEfGk3KPrZvFPGvuihhC3GzDG553hkro+vJXH7
gEo1VEyi8TEIZ3BtQugfLHNcwieRO+TELUIJI7q1GSg674hFf1n+qguPi1cumkep
PM4tIhmDOAvGhCo3qhhC7kYEmLOkEEgn5G96C6pqekubgaSSdMEKQPgWUP01mD3s
WwF9RlvVZqAVZH4CoMdfaQhDd+RxvSY4qAzyQv/Ph1vLPHYBnZRS0EdRWpXWn2h5
l7gFiXzsAMdiDmixJX6ndhunzV47YyGUun3dvVd6DpcdLhquwxSrzUCqEhYiP8el
xuY8hcsanfIduWTGtEiwIDUBHgYUmIS7xmWN/CMJFJ+ncL5yazehMUhNlrbNZEBu
nYW8QSJASsQ3QhiEZH6MslW8oFRb1vLxTZPZcVpoOHtVgrjXOZIhXvxuLgZKfKIr
xnIFbWoF2Bm6R3kTSHcT/6l4bYOunIyIqb4c6t6laieqvI8Nuh3fbjW1a2btDjc6
IPAcw4hTHkbsvx9VDf8BOF1DuUJzbVV9KUSaC9YUUjatR+opDrpqzDk2TZvtWiUd
yAwhC76DjkmNE7fGkf36cWBU9SGDhLFK1IcZaCTv7WfJuw51ZZxIJbaPfRNKItPv
izrSXv2xd7u1qnLCSNKbXA1TX3FGI6vNnpfE0ODFs5EeH5kEjGv5AeiY7Nj7+D7l
ahYe3Zl2Kj7kEA1bb4/allVI/ITolmPji6lp2NPqITR+/aZqqHIDLADd1JeCGCek
9lJ5coba6QRiMlV1UuXAmAOoMVSyOwgLpAWVRqNCc7NcIzyCK+Il6lWKPl2sK2Mi
F8+ffAoOsfz3NcOFbLKNrXPRFTb4Qkwfaw5ySsgNGHGMKIkpB0UcC96DYsqRLbvJ
tA4y7Gw1BI4C5zgnoGtXaJlvcysMsZZZptgzIzt7E6wTghQL/Q20ZrDzEkMjfmW/
VErjj1gnaiUnoxpmGXkObopN8MgWkQEvWjlEsbu7pD7CqZTZYTLZyu1KvSDdDp3p
JK96dX0t6LMOBRVUW+9yX7NGJz7MqM62pwPNNs8YETsv8fiaX8e6LdUVeXkB2/fq
hH4GdqlK7Fsxs+vZ+v2sMC7cEhgAANCenMMyaecdOGUab9vm5g04/RJ3hdMwdrcX
NjAxGlthdjMHajKCvVIUbSW54jvO68CI3UMdSrjJZA94yZXDB9bCZ85VFh5hOx6r
EIEZFmTZT99aoZACzprzj8QjZ29ooH+KyLYiqLLEdnGSWycJPYH3Lx6vZZDrYCcW
DjOLLDm5b+29X4ss/yuJLIgLlTmZj5iffdS9B9uqOmuzcK+Cn7fUJF5o1VdEQceE
OekR9HtYwp41zmsoei+kPoI7a2jcoJzpLsgjd5eYXIaP1PLLdf1tO+JqL2bvlVVC
FHF53S89cX5X27THVzxBMYfMOFUUvtqBjuGgrEBoWaK+V39LtHFnI6zENaAYEtYZ
91S70zcJ6ZB0mh4KJF21T0USNkiuEUqHlVEa1QiY2LiS2JQK669F2GZpLXAW/3F+
vha9kc02BOh+KdMoUxKHtXf4ufHiKkrsY+wJlEytSxrYYYcHb2NNMsLhmYp4TgQT
zQmaT7wP9LzfdLsoyTgBdFbhJFhyrnL9d3v0j5cz4oFCL2HTSdb2QmsmEewLjRfW
zOZvQOVoqYrBant0VEw2zcvzgVTOH2T12icKb4NFCzzCw4XtwUJGaJDgmabrB9xC
EWWV//ZXb2jJcLyIJm3O5WwjUhB6rgebmvvDq79blVtGbVXnhA+cpiOfemUX5Qqi
GJqLNMGdny5il+dikPNC8SbDL2Uv6cU3hayerqiKe3N3QB5UZZ2eYMUjAj9T38GL
VinQB4yZ7zeRaMinoAcnwL+3RMwPO7mo0Fg8YhIZ1lPzWqq0wbJAQCd1gICJAjYK
XIE9zKltYgLuGCqLfh8KGEDBYbI+ynNCijBujANWtxnsjK/w1wAatJkyYtW0NZZQ
UWzsZuIXQeTxmZgcED4pOWeAV4PSEb51gnY+1iVmk0mjDb7sctUxDB64AGP96hD7
Z7ZU6Af82b5t8iR+sB4gCNUSo55Y/LQvTxJVF4pv0I0k0Zz9XkBVidfx9/9KiNbq
FDS7pB1SeAa7d6Q/bM9DKHaRlptA7tIUITLQ/Vhbzest3X804r58vrkkvBWRmW27
uS3MsqP7TB2Yn4U95bD+5EnXAizeUYVzCg8pD0KALRX04zKbk1+fn3Ak3a3AJx8v
Xp97jc+Q4WNoDk9OQdRbFwPNqcKqzqZd11in20F8CcEAQ2vp6uoBHBwyS7lggW+p
tibLSYSsBMnUIQ3rX6fTjEhW5yp18/pL9re4++/Oloehvzhhat5cwLexUAryB/CR
8RFv814FKRogynERl8gZ8aKnjr1KMbYWqi0DJvU0ueU2IRy62uVWpPmM0RgyaQgI
3hjqXsUnHROoVQBrRW5PiZ3YUmOQUd0Qm+cdW2MkAsj4ICsCBpiER4OVDzqQ5rZ/
bzp2kHxyN4t76T8F2IviLrH0l+J2TtFbTVlVPuB9VatPRyiJI3vJv29OCAq/9Laa
tnKP9qm84tzTlj0t9JXFCtGDdPGG/9X3w6Pw0UVWwTi122yZXFIl1QkeoUv45lqs
dUp5raPUbqFxA1CaTvM8eUtKBoIta+Hl+6gLxlKcPtmDv9Dc+iaeQslottqlEGU1
qpFJxoanmyJ/NwubfzNcaAnJKPRuET9nZaoyY962fSILLlMumy8U3Z/33eL80tS+
AwzZT2sgxzz9OJChNBm6bwQ4QN1XedrClYMDoRWSZOGXHik+AF9kjXeJd6xQJF+M
T/ITZ4NguOtt+YmXoTVwIjHNk47w4OGVHjFGjOQ96TvZl8YiwdkqAfh0zmsrNdm3
W18/FhnFK9VAaqJAh92aYn9OOBpqYI4lknVrAq85gjE8OO7Z9UFv9ow/z8q6l0Cc
ljt5JoyKBQwvQQq6b5Hayw0xk38dLT3kyOPxoodtGAnJ6ZXAIzvRJGD07ZuWc4Sc
FByHJWueddUs914qJONEElbm4YG42880TVGa8m45Il1HZFzC2vGr4lwdieEjW89w
3ZiXjvZkehKzJiw87EI+zaivuCsi6wDTMVeX52FKeaODfdkGa7jp7K0IeXijOXdQ
wSRfG1OJnTVrQmTVS6ZpV1dFpDsVhm8M6NJG8ikoyXZp0evzgh0RdgU1AmwsLz7A
3onoP8cgkq19iVKJ8IY8SnLkDWAB09pA+6K7ltSaEv0kWEvxP+K/zabaRbyl7HNv
Us/BvSt53b7x16Unpo8wkPe+6c0NZbLidyYXacPhDEJFSnVgIITatmWev7OGNWI3
vYxYqJa8AVVmNgFTgwSTsAuzb5/xZpqv0n2J6yif9jdMb2PLcOo86g6M/jU9Oa5Q
tp2wm3uI+Ph8kwRsb+kkouNS+1fnraQaPsTNA4H9HrBPsmdWz3BMonlz3YnONDPJ
m3opVl0ReQJi6ABlYCCK+NRdfIjlXbuTNmUjzym1lIhQuzMJ9cGIvzoX0R7MQjCr
jZhOHvHHMGLob5+JwUtc9yeTgslJX4Yk/xaut2CCGLW0Y8DoawEIpdvhSiG/TrsQ
zWZmdaW3Lo5Ix1Ko+bbBO2H8LwqtX53+hb8HgGgL0JQiThgQX605EoHKv2QykzP8
V6PH/T8aDSiooA3mQKiAYBUquT6DMknlnRu2iAMFJiIYEzNPvZGYc3vGM3q+rdN1
rG+gCXrOCRUSK2CJBCVJ00ljwWrwDFO3wGACsHS9cEN9tBIljFSNAhcOfx2UcxHq
Vz0eMN7wLsBzCgN/mLkuU4DaGkVABtiIIlUD4LsziYMc78bUJ8jXOLVjho9mzzvG
T0iLk4GZFNzLU13D0ZN/8WaoaYRlpDTqa5RkEbMd0h61Sr9jxJdNNhDtiy+MYP+H
nZIBXoIL0RhmItqAIZ3FGsjWw3z7UVmxyr/Ss5ijiWth3aIPsGCq5n9u33bVvLGE
o0kuTl6boYcAdncEuHIV5g9+G+/ZeqAx7lwMPHYkOfF3SNUu9BLT1twPpNzOmQ23
wUGH4CwKNffzPYNPZnZiUoNq6VHveEV8BnhjJeE+WPSVkxLaHSElLsVog3aAes3L
1CAfpNU7czcJiul2YRYCffTLdNO4u6d3STk9h3H9Y40UlabtkNN2g/0+tTBQnifs
iyGRANQQgcA8IyvRxLF4MS/0IMHdFaYNGkDd5YggEYURKxBCP/cdFWeghlaHKEjF
B3uRdcLFDLQHZ+URa/Lp8mtXBtluaMM3NmAazObTtx28+oJdn0XB30OdYTajO216
fWxW0yNqeQmpwixBABKiPoFUHALLTqmY/4cNVr/RZIbTgG0pPOZ/NF5l3i0cRA9z
fU6q4oVCcr24Hha8VvYwX4d+gqyfeDvz41SLBCSYJnhHq83nfacN92pLO5foZ93h
J9ObyNoBSb6Z5ju1cXYi4b2F2bkLU0yeur3kbsseyKx5fSBM99XAkc8X8gptBFL/
OQ8tA1E/XD7+ZcxHEL2UsZDsguJ5KyCM/DEAwHrG3hC9/6UyeZeWLD4Qe5huhdrS
82Nv/c7Qt6IuVfEjw+Xrv8OjbcoAA3D44wgA/u4fi450cYvuVnm7jzRivk7mQvSy
l1dvJpudY5H7UHOmqwYb/rjDRQlTYouibCSsONS4lrXUpcSLYPHux2I8qdCy8t1U
u2eCoXqEwI/wtd4tvXGZWiDufyI2wXTCUsby9Sen3PdI3Xzgy00lvEtipZ8KJrkj
36lSL5MaUoncGTaz+CY1YThiCOadjHEtS5ifyeZvREFwc7RdIR742+zyJ8oYNdbn
x501eZJ3WIe45Mvbt2zvF/u+2j/VAH7FrY41oh7ohwutUXX2fzdezRG4tzk+bALh
gbyXazjksc633VV7EF1hWTXT04ecRVn8Nj296pvBuqwxaDs6boreuDGJ5DE49vvw
wvQYIoHAtWyU3ZFrFZ+hCRVDXjAeKYnFaeQEg2CXlAqFMEwbKViQXdaIrE2nFwPR
ugGixUioWKOqqQ9J0LARZT7B9tWNV74O3uQGV7CM0lgfRYUr8vzINu/RL/rOHcFo
0+cDfEDNg8eG/8D1svZYYb1JcBmYTFMPHfX1vizNHvSek4DSRoX3GLO247aVugXj
TIarpg6TmfuHkjk8RWpxFFL9Ki4h+PRNBo4m1WO9vWXUgTRG1vhqLw+IDsicM944
eIJNbCS997Hd7/4nkT9GWWtIIntbSS9Q3Nq49bWLEaW34ZD7QH5UwMdn8K4B0Pg2
dUH5gpkMj/5kZUJCZtrk9ST73jL3Fk4Wq2uX4fZrZCCbh0GgK82GE01kq8K8dOlJ
yEJPFEQzyOGw1GBwjo8zHAzk64E7hYC5wQcx5dG49h0lR4SCOsooqfP1QrgA8z3C
sRzPIhQLv7zho6cWuqXULKaueTb9Xn5RuRdvpgY7Ju+jJCzaXv1LjYaYh401nCqe
Bl9xEJZVbC0UK/ae2LZeluGhsij/hc/BZ4LKXU+DchAqnQTX/VqdimmxGFRBScNF
ZX5ykokbsrdEh75LNg268A02IA38SF1FlT8J1OvBRiO6rOdeXTKQck3W0KdO862/
wIM18peQSADTNK2roRj/QAdRTMGYH06/JwZY4ZNXr2Okv+BJMmwpO0sZgmv+r2Bc
1oXqGn2pWJ52/JWyOm69PeLXZiqTwYgn6Qh1aSzxxVbcpMOnh/oWIarnBl4uYmTG
03P17/QZwl3jFl5CXq7XMsk4nPdw2BBlox/s/Kqm5CrHO6lXOMEQ/20vnKyTtRwB
3ulJ0jyHEWff1yBCAJ1+xgpAMaEPHAKCrOmZKFsQkSdwBPrExGOsjU/AsjbklV0P
nuzy0S8zeifFgppjYadcc3ibC93sZz9gAuYu50kwKbgsuZOI49YZFEeobXXny6J5
sqdV83tjTuf1XoGXpxTKytiZe0OOrUJGRAS9cf22CKEWkMX3gnwzAPVU7kyxuCS/
kETs/pK0yXhfiLxuf+sM50GC9VWhvWxvEv8AhngSaPw5i5FI7ESGOHrTlOtuP3Vg
kzX5S1MjK7vYEy1GAOraWRa41ez82gXEOvcl9yjuG1vs6yqkw9I9um9tDWU3iJFk
QE+AKnT8Y/3uTdr0P8oXGZbvMVXBJZzaYMnRQ9ZnXXkvb9XuL7bPWED7Bj0YwcSV
ENYuFppH9S5SFu6ZsCcJhFE6ViVLue2ISRD4dWNlI2EkE6sQVrGWdGxl0c/CRqys
e7x77qFvFK8aja+IrTGwsH+/E1lPvfzce0Z1kWbJkH1el+dkhYwzJPVtaD9cJvl0
3DiWOijA7nYDtzFj+y6l3crhL4/VzXyFXFiALY1f7aqD8QaXF2FYQsw8d6MJCP/q
kaCnkbxnUXbEwvlMl2W5rIDEh7HU1yt/ez9zC74+VV6Mh5Lf/wA/fi9Yshz2FjQ2
lJzs3oBVFZJkh1NRQf8kOkxCxErLRMl6nO9i0PC2n2ds+QegaAEuUofBXVPESbFy
FMmFCIPS5VfoQaZP6xEbz3arg9v/scrS0T+7U3N1f0tn2bqn80Lf6lffi5aZ7976
QFFu9w4drV/oVI2ApPLi0ZKAlNChHbYHgo0gy49GJSvmkTqeLbWmflin4IrgvKKY
r9IoFBUwD4i0eNyqdv+YBogWfYlTTTPuJsUwbHoaVo7cqL4GEU3gmeZBPltKxpl8
wLocJGRUV+GETM0vDFmjrm8UcWmy/wLcZpDFPBan5oyIKnR4UbKZodlgGv6bE/OY
9EAFuNba/KRZDTo722YSV26qioKSXKROtchGKcLywGHzR68wypQ6GPRhPrKADlxc
6z5DElbPRylCL8plDcWqTAMnrPdbmq1oeNjhP25dgXM4uLL3EFOYkvQQwxBjLRgk
9S5+uOchqwrn57LWi/4GbJrOqNhkMJN6fi9GdbTxTRmT9KoyGLNdarYp8qY04ET1
I1cfs7N9vYrgml9cQgfgxbppANrirgTfspfx/uLNKbuffqhLAMCJMNcufQv/ae31
y5/nbKQqa57g18MmrViyjl8cqG0sJRnlSHFGXgfLqdBFyPH9HMp8Lqqdwrki7n3P
7mCrTzWEfeJxCzqK0JC5KVuxZPjmKe/pptIOgxKKEtL55d7ERswyoiPhnUA54u0+
GDB+yHPGJANrTqvtfdm5kkuHvyrhAWHPoYjg9MfVgjBhLoU+mEOg4Y5UUhP+kixA
ImkQmsBQet9k5Yfr/gzByfdoyeLW2BzGA7dqeRIbvK2WHH210JqQmapmr/xG6K3o
6KD8Tvcx8PmwCps+y96EQcELD0NaSGibo2xzZIWjlliIQsUxFPp2kS5ysQZgRd1q
0+x8DiMJgOFDujpsxSGQeQcCRCBEhkd8M25qO4HDpQmkXpbea2KOy4qzTIEiu1Bc
eAby7d1PZdH+IZ1apB0ppy3PHaW0KLKBCSUq4R+KJmUv1MmUeuuu7eBozRWMVdKc
ZmXELN0eI6EB2be1ngSJDwzvGSplphDvAUjOerSMcBTd9iMH2AMqbwgJ0TAkry/W
khSXtwrL/k4BtnCrDgf/lAN1/knVSnu6mBj+qX79BZWkn/aRsKDniPfW4Vp0Rcy6
FFF0O93s7HUkTI63NKzkTCPdD5AtcOH9ybN9AwG5oNLqK+p2E2Cq6ImAZR55ckuB
50mzknlP6D+jPJ0rNVnGcrOxJRWLayZCz6cnC5nHrR9KFuccAgYxYmZEAkRVJPFA
OV7fuiXZz17QdT+B7KpTyY7PD0yp6cBZYPtdxl7W8Nxn0ApNZpOrwXAnwusSBGWk
rVL2qI6PfO5BWV3JRlxOxOTzvHyL4vOEW1F/Br4a/G5uOeNo4DLZarkYvKsjRXWn
7XlF+xbATWg+XEtfEMTKGLaDSb8iZa6MA/rqBx7gxFgs3g/OjbbSvVJgkR5bJJUn
gsQqFvLUK7x/tJLP/RockXhpFNHyloMvFNkot0CDkAMsz8kMHLpQcYiUXCp0JGjE
sgp5W09kez9HiR4jhSCIu7W/uGT9iBsUE/7bKb7mwYwFcdLxZ2E/k7qlorIXSDNo
Xcxu/yllgm0lxfMJZ+iDs3kIh+gUqXkS/e43VoXKX2pNj36d62YFEfeRpFQ4kvoQ
ivD4I5pDbO3IvdchKS22jx7zj2V/rXZ+ZQ4sMkEWABTKKvxhTDOHyaKL2UCQx2Dv
hlDO0rzVmMACx6Qnhq01Pb4zmVxQlYuFUKLCUydS+tFRoKAKA2zN2K5qyIga+P1X
fCqcUz3FCVX8chwh3sQIjjOMPHjkYYPw2tqyuJcP3isNM1PG8CRZ+vBZeKOFwEt/
4AkfmzyCRT2WywUXb2bThL74IYoH6Nudth2UDDdY+r4ZM2HH118hj/pwf0S+4kVb
1DjuZOAvGK7gi1uBJs4b+2D60/kDKuh7xsaGBP8/M9jb90dOBFCe468pF5eL7h3y
6wDkPFuqzoay0qvDQrXJguwLy63JL8VSR5yJuMmvDUMR7pzw4bPsfRMTXvB9dMg9
1n8fdSUVKL2E6HR46YlwNofd6GmAIjtBsHqE35ISvL3eJ/kgs5rqoMXqMywQ9GtW
jha4PRWQzuTH9wQDRMoBPNGrtvl+0oFJScNTpWnG45mA6oiwqlGrmQsbTV/dEGFP
xb8MnQZJHg9bmX41GqdBoo8ZdpeiKC0qMmz6MnuloAYnbAuKzbp65vKFBu1x32BB
lGCFfLXAg/xFLsOPUh5Kc1Lh/VHKFLCyMWpGhg6J94hDd6iPK6k/C9hu31GLdp0u
Qt9pggUxcPScxZzPaZhbLoeL0d+njczQ3RaR0VZoSDE5W3dRDwG/kaVW8pdSls5q
aTFERLH3hkmWJC8rcwPej9eNT6DwfiIGTF7sPlkTzt+/sGVu+f92sHcEqYApdGcT
dfSx/iLNn8fe6OLqBeyq+8oeYxCa6ghj28qgKtFHRyDaLegB6V4EEZEDWULJUe6R
c0wns2gOR95MkMa+CMwu9dXRBebfnTQkkrteIXP/NJzhsZRMj6cHSEcjxI1Z2240
ffn5FRQI6zCrRlOR+Fhf6wBNoZeaqDyuf8vUZ3/ANtsIipft45JsJgY5AGRc1JJb
g8RAod2PnnRft6Qv0qohjcHAZ5RTkf2C+0oQAnm871d6Xo8AoCjPGFUiooakHsFU
S9DgCHAvAV6vQxeoMKnpWkRN7cBGooLtVCkCSEF1Cb9deS9a1kVTmoLCQVLWJzKO
QoPh8E7rrstCcinOJFSz3VWFD/PmHTZzS8bTei5Wka/GD7dbKCr9WXwJ2iwMnu8m
fFPohFJ8cB+0uzpJIR3fPl3pM87vubTQ5hz6hV7jpTsW5BTPjjGe0nM9XzjtkUcM
MLgWhgbEzmARjMwBVmokKUbh0zgbQzdgpE2lirfn3Ol1qHXebnUi+cUIsLJjepuV
SCl+LrCgpCGzBt0cElufnPQALG/jRn3dg4JT5HxfDBor/szqgR22y3B+UROMSYcw
luziJgdJu6Y5iVFYEl2cpoLIsmSQBGV4WmBlsu+6CIJiAwniZ807WjH2i2HL59sN
YMalz4+T/a2xYLHnUmDB6Y8h1pANlPC2tcF4OjuNQkWhA5o28zWxTNx41RoniBA1
9N7Uq6qTKAlPdrE8Zqxpjl725noIvlxtQeeRwJGXjAbkomRf7trT0p+vtryfzPx4
O95QfXkDPl1Pl8n/dgGpsfsEZ6Y7zdd5INFlvPdavICWgKsz5S9mL9sFZUeDbZ2p
zfF8OHoCjmLjvqmoqOyoMpCvW/m80jszV8Oe3BCn4Qi8Rmh1kwRBN8EaWetEVbnT
fWZrLpA/+4VkiwkKB51GysFL9w9oGiyM+6g8qUtWOZXOAL/Xz6/73ZHVi8WtPoRr
lvbNtE0WcqpQvP1cB2kfKsn0UCu22itrwyGw4S5ujWGqI8IV/ppjpMdqB2bGQ5mt
quI++YQgQo3GUKOqGE1UhvKbwkEJRtOKv6dzBefRaPF6ZrJlb0ctWsrcsOsAWHr+
6oN4rPMJ2RefQVD6CV0LTw4wMcvyBJYRcoXyiUdLc4lE6OAwTEJ0RBOs6/iblTCp
tZoiDyCWeC/N1cz+ztsJA/zWdj6+CZ94TpnCyOSn8j1q1QJAYUthUhKJEN/B7URb
9MfLzTBPcnjnONouKf0YAP/HQE14IXb/AbfZ9JV+LeLhEHXBhlyRvVw+HKmoaxC/
e7IHa3Vblpm2tp3R67AwmZdFXNHAiER+ulLGd3VgbqINgaxWoIDPve0WmUemmkdc
eUr37fbmESsmv9Pv9fRpe5TPZlB6ZNRj3b+pICElIy4hIQ0ycOp7fRNrKsWrVP5A
DORq5jNZh8gi/iGbKOZJo+t2em7NZti0JJCOLlouGJopw2f4fsBvFTjkRNmfsywz
9VeancrfzsynhONcjcDiz0fy0oATi75QlUwoJNFvYPXxvTpha6LZQu91h9u5kMb2
g3MBfP6JxbPKoXQiNYkcZ9TIrE5Fg3zC6xaSj575Er7PjEM31ifAw20nfYj9iXfY
lGYskkWTp7Dzsk+xy0d/iTyOmtzh8zGA2Lm1XJZT0aHW0HMebTFom8ZDLpMDX6Tu
m430bABtM+/8BWzS3pryJJs9cPm9a7GfyZCzWxpsQLNXS2AIIFI3NqOkU4/48egc
CY9eFHK3NOrDLlDQ5eORT8IrkHpQQra7zyWitmCembsW2RDESOHwMY3yuNI4XVB3
ICNB0eElMhEWeYIr4X4C5uPW4F2qUYydSVmP2LNmqe6ihmHuwRChks2uqPstRuTq
VQcWnxeAraLPb3tvEFAux2hdyPxZ6TTCKBP63d5E2DF+upSritwY4F0K2I2yYA3I
V9AgVs11HyKEJR3SGJEFEF471apZ7/+1SrsqHBgk7E9rQ17JYOsMYHRMnctI4/x1
aw12Rb/AN6xReL3MUYstCY/ouC1GI9M/uKAKzkcn+3WpUAbB0S3Yy4UfcyVc83Cp
qsUgkXPjS+RQsnJtua17fafgtr/5mxm4kJ0Xxu7ElpSjEkuQQMh4lqIVHpFWJ2C1
0XTIbiBt6whtBhxlRWRhOz8AdAQAR+vTOMX4BFuQDqQEGo07ExMQje/S8W2CMf7F
1IJ2c98Cr1xCgiqLv1uEzbC7f3mmgle2sXLxM/bIX8oNZBULO0fPXFVyyqD9DmhT
7/VJQ0Dx6rX2FkerJwTuTJrLPRccRPd0pM2R/3rztfMbW7iNP04JZ0ZALgbfeAsl
1wk8VM9Svo3Eg/091HLtUNmRor0e+HzAW8d6uttQw8SZ0V/22SNri+gFCzrSxf7j
PvhMH78XFKUVQE+dNsxSRtG+scQxNG7xY2MMwyu9zQxC0Y6K2Slu9EBi/Huto4Ur
6HLAiD/OjiLRNkGnSb9/vIVejnSXrKEHrjNoFrPOwBArf1rf6/O6HCE+hnfLM0N4
h2y8761dmZxaOmp90//f3Esy/SAxRSscHSyJsTy7Ed6E2X2RAmIHZ6/TLOyQ8wn4
oShGzY0n6rKWHrOBgYCVx3mnwGqB3N7JVPM6bdHul/TAzYd4J1h/j336z3MOGhyu
S2ZiMJzNsLr0q+a9o9H83zdRx54Ziqae1c7nIpHwteeON3BMddL6rKXHtLx3YxuL
nzwMealIVz9g1EYARp6CTDzkOIUydtrptDyKDwsxutvkv7JnnPeuQst1b8yw2oox
UefsDLyt2fwf06yeRcLzsIXe6/gL3y0h9OxbvKtV/+qvHHbZPrsNMnmXNHIx+L/9
GvUwT5kfnPaYwdpg8B1w4cgZnIAxXAiGr8l3wLKW/r/ULS3Px5Uf4buze5zhqNKb
N7JN9L3m+VoDBMZ3AbqSJvDeoWl/ouE2sbBiw+4ZQDqksIdayZ7kAX8EVCCkd0jc
eJZ5ijKRw8cu6MVfHroeYvK5PeGskrvCJQbszmPIzT5H6kFkPAksyTyZiAvkKXIn
32a3Wk+gR+ZaUh3zwSzm6qukOPF6HY8gOgW4b8QltohuqvrmomP7g7PkuidZZe8h
iMl7JEFwtjx5mp6N12fKfD47EA9eh/+r6Esb4+5oFeYwX6kSU23unqlpm8b3TZ6+
HHUctS8sieA4rmiXOpiH3EGWsgZ5qfeiyheKEhbpIuDDqclFBlZudojfSBQBZnEz
j4ZdrNcwVcO79Wz5MMnWXYVGKWVCe4d1RQjsvTwdm2sqp6tFhH338IlpfanN0ec6
+CxzT5W7JwA1HUHZ+ZzVhI1QJBDBPAZEFiD13ucmLqoge0Em4ASlIJ7RRFhu5L5z
KL/3buVqUWkGolSjNTRT9YGLWt0GjpiEHPrKpnAUlJE+daXBe1jfhdDKIQo7zJQc
3/Np5YuWIfXyqWZMYWLpp9rIfZ5+83GrAppYSiiw/Se9GYMZwd2jR3qoj5mfHyXg
OGw+pJAC28THgJrItTox+4aSCDYDsMF6ephRaFAYICpDRCivuM8/I/yi2bwW03V0
mfRN5led9hScaCL8Qd0EMSoWkvsfdzVpiIu6DI8A9oy52GL5o8mjZrH5EU1tEfZs
n3xZpNGHLWSYTaTa5/8nCywxcgiVHozCA0zsCRJCTf6ylTKG2MDEJiGEiOMeZGgg
ToRP8lkfMzm+tG138IFgSIOwpjdjFCBi6ECNiSvFnyZqp9PmxfTxhUD4P1do0YOw
iq8XJBrqKYbBFigKTrxWKuSp9t/CQzlxrLNHRTuF6QjYTgmO6NnRgkIxMGw/mFOl
FsXusGbfzCRBW00/79aITQ3uagF65urCC6fgjHHSyTpI0b+kIc9Xf5Fd5Nm7Qb7J
iURf0/N7JX8tRt0LnT7FZ3K3F+rV8FbFUsrSU64x2QjDO6xhmC2nJQuOHFh7A4bi
RfxYG4hV+ur1cDEi6LceXicy3aUI1COf+oKPk2Te0Srbpj9k6tbD1ljrvOwStOvo
MiaYTdj6hfNFKri4hnxsPYZ7V+9PGTQ85Crq2Lf3iujb6000W2XXPhjv5fKgYYzx
n1oJ7gNAlWinKbaPa8imP2ONIQWylXVCurnUoP3L3sgIlC1TVBNBUSAnR2tWFB6r
grrGON+YqFTETTJ53fvOQLZIek/BsU+0UT7V72WY/DP3GV11HOpClI5aLL+1rzMm
xILXKVqZuA6AyEob5hk6MBkyGFEN7Q2QNtQQZHACjX0XkvxwPvZ9b1zJnGbPtsFP
uUVWvV/hfnP78c6sMj0VM1jR1/VuI0JKqqfodzCudOiMDtnhF3COIfJHcBrzt/64
hx9bkLZdcp2npndnCOThvBPKGVI+5fPshFHsVsK7ldlyLip+czR4/oN7jr70psZC
FIwP2UgVQLYNHFca26iaP5XUj3s7vGJUdJZr0dWk4aiwfIBelQAWT6WDjar1ReEI
++9qbll+idixrf8TapaT+DJtNqrgtS5qxZcPNue6yYh16o1x7LwiyguDoF5ZUXHi
G+styvVxL0LWEsBmNX3ksxwXfCqKIGJvOIFvAyoZ9x/6lghH1OWrKTlD3VqhZARW
EyQwQ0qnz80uEHfaZMPArr0S+GZMZwvgITWMT+ZlVz0Y4XuUK7ELauCcqSvS8aBw
olLw/zk0NPazpugIEShjbLWMXFScOOG4zkWaxg1EKQv3zNfwwL9UybQz9d0jW51X
R+JdL5eTe400/ch2W6kPeKa+ex5l/3NuDq95QyCaRvUJg4UOX9EBB3y+sXryFKBu
aGADTZ6PX8MvWZSlI3DcBma6yDCd/fVfiTOa02NZ5iivb17NPoXvGtNxFnER2MZT
j1crcthgWfi4nEy2GNztNpUJriRFiW26E3t1ty3+lQ9qQqF6YHa27fd4zOu5qOZg
LiS7bkJsuElxis3rjHyyOTB35tDZClsIl0qi0O+dGJvyTFsfzYFanYt4hXfoG3SE
ZRk6lR4pnqjXm1AljYcwUJO2ySybY+KWT0yyzko5wKFa83oby3l32KwU45j1WEtl
jCnzvTPwP7THV5sJ5BE8KNxjRX504LmJDJnc/S2reqTgnNwyLCyDB6JOHx6RByQd
WOZ5bM4u+caC/AYsq6CdmuwP8wAT9C+QcxKqbKR+w+3A3Wn2/1CSBAlShQ8OcnCk
2JRs3IrQENUjMxaAcx3NuNrBBl6ys3440Rc6Ba60+TGFLweXTRIETRM/xYTgAEuh
eMRlmBMj8P9h7kNxgg7DVYCqWwu7sU5J8ltcdaenbodhwCjj+VQ84BKEB3zbkEK6
pUmVbHrL9m5a7Kkd9jYeXR1/GJ0min0KQpuKl0VfW/0fak4V9eFzfX6VxSm8hf7/
OCo71hVcZk0+1Ra19l3npb75nC9TOkEc0VJB70E4S4pSNoukSI5fXWMRbWDqh6h+
SM0qda82KZ2Gucwkj/BkVNLKWBnWM3cRjlgBdWQnuzeORxuqlyHBebyMdiDdLzYP
Xs+efavWvGVAHeEjYUwRSX4zeJA64S6RoQvagL6UtGDKYw0yKFJsyQTKcCFXFsVg
qpVDSsykU/ejrzmc+Iz0d0jf8sgH2hpVkLN1YE2SygTHN4jlS2sylCSw0yu7U6Iy
vP1vkSolCSKvMbr2jMBfxkY01vjHtitHoyBcHvDjtxxfaUB5tSysp/pdz/w3he31
yy/vNRaclBi8SC/J/j2tPVQVUHI1Ebr95xl3AEjWI+6y9/aZkBEzouWUVGNqT77y
yPV0H8Gk2Sg45m3obvwzoe1mT4nUeoiGJq/BBpLz4swLWjI2XjBUAi8o25yqbo3L
L/BDZTFz+PtomyaqgDaj2q0xA9z9I2aX9GEXDQDh0S+hkA0AP7/0OTcNLIJw77Tl
uh82IjeyqkI89EmOq2CCFP9yLqk/qoPhnNi0WCLcZzw9dF9wk7WgizlfrvQsGAL4
GH3f3gcBf8Ir64VovsCpcvdS4IXosUU0L3OoK1wKCgoGXibaZ+cM4reoz4hFubfr
3iszcBaAYQAVxGDewOgpwk9LGn/nVA4t8TVwFlvufknNhKdG5mggOgfxveq7BseN
Clws6u/yBtyMfV9/D2zRJMKY8DUmyMvfiHiF64NfRO2oWjSpheIazzYVJntEipoT
WPFrE7bkjlTBctQy1DDdjH7C85DTOtRCMzPI/CpQexXuMoLm+kpXlQ4DolI5tihx
GW+qaoX9tyToVP5E4P9Al5c9JAlqHqUaF7m6l1DsaMKPOVY+EBUOP+tkk1SAye9X
K4VWG34Bx7XZRLUQJKlByEs1oKpjlvbJIJK9IBB+AzkfblZ1EDWcKv/MSPqouaNE
c7AL38w3knK2SC7h7ZnRa5cebohOgO7QpuiDbHEfiazxTt2NUaJ+/2PmvxY2Cdrm
tryDyn/4iotnCURPEK79A4ReFvDmbT4LM+JVB1DPmrhSYjQzJnH9aTIRms3gIeXU
VJt/ffRgUG8GNaNtpcEBhD0ILBnB0A/GioS8C6OTuiVTGZw4NTXoA7nh9tO7WpT6
07QlgnGCyZhtxRUawoDbrbNkXl9cFQQFWeJRp21z18Q38RdgVyd95ns/dbyiLStS
CzV2OLiianoDhV01cI0M9rbKLk6VDqbFHPumGBpwlnHLe2mrvXj+XyIg9cV8Bsct
eAdBV4meIwjqxE38GShPiZ8FztzxXsuiYV9ILK3777EGDy3A1kFwBA3mxx/xFuwK
zRlYsCzAToSqvCUEXPuzHkyp0Jzm+miPoy5h6JiBtvUDMJWUxoS+/2u74BbVtWdQ
5rtMZDJwuuN2ShWCwtCUmd12z0oXj/MCcdiKui1+A92lvDaUOAdwC9V5taaMr9zJ
z8HWddw0I0uPTIG7YR2zrM0r7B5HhRAqT0499pjPlHeyYgKqcctmRnKC9P/WWVGL
MYxG4PoR0STdNAbLZoTGAEXpxwIFn2VE0AZ/5KrCHZb4d49vx85sasO4jtuMNlSw
PdT/7IHwTEyNPLtv3i4w2fZAqotlOadzFfUUSkIR9hu62yeW6cQWtWUe7Mfm4S+Z
nMgOkPsOEpdCDB8r0LBvSjlrS4sXd0xVK0ED+X2TuM5NR1X47hnP8N8mCr3YBz3F
WDne21xVoCCtVacz7YYISKhx+n/VT3bZygfpgMpoWHjhfwdUVKrMW/LpPoAhWz+N
viMIUoQeG2/QWs7dVVHRzT3AYqJPOaolQewa/6ohIcQkuuASSSIo9naVsudsJl4+
Z11spOVlAxbk0+zNsxWMCNIRYulA0QGpgpc2pqiUSInstAOp8iz9Hz6EI9ao0hTX
TS/cpIjluwyR5+KwrG5yUFwZJDd6Dvp7+N4CRG2KMlAg/4BMIDxbn5qd6n8rqS2T
iSezqeplsZDnlnA0KLl24tve0K7V6kGNS6ZH0cVaaI2eJFF5PaTNC3r+GstpKTbI
K25yhrJ/w5AtBq9qZQMUOB78bBywGSj7IvP03jf3c0GY5PW9rGgHrYzL8y9m/DN0
gwZBZFIYyVcVjhHXXHLEXcH9+lIF2G75IUekm00n2ZjhYqEAf2j1qZfVRGj7vsVM
4Bb/28MGbK7ubIRf/2FUadDa5TyiF4T7UFIGrsO0USSb/RVQSQToyJRqwyEeTdPH
k+3danBVxSQhiVxwcc0kTdvSmtLghkAVJMUjrkAk5S9o1iWrFauBKfE6dBJg+3bg
qn8h571o/OdVL+D1YnAZHnxFhKYseExN4YZhHzdelRPXEiEBnw8pizFEkxRE/R/t
P/A0unLU96ZFvxQn3sqZZ35yA5PtG2sLi+q46th/WQ18Umpy9hXE7dFV6KsmSpGi
GzJ15XwQ8aGuFhVpb7hu7O2NajoyuoE2s9HUNhv/tvLuxx3++fEvbVdFTfbM7X1g
AHCAWk3D4hGU7pgFKJukgjg5i01V3pQV41RDBe/urE08W4w5WL6MOgvybXjnTEzx
8hOAzmdfLp0w9f64WjdjYB5iTCnRMkv9ybZ596wn2w2nRsK7k9k6HQpdkRnnCrL5
Ij75W3sUxhKzQ4t2DUlS1pZMH9KWnFB74S8CbVNMfpNvE9w4LsMFBbaBDuICY1zc
qmrT1Y83FoATiLf6XvWeHFRfNHnZWBSzOPObvxp9rFl5HfeO/LjfLyYhcCJRt8jF
OD9sEARI6/Xhvniav6d1Duonv+yUziYY8NHJ306uWSNYQ9TMXWRKcLqwyGYpaYDq
TDUbYL6lbumxvXppPsFh4CpypEqx6P5pyQ+RPy6ER3wpwz9L+hdBqizlTCrfQ+lL
CB90eCTSbkmFpDNSpJfTaAmew+7SzedVjpHuM/CsFW4catTrYBRlMi5A9MeDHxPe
brB+bDtXiAtFKEoynM51vOKGCaHezzpXYf6JOf7No3ZxynjFcEoJ/twyyU6f7D9M
kqaTolCIk01H3QFepAKSxpyrSh6qcFaBAxa6w+nlTvnshuil8P5KvaLwJW8Z3Tq3
sHAWEL/nRr691FQHNE4p1jZXM29wT6GC+XiQfDSqDRWs7WGdAwdLLp2l/7u4kt/e
TEHXlcx3jJjMbIqC5NSG0wcvFk/KJTj93RlrfMzvJAE3nulqkb+5Gb5PNKUmQLFA
yY1wG1jGCvORtZOaSlGItUTMjdUJkNlCH6WxMunJBopiTA+I3Yn5lZf90OhJjH07
xjougYWTEkwjbkX5b6Z1QDDtMo9ldhk+vwFpE1cKt+3i2Kv0SsBB0FWyTZQueq30
AMRC4WDBCgZr0WR/bNN6R/qAiq8RhBcf0i4elFTqWpjgL+5Iwi7Bdw80AKHW3Ka/
Y/doAopgboDuNmgXu98jvZVY8w7rOsd0J9+Py7tpNgLukdwtzl7LAOlHI400YUG4
1Q4vW9qYeU63jNRTPgrvk1pVSbPT6cx/0iS+j/3daTjclvhjUApw1vQnoARBc6f+
9ZbTiJYUnt4E3iIJF7cgQTQADZ7p7BbJS6xIYz731L6+C5EX84O2BxDD8n+nEJx9
qzESfRKfLgdb8VZILJbVIgkSLq/tlsJqUOU2xLEyoulnFHQR+dNjkiibh/SyZt+F
58nbN9cY7Cg9Lq+sLJsXiRQm+BWNJRJ2gdOfNWbccMDduIxnZyCZl1q2uJy3qX5N
/cNZ7okWPmXg2aVgIhevFJtum6scBfXXffYpGI7z0iYKhBSEnWB53YyqodgJRDeO
S2Ydy05zKefRJOWkJOdKZXyB1HIt/EN4d0p8rAZU9Lvek5QjzH7dDnNVi1DsX+NC
CN319Y5k8jdQW1FUWkyZ2R72lo9NKIpbC8kBaZhaWVm3yr9J8bAO8VOE0tQx+a4b
TAF8X1N8Gqclh8gyRgiInriCXFzFP/eGNrPPlG+AV/LnQ34Ia99lGbEE219GQkWJ
nXrrhaGPgSrK1/kmwrQAueOPQ6CCgqMi9TGUHonvRdc=
`protect END_PROTECTED
