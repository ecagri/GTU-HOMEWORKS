`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xIjTYUiXSoMJsqWy2dra4fBl5HMQYvI/dH+5D2mzxOmFWVqBDKY4mVTY/Gu9s+tE
5R/3qwlm7ivjcCw9h7S5ZLTV54nZ1b8srcS0WCbfgrpsJQdHopgjItEsjGDUojsv
VPn6ExdjpvaCouJ8ARs1SUo7P7ROaekG1KfGKa8EW9U7ImFk2JuKLPGJY71dNuwO
tF45x4Cj/dGtd74K1IuLlt3KjBa1NAdrNsw3H7YiiObhh5eoPg67gae275zyOXrH
uzTqA0Fj+3YYRc5diyOdJnxptYmwZg5aWokilam9SfmdAWRZmABt3IHOmPgSkLum
K3e+QHWsOGyVBR39mB6NKgWUA58/5GjW3VJ1Hquq9fEZiDNwSD8Fvik8YQ7tOvkq
vCV4FzmcKBRMq5FA1KxzYUCmyFJAr9wIpIeRaYp2w7UFJ85NoqGAnmu4IuV2HepB
upDuBNrw+tA6jOSxBMvWQ8B0OsgnimNM/zpTkd5o7Q79WsmaDtEva7W74lU0/uiz
lcAjvU8EPys/JN8bL8lXhED5yseZvPUOfY9cJ3RCPUCVaR0HS8I0Nc72f7q5xLL+
Dq+1TZG2/YVsStqU3oxhtwAg0bX0lXtI+vyhYR/n0RrvPNM6nlCLzA4OFPmfOXkT
m9YTGTsu36lmCquE1r5ahh9eHgVchueGkpvwW3aczK6Ll32iYSYeflQcGf3LGPTj
6GKY4KF3budkv4Nx3r4KYzPNlWecHKLPOy+LlWVX+0byzs1KaDomTyp07zGVyVSq
hCGRQSByl/cYhA4n1WVOXMy3nam9v4sGMlF2UQwt5CF1RQYP14TgdJjlQUYawe4l
6XbyUg0f7y3ajYab3hi/swp8eWLsOkm5676PY1HM022hzZNAny75JvNoyqCpF0Gg
517d0eTDkG3EINNpJtEqzS1tGvClXNjBDrWJaezr5SfTcVggAXECqeQfhpfakKUb
N8ToMk3eqGKI8bFbMLnMcQpryx0zbGb7TipqqQQJuVEN2D6g8ITUpLbdBhfQSZtj
EvFlc1N6YKDjFu2VPh0WhBO6T1rgIO1kwASxQtz3wuxABHloZJSpZxK9HgpMKKz9
PRn9f26fX9k4VuRaYBA2YKmiQZDWBBWHfw7jAFZTQ/Cj9BgQ4FvqpX3zPOZjtYkG
QYtnG+x06zr3RwHu1OrU7Z/SMOos2ELw+vwOworLEwStiuojIfSLUlWvvKlWqZW0
`protect END_PROTECTED
