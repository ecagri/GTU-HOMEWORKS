`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0bTTAZkK8CGxe3FTCMnSIb2rrql+5u8s4leLc9MTmIltmqdhuM7egsgrznJGagfJ
yNeIycTavRAKAzl52C01RfsDEDc2zpJifrbABHJmkYgFMTEovU5RlKrRJUrP8whe
4eiIHc9WIr0Z2oc0gQVYx1svB3SMhbK/9xsJPOpSOPoutfMQiLqPwpyc687/S1Bs
4kBS1eLGFvPU+xsFPK+yarwZtFpCTw1qu1oG3PZOAUsV1DuvS7MZCjwE2K3m8ka/
1H1euHHf207IVAecVM3U2OPU7RXV0egCLQNNgKeV22zb7dfN0ePOG4793ZdySwjM
2BZbW4USD15vtLExAXdkupNoVmMfVH34h30tUGHalrbLqSnjXPh/UUQVGZtUrXMP
fDKjQXjDs3iBhy7FrkS8DMqvXEHsWC/iD83eOcPXxg6Vz8umanG7i2u/UH5Ak7Ai
R1/gvkrFHRjc7ZthRC/UCxgAp3zxLhX/n4wiml6RhJKD8a9JzxdUEyWGe9GV+SaH
yrKlTSH97zcVjELuSEphhzvMS5zoG26CgcEamUogsRy5uvugGt5FeUH2lNIt65b4
fTaGNLXlAvKwDTYVpDGUVkHnVPVmMAi9OIdxN9i/nRznyEIVsEd06nEJMcggYwkF
LFRGP5co3CimaeOT+Bw9XqAUalbw4jXiNDy89DcR95qpcTHtrbA//SYLy0Z/XCTO
YI3rwr5xqkJICesKz2zUZ0hNheER5nnJhQLlt0OfqJ0Ey6cq8Olmfh9cJSf9f+Q/
WX394dK4Eprxp+saFJqAduf/s021WGfoANsYL0lj16In1rMJ58s/Jc0jNH9F2+j/
ZA9oEjVXROHeSfxK8rQ+PWbZnHd3A+eQYBEb31+JX7Xm4CvBQ3O8FY4GIOyojV0K
h8zlLzobTu7ZTfOgCCTaD9ra/h7Cdvs0I4J+Qnf+3bM=
`protect END_PROTECTED
