`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YzVFUwS6HsPTHPHHjtylS6gacIQ+9J9tXEWu72YuIOSbjxM6AdlEuGFU0+lvFCRZ
SgsFMPtaMAE+D+fB8NV56Nxd6Nm6KFAMPspcnfO0kKCeORwQI7At5qCdFouSZ5pP
KpAHUKP8OxVp+pQIIT4VKyuWsriCujkJy7Fb77MPw2rK7HHtUheDwgQt35gzSAbS
KNq4q3R7b4+0CsO2aMqvt4ibz2Le2ShysBO4NkbyOqNPMGgCDYMA0uK1UCDQq3GD
971OvPsGIhxrUuBAl7X6tHWLCotlEigIcYKwuG6+0Gj9MseYuG4XkugJr5pvkX7g
CggCGbtb8qyR97XTL8ha+rYFGLF+Xn08CeA6aCi2XGu8WQ0Ryy+AwtjT81Z7KkZ7
JPJIVrvBmW7ozVjPZFJIP7NpAtS80dYYPtP1Fcad2tt0NpkwlJQZRaQBxrLlu4VH
a21NtqRx3Sc1Xih+XoweSCQNdbgzy8WyvtdI8rixuGAusw/a865m30nKIZT/vF2z
iWxZ4C9j2o0X70BSiw0G0fTwmIFtWGQW2vSI+heobJVCDz3dFXOx4azfr9UlyURa
RToDB14KxHwftGrzvGS6jQ==
`protect END_PROTECTED
