`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DXNzZZ88+LwSE+TRNQX4THpScRvCSys0bS0NpbpVxnNdzhTeqtqzP8W8l7Zbq2Wm
JQ1mIFxPgG6aQlr8CZC+8SQPuj9QYAIGJv0NxR27mxNLTiYNOCbmnS9b5uOhjch9
BnVNKnEmvXi0FFAq0uhN1hjxg1djNj7PIb144Zh0UD3HwkpWwf9Xw0USd/lObmSl
j9DmZ1sVUoXR1lEGD984gc7DPj2mwwHIX6lmTL1IyX2H/hNr+k6QWb6oR7aJosip
/psoydUaJp5Jc0Ik0niX//ohEJclyfItiJJSnp//mJF7e5E+nN+HatfZT0fBCv6k
K9IvHb6qke7mxvkuLqtGP2M/dGeuevQkxh426r5xsAaA/iOX6KfVgX9WIeM8YAF+
b/qs57jLELeSNHp7jvQiPGbSpqwqad6R/7rpzmNuzci3Dng53xTYYBXMHIvweP7v
krHSUcvB23BhVkrSC+X7pKnUGOR4Mb/SjdwC9m015XiwEiAU+RX9LYF6kSwuDX6Z
KEH//bmNZfkP/ZBYez7rqEP8YJqP8OAfoKd62YB3KB8IR9T/dVQU1f5W0/NC90r7
ddv8J7lXevDSBTSU6ogxbyuqZKSacZpiSrASj3eLG80oXgECc7CeEoqPwM+iAIVM
+U/R3vu8Sy8yQYIcmgryG3tr939UX8sFN6mjoYzA9jB+MuEAsPZ7uzw2yosWsS+G
EvBt2COZue+dq2g6G6izx9M44+f/d39I54ZtDPEIAUeNnVC33HLkRUoAEeOsvzPI
ldJnCRqrJsF2xB9PFGHTTzuNIa/TthXudPSTbf+D/Oh4diiXCV0F+Sgv9Ob+2sof
ElUxiyDtrZTdJWtxg7wGWnUoPY8DEEG1X+G841UCFAT1Ng8XMzJz4sMK8gW3Jl1i
v5WXZnYDet3x71n0FztTmA==
`protect END_PROTECTED
