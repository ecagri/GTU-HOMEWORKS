`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JI6pOt410XbFWEw4/zzJ7dl7p2aNoI/jFVe1Z2IvhuIguAHI9um0Ep5At3KYZ+QZ
yysIklSlVW2SnrBCtVhAIoFX61clUHGtJv8oR3f2tUcLgPEjQJYFS8Np8TlcpWpl
l7Ct91bh+tfIBLeCsh9Ns9FNfmCZ2iT181oQ2C4PdqpC9zsQhowXuBk2YZZ0REYZ
q+X+WG1IoezFmHAUCEe/nNf1Dt1vYdUjkF0WoXbet5uSRikpo4J9Pljs11XAjm6V
DvIddOhqa0C7Jfj9J/Stx9lUenTuNZQ8/F/ifvSjzfcicU1ic/PCwGSLXeTFflc9
pzzRzCjS3l/6KA5JbdglwNuqHoBbIVuVox0iU3FaTAug7h0YxgJTFMZEyikYP0ba
q5GOZVg6jepUJPJH0KP1v0fAtX3ecWU689zhpsWCuGeEhFY2pa9urTGbD5Aa/v9m
/mTSEj+kx5/IKw1HTyqsj16DGoAwFj70vclM5xht1B349xg9EfF3OVGz8PW6QqQC
4r2wSTBld280T7OzNOR3hRLpJI/ECKJkwWvE4ZD3xvQ0GbA8WRi7QXrwI0JyTdiE
fRaWRlYVo/gvZEHMIaceXheShmrXvKizhSTPSfs6ANUY+ShLC8xsmgjlL7YK364I
RMdcHdNAIPjR6bcyO4TGfILiFvykKHyLA6kRJ3McGM8=
`protect END_PROTECTED
