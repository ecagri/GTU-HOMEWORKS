`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8X4HJ8EVLZdnPPSIXNY9AKDwnhjCCskUD/FrKas0hdks1GaBofdnNUCCIHBxlJ/X
NL4jsP7sX9vx3CsXKKh++3vITue5Jo69QYMYH1qnH+J2iRWSYutaxolqS97w7b7O
X0OtZX9mBEhiXUfHthcmWEhIX88P/Ocdfdy6JPwY6ngec3o6HG4poN9yjnwqZLZ9
hIKoVSFBbQNBaX4j+9LFRDQ7QG90o5HLU64yF2Ka9egs+BIfxVYDY4VSFjN3SnT3
bLui/kf/9t0cZZo6peJI5LUNXRf29jWJdeMOwl6JtsuvyDqrI4AntugBMotoL4si
bw1qV7LpqHYrKYL4hdxZ2kEZgWpdU+lYDWtzztmANVUPVNTByiSvHScLSoA+rCIc
iKOfmBCF3Zh4Sm8X5mJ96HKASa+6piiATOjy4dWtxwVzOmvo6My/f4jObIfJ8a4u
m+GNadzEyFDyaDBuwPeFY+yF+iiY3soeXQ1kvzFvKksnwZpaz7CyP3AwUioCDSGH
37w2aYdDuSQW836pUTRzNLhZq6bz//IJ4jGlA+UQeY/GmxX4sJWhXcJgoW6rX2yl
Z44dQNFIJplYU/22pSkdyemMUIN8nSQmcNc93K+1QtfqrKhLAMbnlHlXtFYvA71R
4AvFtsSAqItY+pZMSz5ljbUNMwGwdBmPj5U2G4G90SHATbI+K4BMdUoM4QUph9Yc
`protect END_PROTECTED
