`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+2WAGXsTVvnkXxjEDPhuwBOAPN8MDSwszPbSt4lsVcfKVGnn97XFD5balCKAbrrv
hDUioNdRCC7v241+Gi6jwv1Q1AF4lYIsyV+Xc+XsVd3mtUGYRiFt6tUGbAxqCDfS
+y05gNU2JWWoX6cShzZ8NYEIvmng22XPbg4+OqZ19zZrzCAaM4vFlU9z1cGP3TCm
zCp6Jwd29KsWMHtbKkJg+ux5DGXd92h0hMovdfdGTI/Tjg6BEalIKjS1R+aNJada
eMH9SqGt1DXvdJEzDQDbcgwblnuGmCMEfhgOIXTnWaHVeKOeMn/mIEcifoeu52eW
/CaWY2f5bLU+K1VotjG4PTSzRxaFg9ivI3l4Fh+2+1CQIfnexe2IaHv+ho6lR4RK
g+7YTTW56vJ9U46myh0LHqzcQ9xT3KfdowmCVMDBtJk48GqSih2tLiQm6jvuxnIF
RXLWWGV20W4wpLUi0vcCL3BkEInC+pCB+uFp1MovFQGUGlxSmRwHjD7hvYdajSer
6ric9JQbQmeYM0kFnjVB3Vw6FvyE4rRxE78+Wab9y93h0xZJ8JYmjbZq0/BXPBlr
H1pznryHX7JDbqUZiJQnJC3QNyWcS5iqnmLTx+s1DwOEerP25mpXv8HZFMOZ4QQ2
gX+CMoyRZ0jKETal5YpHVQ4GIfAMC5dCsaCIwDoV/GoVl55SYlUJbVsKmOLZ7HES
8ibVFo3O1jqaRqIIwMozWo5kD+GUznxysAxDDq+zDcOP/xM/UYjG5UTAM9qLX+qL
`protect END_PROTECTED
