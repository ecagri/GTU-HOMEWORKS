`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pEimCcKgmZyD9rqY6jGQGohiRgSXXGnoStzwUbPV/Wort6M2HCnTQ3rhfu4MhDQu
AtjmsfxqtpuhscsdJ55Sf2e9YAsgAXz+UgcDGrbCEg+JdukywNEeh+e3smTEC45/
lWC89D7RsAgSMgEQcENI0kMA3YuOORAfdWzK/fRKs3q1wePZvhZHUmVVjrM7vG7Q
jlbiAaGxqL8XgytgeIAmgFe5g3fcJ1Hu4s4EAzXPL7r/HA+3jI/uiEhtztPu5SMw
mgApQUvcHCpR+YXYjyE/iSYE1SO5rq5OLmbkb5j87eAHFpi/yQRPsAK4u8jyuxcD
hJPrmzeyJmfwqD7Hc9rlziLDSYJ8lC7sRuMuzx8SeLdpqIEhKNyZ+rJAbBzKoA7j
a70huKhKpRlGyI2/9zAl83J7+TMu6R9WoKx4Wjq52fJbFhSuWdtbW9A5zJfZyui2
+DWqrbDm4e+OMV2DQNye0Qx+vDTRbv1xP1rzLqRoD3S44a5RzIK580ZCZ784jWzP
jokyv/C0s2K353nGd+I8+usx6hmNuDDurB1CO0aQ+0cUiLX0tVZ3U6+gza4L7py6
gbbdNe2fzxTXeJPzIljnNPb+CxqvmlbmidwhtK02kgggt4hoaq7V3B3Hh4J77TH7
gz+j75XqpsEaNAK7blcshMiOUHoGJtjk2s8Br8qUKtEN73uvr4M8RsdnhvtQTv2y
`protect END_PROTECTED
