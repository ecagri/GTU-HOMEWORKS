`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2P4JHkL9gaYSln523P7IZthWu3W1BEhKhOye+KbMtDEmdHPF8U8ZyQ+PpiK3lK3C
hLH4dif3x04/AUYVK8mRDPZYe1b21T70bXH4CFwLkCfiZbKvmT23cGg8JeGak7da
jO02pVVNJ+M51DVe3wm8u0o6SemrDnp8uAPQ3LlvPCvhZVlSOauhciT6C7aq6ZF+
a6mTYffh+rN2J5S0M37VKtKpj1KL9pyH9Qypn8pNaadU3YNKP5Fmp8pHyCL9VgYC
jcLHUc6IdEFyRU1mioZHEQppNKsL8wqTctuUT3kqotma4Q2dDAmjPnvsLtXy0MJR
jc0Lw6hQQMoT3y044pYu79EnLBvfMZkiPkAf/v/LT+Fb0JFPIWfsyyR1/NGGpIAB
OF3oxNOjIPeva4YavVWdOOmMICxdfWrSXnI5C5Pg7uJzZsCfjd7LkuIH3ytVmocA
fitKnBpu3sZ6odmjvqk2k6EPWIduOZDomxf2kUKgnVyWahgfAVBboUbReIcgB4o1
84ZCqhW2KWbspJapRtM0dPJpffJvRlWy3Wxs9guYGWcx848ouQPRC5XPLWJdc7q/
rmXWLwvMAC7RsMYVsELDeA==
`protect END_PROTECTED
