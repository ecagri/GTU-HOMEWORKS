`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RdSj3aUQ5Ger0q/4ngpqQWW6Fa+FEvcA/QgjyEzLFnU09ivzMDGwcjOuT6YsKJq6
60b+AOovPfl8mpakcNVZ9CIetEGFpaEVtbe84YrMjzF1OS5RIBYe5I6DrEkNw4Xh
/jYEQgNA0mGPTecMqA0mtITCnTEh2hn3UN9Ru+pa4SQEbWIR2+FIS5XfYETYFw3D
9Ogmy9dT+b/U4j25LG49+iqtgpzeMR/LG0yz8zNO1RvvgO+BIgKlj32O1MrTQTg4
aeGelhxswt0ooufXwBPA6C/xMw1MKVeLQ7KXM9f8K/C+eiL/EcC2R9YZV/4WnhB4
Q7SQ7PPnw5Myn9JXp4EqodPtKzPu6yoWbKEPsFLAM77J2ukEXlbsrsj1NP63NN0/
tfM2+JPvcffgU/3t3jSstpDm+SpLDns7NcJtGybRMXG/nIc7Hb/350KUvyTwy2tA
XLsopxYfuSdwyP7WFvRAbdBa+q5+fR7AkX6zBXcXOr+M3y9p6iZnUIgQ5chYOoep
fwfiAMw9tsYY+Zu62I3uaoakv/LwBRRyNyVzZNPo6cY613HwMQ4ZGtTPx1GL4/p2
WgTyc6NIbulQQVPKY2Cf1cX6z7ZpzA6rfqZbajvl2RItgEcWe8pSX+jIb7mfvBQw
XkJtpGFJIbqzrL4Du7VUAfU2FLswEP4Jtgc6cVsPGk+7WoZQ+1IHnaEA1zSXBhSS
9ct3ryOr2VthvyMcbNCf8Ql0Jv/aswn2HTi/QSWHiQy2fPObQEboXV1aN89/m9FT
SM0sEh5h0jkoU1KW1uz2OY3yf6vMHAD2GOyJbMHFbKVFnsj4GWeA6NWFGt82WJ2b
FeEyZCHAo1bn2qTgHwGTROfZSMmPCQeqOzJ8FxSA3nsL41Cu0eKK3OpVQ6BD+pj9
hoG6A55IQL0hdKO+OXyfSG5eFrUucn868HyphVkJNr8C9fPNFcp4tihnomSi8eox
hYWaD47eKJ9VmpnJUCOrgBeRjkAIoGealrj7ePCmvNkEe6MjUfZMlTup5Ii/BBE4
alqbvmCbi2iQkUWdCg84JT/Q0XUvIdE85WTg46HAFQGUekDNOWwgIL3JhGCJuWjh
kZrIwKMF5TB2sQKJSEccfen1emPAhVNQdLg031fknNPRk15bHmG4JoOzXt2K1629
+O5yEVyd3i5y2h1HOwVUvKFzzHzNF4fD4RaG1zt4ytye+mvXZODAu/j4iB0UgBCm
axm7iP23lGWpGwwNaBxQPBb3JPDfhG9HLFMBGjNTeokhp2UNG26C6HZ5kHSZti7T
QY6Tdvu6ZdRMEqbIFFjtoDOs0RtSrMmefdZjsyhitUutHAA+JGjLr4cSl3s5U3fn
RFVG0zggDWNga97Mp8nPCiQ/7EaVQMvI6ZfRWMZGh01QdDeg8Vi7XITUuuav1D6N
SMAgRP1x2L5oUTxi8OC6CnaUdnKoDYR7MtnWXq3CheCcOvVjxSkWqdR+xqUzcy71
I7Pz4ISOpIQLLsKuheHdXbWVaUfVeWhzMfWzlCshLJfFOmjlMI5adCRRy8YiK9Ht
qV/bW+WeuMpm4Mblffb6r6/6RvNj0ZLc6Tn/uEOS+VdoJ0Bn7GZrIXW+bLDWHGfM
+CATx4vjGYWzaaqExJ0XVCxVO2wh9pXyIGjHd9RSirpBmpMQZbL4lLcQpRwm4/Ow
QjPGqVFQXYwLS4s6bCUUAHQcJjwmi8QMU+dyVAsK2AucGPdteTWL9TAApfuSb8XC
UhFwBNeOqPMW7YlFrONvgAeO9ORfd0M9VXH0k+QL3dNT5Ia5YrpExaDpBAh3hty2
Gts0qw7Voq8f0NTtaTYvrFxXSRfLzlIO87UWfR5WZUbXR4ggpMZobZSFcs/TsV+F
W0rgEt5F/PiZ98xJWRAfo7fwbQtfBbwoUePDGLkOSeld9EjVSVljec9FWc43jJ/g
RwJ4DMDkih7U4NZPmBmlxy1bvGMrGri/RlU0zaECw4Z6DXHSmq0DqcP62A9en238
/wGcLy47swCJ0JpbFYi4UqVT54qM2MBnyTtpIHEklZGEfCqPMHNQsWbq3D4i2Msc
IuunUSZVB9e42m04iWcU8vqRVigPfZrEkF5w1cJlr/b8qSih1jMLBBaV/1oiS5JT
LagKVmHUOpniWhNilHCLFXkd9jVUmsK5YnI+Twyrft6tSoxqLaZ6kCN4cYyaY5UJ
Vq4VGaN0+dCGr+Zsps2fo0TgOb/EZM0RyjiRYQqQYBaRJkqwbVsZbu/fYcwUuxjI
6ZBPufldNDFSrFjdnkXNDVupPhvux3J4/K3T+65AZTOMLsQXzGExSG+X+xJN7kcA
3faF6v7t5mL1eGaXoeKY/yfoeh1AoRbaLpMUQF6ZFdiF1hf0UnWjIv69iurbJ7J/
rWax/s5556oVf7BZzJp2Cy3SkzHqhdIgaLcfoXXDJN8jA8nfAXnjWWeBTMvSWOw+
`protect END_PROTECTED
