`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IvVQ6TG/iQQ9Z0/Kz6tDoQeMSBXcPS2mXkbCH9MlsvGUG692hOOs3JMxNDPyr5IV
ic6aNdKqd+DYU8khcrc8Z2PP41Zgj6vUNVDrB8XJMcJD474rgd65/ahhCPSmMn0S
WkwQ/BC3pL4qf/rzi088X1gSksNkL84wI1acrBvcZEZg7N6UGTh8v4MDgRhsyhJa
jCJqjlcqm/95crEZhYCreRtJPpzyyKz6Z466IZIAK9aPRMo/51rtbC32jCxeCmSv
8PAnkapthgGvCrnRq1iNwqHUu06GGQf0hwK3bFycUnQIb5wkgLjvXHA3kUPjVsH9
v6s+2idqB+IfCo7INMbkXwntQaa7dzcdxCwHhmP42+jG6DtCrIRTk12Ca5QywOeu
i/9qHuFoPZwyUAEOHUGTsVfRePEiLBDOInTBmAf9dJ7jEPlMTuPaGSEoTo8J6ewT
YfOGZDQzr0kpikXvAJHwMwhMGhOluQ0TYHE984IZqJipt4PZRplZxOxVevhaScGL
9mRcpKt/Z2p3xKU9CvqnTrqXgClVM0fRnJUsjxeIqiJKCTdeUCm9kdcAHsxzl1B0
wJSjRKF5nODTWgMwggpEFiCIzSJFch1ubXUFI6fihy3bj7OZ8n6K4yBtOAnfiXIM
8aQOrRr1P6U1s55ASK7u3fMwjDuZk16SQ9AY6USSLyOHFgfc2E1RYqUGpwlDRquh
TKArdkPGYG4BfjnwDGZ+TlLNu6Hh+CqNfBp9Y1E5HelCJ0/O3DGnlCfsypibumRd
ms1D1wwkGTBd76R0K9IYiiwEH6T10xZJ3GtryszagL0OX7ti6VATusm8RKlnkXCy
1kc3jsxDuGAvKAJvZ/Um7C9K3EPS/pQ3CGa732lGuC7ptq9u2dg6CJs1W66R5qCF
Yzi17F7xXeQEhf97cLMmcVV99+rDpbTw69AdRvqxawA6Y6CU2r8WMiInJwDKskIj
1y6gVQjwUxj5/r54p82g+tYc0O6rb0EG9+hMwxAcoBLzJaqEf3sC+BV9SKuGR/tC
qUcjmEWtUHYGLU1Hw+jXZejYKZywVhP2zM5f3Egt0/I+QLHPh7WdvG1AwHwQI5O/
SeRF83X+SexL2pAt3Vsd6ykUax0xdv+jfpXPNm8WotKNRlgdOB5is69m3pevi6yb
mVreLIbqctktZ+gys62M9fCjTYPZrJfAhAizmw+EMyN4ATALgP7/Hz9LMQFD3jHc
m2fKdJhTbbz3tXIB5+YC23iUfNHt4/T2dAbBp/hpNJifeWo1yK2rgNh/wwgOH1aI
FCA6gV5ky27w1TgBoV7aHtSmzcpxjK7X705T/vDVnO8dFUoJIAM0DyBGxvjGdjhR
ITX+vJgnH5arFv8b4dpIBBI3Awh/YusrwWSmc5GZCLZfkgRl533WeiQGvjmszWKN
6gvDXhC1fsZ0BXNtq+vOeOgX9SugdHMYPnIPDBJral9ic+hl02u5Z9pRkQscQJCt
sZ2VnCCgLZnbboP/FUkyc3dxAefBd5qAPi3BdQamDkGMPghi7tw7QeI+M01nawtS
jqm7INnfvPAkTuSqCfdMso2HaLqNIW5HY43b2UWAWHolWGC0665FsuhmpRUrnko1
5r9RSJ1k7pULPjXoeqhlCytHv5ZyfSRKc4QX9rWtSBGXyvCq9mtxOg0TQhnhbfCb
ki/RKjpIA39WgmDUiZM2R5jPp2GmACzMKcLgvceeLrM9lTFW8fQdYUx0Ec0J1rtI
vZiDa3LnnIUmAk74tmw0Dr2wfzbx1Mag6d7IIjC7a+5387l/mdRfbK2YC8yM4ZsZ
eRNW2SdBU9frajwOC7rke5cGefPttAIbV0ex/on6mmZ5FdrGBVu/f2w67nRD32B0
xPaOg4cNPhEzfAEyaTG/I91si9heYRGIKApw0ejnwxL53y2Ab9PaCdhliwjfU6eE
n5KfLJ1OKrWcITRtkoZ/nanbNg5Sv1etf98MNiy1iz3AaSAvhCSF9ussTUUTU46J
f64fjvVAsHNKl5n2PFCzooKXqvJeop/R2s6e9XIV8kMrtVlh2fi3buDYnZPj8GwW
OsPPRZXo/q552pNRzDZUvufUsTioCg5UXC8Y8tKjN/5UZjlIOkHN/QOdM2vIp6vY
c/sfJnYiGIhtVUw4h/FdcSKboClKHh9et8mh7UZZqZHa2UMkLVxcqZ6homqBpeuW
jY3ILoYiK9PG2vlXzGu7ztr4hHqvJSWpWSN7mXk2sR8NNPUHYNJp+z9UTntNMdfA
RrR9vhqbrBbJR0rgacqtw8she9+QayfjKBkb/CeTSGumEvepXhCBzHtRKqZBm7Yu
QOmAF5JHroduXCNS/6O78Ykkfm+fnJK+kWcxPOYbFmrWB1wv3mr6hn3XLb6szM9w
5LnWpXL4DwM8cA3FkCGIh3xlLkjL23YjXXCJdUZQA7WD82NievZV4edL30vPD4ZI
gLSWROsCLwctFrJet3tUEM12Vgb+4+cGn8kLzxvcgRmSSoIJJXW9ZfDXkl/2cfCv
duNXsZ+PFOuMBwvAKappgjJiSDDmXiiqh+WJclsaNogVOTzQ6lYTKs3cPXyUB6y3
3kHcDfDMp2ipVW7Yk9xLYAuoINOK7+aEV8AUKso7Fa1+ZneE/qmz1OLI28LVd5yw
fECoMLv35/r0WxNZGkjtiCErCegu4xXHa0vO8UzQVum7BmG0qYZvVmpJCmx7r6Mh
AXTiRmJhosjXdaDvV6QVFhIJLgtKNNtOdhsnx3qjfOxzWPodz9D6RxZk6Ts7l85b
u9JtTRwZLDmo14JMouihH/aqIh63lHaTvCe6xVEPhPNVufEhDYbL8xt+YOgvGKhN
ug/8lAyPsWZXrLx7Zh2epVZ7qzathGSALtULhQ4mADQYzjZdsgRs6Sbfdz8C/HWa
5tocr0L7aSddEIyRS8/U8lI1Fze9XQEG5vXHM3oaHht7b44h2cpCbA+J2WdO6Qm6
AMJgH6zQBXlujcR5WtF2xFC9uAirZ41Nz4h+sCC8mJZGjQj1lLGKbEq4AB8HQwqa
uVlqkqTxTYuCykjZWWeNn0wNJ31UoRRVBaK2yDDHGUPCRmVvWFlpMFQwao4xWMtl
jTOc/fPICkfhTxvOVQuGf773pk2o34JimXS4iNDbAbTH+Ex2Bkgbv41zHx5ZDWvY
QdedahSTImVANgoCcWwbs0B6vZ9Dg8EKzBLEcf2sypnRQVDL78QqZombvQkhHsDG
24HxWTGKTbteIh8BZ8vAwHa6sOjr5p/rKOhqTNI6iv0pms4HC0dR8pwtwL69CQZJ
F/XxN0d2g4vJm4ihKOQkKsP+B4hjK56u6q0c4glxJRrth3sOsSRzf1ZUBbQuejl4
3kuTKXLWJGrJ8mLzoPydBHhoWBPPqHUYy/4TAfMsDXO9SEw0Clu6yyr8Ptp2xWFl
AtxzAvz/UTuE2yJWibYD+6I5YPsecvvKj0d41q5MMdz9SZVT8hppKxYVBTPr1VXE
5uVa9xLvA03VqbaLdyuRGOvBl5d2y1S3AFFp2/JBTcWFA+cUluFWzkUiWiVJSGFS
5L477jrVl9vp6VEeWLCeJbCxBDultZNzDaHSUcNCd1F2dl4f7iwG8ec87bX2bA+5
8w5hOlrDzP2sLaYxasyBBLMEAJE7BM+xyQcT3U2ZbqjM9ABNxDrwWOeV9HXtPHK1
AJgxxGHwIxxfQjeJ9RfySw1a4b5+0A9sb3kKQJc23n1RHQ2oxsXhldMotwbjtavq
QSbefSUP98jVXxfnoGGRed9yBWReXiBaNxwEaZWpBHxoNLR//xeUDicDFhMKd7FW
pAFT9TgWxMKyacN4UIvtiWPj2voZzVl3wSjTN58ciay/5Fx/h7s/A7YbkQBGafem
2IfMM1yWWOnL1hyJYDgbaw+oDuEOEclNQASWcCXCR5CcAmnR8udJ1VcUuv05F/Q0
t+f97V39XuZrsq+h/1njN3h9IgPcE2xQWfbSDXPl86w70RHpMtCVEvzSOw0wP4wx
tyxvSA8vRv/XhAQwU6ZtMimQQ8mtgyZNsT3swS/dtrjIcHIN33TERVikX9NA1YQ8
iK/ocD78WaG+u8B2OvV2bdPs6cqf/eKm7caCyLl80NCUhls4ez1dKPVDYbzbgXvD
gkFoWCFmkgp2tDm4B9Silf2YBhQlmLWrH0mO0D/qXhbeugroggCiBemIB/N/uOQA
4uG7SH/WAg+HH0+rEmR9p69Qg4JVH8dtEqrzYp37DIBpBNRdQceupVOQQ0epXm4e
v3tYE231qcdzAi6AAbZuuI333VKAu13inxtF6Okyq5TWuL0p9/qQtHhTYik2CYqP
EQvzs5JzPztGjKpeQYyhNEjYEI94VExMIxcMs/tJATqwPWJjPMafyOff9MhXHpBa
b7Ge3qA+sAKygZAbnjS+ZoNT9PmoAfNjSaU5B3RwdycV9BZTMaDXf6Qsu9ymMgyH
mhfVSuKlq5nsnG+pXYBD+mKPSvetD7sCzYFYzAFiwpClQY4CVOcpF48IUB/vTKjP
Vqjn9tQ/ivK6DqlpbsuI9spoDXvCT4XvR4X6dpFlL8U7yM0FgOCZcWktnnuuYF7O
c/YOXtQUBN0FI+xPDxWVVyxWobcBf+Qcq9H1De44Fdm6dGoxuHTRPCiPjimhGS7b
tw/tZ/ErnIVFpbw9LmqMIw==
`protect END_PROTECTED
