`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ozjm+n6Kv3uwhvNZY6pklaqtLCK8Yi8qfQMLez+ClPK+4w2pJCOkXdCqGmYcpkZa
beDpQooyZoQurpoYbKrlo3LnwK47GYDF6oT5N5E8DL6LR++TsuOK6E1cCx0W47rY
xxVy8pJOaAO0DjEK9QOmcSt3/hfyIUV3QCIT4UMzx4W3W5LHpnZFrGBa4luvVARo
s5HGAX955+tyIQSXd6tuzxTVsbrpmkVq4GrHkAU9LQ7c1gM/GI0xrQ4t3xvZVFHj
E3FPWrwJylfv5abbbYjVTf2Sz7zUEt01/RIDE3tbjUCRlXEEU3+RdSYL09G1J6N7
EAqomHsNsowLKibEdXQAQoIWpRTWL52m/tT7qNeE2aamkGBZfsxXOUSYmtUgkywS
4N3fiaO9xgh6ylgD7ww3WEmBdEZ3kXTI9rndkFssHWTSD6bpOwEg3sCXA/mU4loi
qaEGrNHNejvtzty3UYIXLxeMgFa2dRj7vZvOEDdbq4VtgccMz+/a014/9+wxVbn5
O/SUMq1TrwSl1ATkg2iMpRfBnKGUkVoa7LaeaWCBikAwtmrRj18Lj7DK73FRRk4u
20aULMwjNGMAiFZ3CzzAbelIdLRPopMZnDNggWUvQ8OYpReaVD6ED97T+QsWpl4c
8fDEqXUcqr5adaKcRSuuqaGxoG5KIsYK83ymS0QqRktswvBtoagOtFBX8t3Rodh7
06nfi5Omz9/PhPbTUp1f17mx+inPUcujyxthWHReCM786NVsnixczxW7KQlGK+x/
ViH0wweCsDmSGuwrGnl5sHrQ40nDrviZTahaCdYyjtkv4t432F/EcdsUdLyZ18TQ
GlEpZgqJ9dYjVMxtQjQ02zkvWIafXORDeJHDoJX1Uc1nKbAVUUEO3UHEwnebuK3r
cZe24m1EVu4BDnwaTZ2U+5uYGPLCGvEOk/Tvd0YsAri2mrTTiLbTeBSCDjge/5Dm
FqzzDQQi2ZCy4bsC/B6/XvfkQ/oxXs1vSYYOqomtOTNH0am/qDvzXzhYyEHQlPwK
ef2Ptifnu4C8SbH3eDK264vNX8nxRprjxoNNgHmq1USeDYDIiEaatL0aSrvpEwfO
Bl5LZqAxSElgoobYKru4ZXBtBESlbr4zAMXgJQwnBQwGOkaUPUm/H4yZ1oMDZskS
MyyiG4f081/5hmprFEL0/MUvnR3yjziew0prYccTLN64HkKk7Ho+TMa+VUZIki7X
4hWEhsEIk3RPyLqQa6mvwBX8pCVeLvGAT2oOtPRTLBsD0mbSziGtg5VXSEDBcMJB
trLyMyJpwDO3ghpbY0QqcSDs0SQy3GamZhgWQggCOWiFsyP6e6A/mGVoFeHehzp9
k+H8arbosI4NF5cDSbfZQLfzI8YwHaFTuxfhsNor0urc7N0q9CWdPuBueP+YnbsI
YO02QCWsGu832zdddAgoSfD7uB2PVihKapTD7rfiKrufx0bMTZ8We8CZr9VG2X2v
JFgtJOAwCGzxGGuHY4DH3n964PKbM+up+w//c1JhP/dgPSgO+mkM3bY+BDHpL6hg
VJx/CRiNx/4ml96TdnzAj7pH1HSbqRMp8cFzz0B+0OB+Vs40CIT+j4jq6UnTqqPh
8bWZRJaiTxkjGfQsvsvDx8mJw6CfP+hv7fOnoKZjcnglwpneGdDzHr8nHQF/VzTG
0HW+F14eKLe9dc8LnuanXIaC8dyB2bsxi2bA2X39mme6RoNz1PSY4rbj3z5Dfe+6
5TV2qSxbCdCmXYWTx4ffsG8MC/Uh9H7CyUovFIgq9lQNCmIbFLct28wYXlXhGeZT
FvlYbDknnXs3r7HBa4b9pEQQlVMlKzvG3nBv96b6b/CnjG4A+/JUmBDNShgWAPNi
0cFaEDsdb2qIGduCoOpGVdRsS31ZD6ybdjLeKMIADMveH+sNTVGbje992akgVBY9
yqk8asiKFMZZHUOESriILs90njMqZ4zX3POcrs9qGEpxVH3pyOZrKdmpW3CZWciN
CkZcek/Ucwc9dL9IZpDekAugR8z35Sq6vonUYuHwpiNMhVS4u/CUuQ+Asw6tInhg
X5g5BtAcWvLeSrZ6HZ6giGNelXNUGT3ml4LHJQxN/e8+6YQFw8RmUW+CMlj4dfoq
ifGX6qgz9+AVLHpu8OqV8hv4Y5LIQJRONeVBGVFQQ707cmU28jNc706FsvwIYMkT
NElJ8kqdb7z3BVCUZblDfmEGPaOeQ87KqVuB48zyQDK8N7Q10YPSk5A/cTrDa+Wa
7vXcwQ8ow3rdb0HZCwZFmrpl/XdzG/KX6ly/Tr58jo4tuiPj2xsCiP1wdtoDedrh
1trdTjECN1EQFR81VaHkaFqPTYvRqGsG6pP3CX/g4Vo/eNkDI7ALLoipGS/OtFJD
NrCzRm5bBTaQ3uPpNJPuZzudekn7bJl6x+lxm6A0aCSiU4oXi2DBPEoJc/WXZPbr
ZNM6cXEPCIEPCqYGtM2y9DFUO89M/VrRmYdElrvlpEjnp05uaDhs3zNP4O1Qbk+p
nQkTMv2rg8AhH9og0SZ0gQV0ryIHMu1pW/KKwK4vMhhyZzH0WdNLVx1Vai1MpNjJ
NFSDcBqYt3tEmQ2yhQIQXkUPsR7Zh21zSQX0zr1q8cqV1QjFlm7bxPMLd5Tnf2Xd
AcpXpQyw158lP/odnYHlVo30Kv0mYrzCMKoZwiJNWjF+f+cEdNNjexcEUN6Rxs1t
EIsKXOH1CoFLeAIfyDf1ug==
`protect END_PROTECTED
