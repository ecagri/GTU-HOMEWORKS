`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
do3jFCJuu1wjdLTI9XmRDqPfOhHDU9/dB9b1F9RqM1pKzOJkoocv0vEUVgbH7FGg
Wd7d5Tgtg3PPDhqROjEcEhpLkybLgD1Mq11CP81pG9HmqM5aRP+nPa3TnBK7vkxP
Fk+wRWFLS5e4YNRSf3XshMP6jENTN/JTeVLvV6kG7hV7/lLiG7x6i6UPVwQV3oN8
s+41TuFzIbEQCVIvAzHvgEGL3pDW/GUc+6qtm5ZA4oOnPXnjvcKDLXxwakNXyK86
r9liMSeYW4nyaWrgrmzZhaiGiv4dUrq5yFOmL328igu73BMItHikfHZ8cDW8Gtze
WYjY5so8NiVf5urFwGNnFvNYhsWSowCUJALXVQEJFVqoeoV6cH8U2T3GfoS0axmM
orxXA/XDJhHZzGJ54pAB5BsndwY2NANqq72MvMo0iH5A5ZVq1I395AFYpoGh1zWf
oAgn8kwHzP7XxWAK5YWjQrN7lP4sErDIOvDWUjVRlfPZuRtQ4yyFlIE54oyPzrVm
`protect END_PROTECTED
