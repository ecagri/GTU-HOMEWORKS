`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
potalIDRyK18R2smwh+iInXeiYfep7Wa6C/XMTJv4mYC7XoaUWKvcVfv+NTsKitS
wB32WNZUJd4jBfoHqC/xRI0Wu7IFoZ/uNNl2uYjaU2iSAwuiK+KmYuczhd7YGvDC
N4ClUgSqzaSt4NzbhtQRLpHuVNfuiOkgFLKG4y3OZBrszdSv9bJoaDYi3yWWch99
iwbV4jk3XzYJ5sV3UqsYUNVZ/9tNnkpv5veamDUJ4sfQH2A2PAGzDnk1ocz7n6s7
QeOkJMym+KCATnlthTl45z319ILiWqpLL6J8XQPADIKig2bUyWEch1xPVagA81Nd
P+OF0lSClyHYG3Ew+zZ5/NDWIcxTtiXmEZZMpekydU5UjSHLROsMIiwkEvVDS5PV
9ibTH8pae/hwLa0zOBh3qAuD6xcxPj537NC+B00hBA+Yxuo7W7BHDAJl5DGav/aw
3owapCpM/VXeRKF7sIj0upVNfPWmEakI3gxix6oS9+8xIn4yzPT7gvNVl0V1qAV6
BmohDiEqPYC+sYgUvl0ZtHjC3ymDjX5qPHvjK77FmTYlsj8cLXF731zI/hwN4ABl
uioswCVqWSb85Qh9RHn95WnVwlarqAgcaV4aUx0a0880K0naZ0WxiI3//xJG+jop
3qIYI4V0DAkudvdnvNCeix+zkTZTMT8V24nDKFijGJRewpdjcOzjZkRToMrDVxv8
8sdDFHn4kd0G9FuG4+KdrAjaDZaPtT/dnAJ9aNLIRwh1xIs+2dsiG8z3lm2z6ETl
IRUuVS/zvAkIONHJBP25Gom7at4C8oZOlfAIfwHRZLKhQ5V3rQxCROEsRuIPN1E6
b8zT3kK74dDDoY7Q6UOu703acpz16orCj0BwhYb2TSHDiUgdIs+me0/NxoISEu3g
RLVSKXswp+qpy5xM5sFWJt8CNxE7g3itWTkenu7pThie+kfUDToARQjGwy2C24y9
RIowQoI1IGZXPGY7OpxTqYqZ6tHDmw6ZBG7c8yjzKhUiG9srerbrsUnu+/gfpS/P
H3BaaT5rHFuOHeMvMkE1b8DTO0oa3R8lP9twWb8xqJRFwQljbIq5J/qQDTppCWgj
wSR9Edvj1YaMW2KV9ysTDoAM4ZZwUzcLQEwLv/h4W9ymnW68XR2LlxUB5039525m
/O/RCxrREzRxqwE2wtko0mbKI2A018vOf/RKVky3s+BvLQB6v1p7jFWfUgiDjLEb
G+CJfTvmuI45e/o7TFGf0oc6AnkNGcQBs40u0YU+g/8gxetWwl2xcuyfpi3SZe2H
k5mnndKeFybdSP+fzgJaI8aazSrwZI726ik54/KQrl83k2FyHFyszYfiDu3pjxUx
Lv49/vfIKm3HbS61/lbqGc4s0CWfj9dVK80bJuAgbWNZdZifO32IS9NhMFsbKQLL
I7LN6FYCgvV7h3v8Y6e6xm6Bgi+p2RSQ6PUQZkEFq/mdNEHCzn4p4SiEnuwmDCRU
aWbv+y1jbxGanIOfUwhtHE/sXVlCKByYtN7QWg9fH2LNDpY02gNMs3QeA9llS1Xi
OhilUoBCQBfGYk+zK/tM006bOjyjW3WU3oHAcN6IiiUKNqe5UoBzaBLBJqqkJLFt
T4o8sMnMr8qd1ejSx04GZ+R7nSjmhTD+XkMD352nNFIUp/eXQX96mXszf25ezZwy
H8yYEec0BKbJDtafJIRWKilxRZ5LHRaXHgfWk/ky8EV+6QMH/E2O5N846O4CpOvg
FFnwJU5oZ3LT1/CuDe27Bjf0lknjkPlXMF1l5b20yqqvL6IrGpi9uzmOso+kkCWs
W2ZJhOZvWtArvhEJrA3JXh88J1GECUPlMfNAlAjzTbKX+WePlrbGdiEn/7pslqvA
8i4bVjHz6CdQq0dNFGlFQNbCjLwcEth6V1j1EJ/8aeq4Naxf900ZKjA7doo3POhl
zkmrFsRpoUtkSh8cwB6nlCmEAiu4eNPb1VQ/rwgNHyTp29bC7lWWV2JqrxlhwKOq
Yzvl066alpYS1fk6vh0qmLfp+NYQIylO6ASSNMDFcGCRfKMnNIzQ2igDCwORM6mL
rg/BOGHXvVlPoOYHSsQiR84oR1hvjWaJtx8y0rH8MdLbWbblFqMEjPK4Lc6x85Ir
xuq7erq1E4kjwIt4MH1qTtpMC9p+To6e0cZdC0iva/MilQDw+e4Nz4vbSbKjeLvC
XDeJYftylbuHwVD8Pg2rOE/RKr00ciA09UIYi5GtlIS3lMXneu2zkmLriNK2852R
YCqUUAAOVIHUVsi/qDq7/pj9ahapORM6jjOXxZfNTEE=
`protect END_PROTECTED
