`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5TxxPdyqBFBeDlw+BAOs1XkhoAkRPqjR2iO4ZMv3R0h+wxTHVOk4gp8mnIoH41iz
ww/utJ5HqyRCfhMg4rrDw/tDBgMMNhdxtT1pDd3TsghY1OQgho3jN3K3piNcT6VE
gwazXK1/Ug5qhMR9bjop5/yLh9cf+6P2+B/+dFxHL51wuvYMXWzFTz8biHamImRT
RG0W4YQxSyxqzPOF7mfxFDQ3ly4b2RCjVrwweBrtg/4ZNjYvdCRp3zxhVSzoPZzJ
tiBvMieCRPmRMyskXxtBGw0eGGvwllr8b5lzBqmk2/clnHpfpyU1JYMvYEY/8M5z
qO4jnyXNj3q+mLxvctJIhnHdQVcvy+S1ilMvYkM5nWLCXObyhZ6PPC+oTUppQDow
bfm3d8Kl5Jp3Vkj1ZIokueeWvhjfOUXq3uZ2eWw44CSXHTHkO+TQCQiRTyKNub0V
kTrbbcRiCEfgQzh0ypBIDnWfS/ctWqx2Uus+BAFuWp1QY/mwc3LvKx4Gp7doxLnM
YVBHeDGt2++fkD1+kc1MJYPXICl93HeG5RDNRKN0Uqr4vXtS2fZYlbxfgP4TEZ4v
ypzfbH7kQiiMt6ivMPvcxx4DAXXetgQGutIjikMhGBdE8praJkl96eTVaX2sSN84
jgTPJgY7heE3LuQsVBspfbLM5OjiVzwYgEsmO00lH0I3QemvfTaII/9erLbjMEuC
9FGw4mFDrm+BIdS6I0G6sfFDEIZb0G5e7OLrFo/k01v8tdh6JzsokgZpv9Z2gXNj
ux2VSj28tHOe6nMPGKWDur8SPEbYnumDZZCWyTbtbzAqRa6tEJ0EdH/ZsHYqZWz+
6nHYBBwa/cqCbvSGCX5Ec3tsR4qlPr2+KLsUkmzaRgz41cP/TjBpfznwkX1xqxdm
rYMzmIH5xOcB0E2EjfxAfKieM8NiRtiRFOxmg29R/f2l6URLX040oDwh360SZWKg
Ic4lghTV8BQ9G+tzJdWklXBxKCRqGPHuJ331FDViIdvKnaJHBYmqTfyhIda6Vgc3
Lb0RxhTr7rCOv97hV8UIbtsiQkoLPpt2xh8i7ejvlcnxtROIVs9LFB0z+oE2Ag2k
E/d8/Ec0knynFnWOW+Ia0rt/digc66AnzIluPC0d13DQQ18idRs+RIHFehY9pnEU
atWmtisbTmA5QDgs7QZku8BKpGbSHzKjdqRmQPe17kbPqxZQfB/iYhFPQlfd8LSx
9ZCtszN2kQnHp9XjaalyD7LV3gMY/Sai7b+DeQtwaN3VKHq2bkS8lrWNboQt07nO
0jLzrGz12zGJDuNWGOch9DyTd9e+a2ASAt+inEiAir13H2bXHzGtzGGT2DJtwz4n
WOjJ7wDSx0VOF6kTHigIASwkcm2W9qRERk0yEXqdRAJWKdGQhA5S3bEYA/nAna5f
lwT77xNSdBUczGK4HxBfj75r1SNZsDhDGmm8tEgIlK7v7i0f8yEbNTSnqiwZB+Uc
I3swXkRDD+8A3Dh+k4ZmONSrbnHcm7MLpeMCyUIf+70maq87M5V1sdNr/uajLkGA
sM7jwGsJTMj10tax4pLu5BtJLsiRXAgp0GrLvmMZxmtVl/bebfl4L7/xMdJWAU2J
Ru56nVpiXPtz/Mwm0Ksl/MSNk65rcdIHl89MVPoYlbksK50cC2nON2gyCFiPpBBL
Q3Yv+pVw8vNqQUtCCtTdbdglNJayVlt97oFyRXDn1LWkqHdn6usqup3UFjRE3aeF
t5dZMwP35SFAzs7ohkmiOqZX6vR/cGmEQbl6ga4KzUinUm7Bdg1qHBoVCB92F6uJ
zuqHtRyWMwqlN6C58crg3EHSs0ndQtWQQN6ztH4KC/YDdO+QZNkTuaa9YmRJuhkE
qrTDz1dWYX8gNS9nfuk7bD8+N8HEOpsBf6Y2Gx4wPpBKZZUn0t1GNonCqg/2ExkM
NKmvWyt2ufiy3JJYwVfsqhuYobc7OVAQclvSqffd23uTtIsxTBkmBTzXIkousrHo
DbWdPcw+LwsM81l8BY8KpJm2wP4UyN3WEtI9Lv5tirsZjd7LPB088HdCpVb2aXmP
tEd6aOEISQFyWH35iw2ddTu08hR+j/TDQAeiQ3l6AIdKd5rBqhDdc0CcCLkrOPtp
+xcnXbZtpSmTZOWhzea/aky/8PzsfVdUupyPLOTJ353by7m1Av83esgIs/Hyhq8y
noLXhOxfV5cnG88qKL7FguRzWNgi9Cy5oxN+HUYZvaSkYKf8xHq86MFNy6wB2NaJ
pMNODw3M/Isj7ZrrzmQjQWgkQpiBpAsr99jVfpYyp8/QBMedrj1gcT102CL7Tkdm
8aj+0fIzYjhQG/PxDAG4Imx5Ix6l8Gb/ltqAjhMMboBUJnTprzSbHr8SFiOQ6znW
5Yp/rijoqaYeubBtI4vyPzl0Vx+lAex1NkXniIWtr6G+bwG3Jpt+5PiBbrW92Ruu
VBFYfqsy/2FmZ5hRW+AVtEbij235L7guuYqfS3eobc8984lbfySkUrqL3k/5yh6w
uPEZHHT7q5mVrc5ihY9R+giBl41s0AJPZfUczW4EAyo=
`protect END_PROTECTED
