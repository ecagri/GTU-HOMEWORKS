`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tALiMN3wYExCbydrtCp7B/VjbuZ8nZfsuwpouCmn2nD61lK2/AJsd2gVT8w1xHoO
CS50YJqBDi29aHt9ErcAByiUlyaAvPOiXeOFtJXNUh+0pZHr3u7rTUNTiiwnh/Ro
SX07Y7C4Y3JEaaXREyVJ0PpI2EpMnt8jJX1p7PnaHfCoX7S/fAC6+HaIznFoaJlm
npHm2Wi5UE0ma9NJbvP8RM3KouyoG02BGexQ6zKd/mAPaBuwcneoorqCEZPeCfkl
5z28ys7J66Jz8/fDRkS/PL6knK7mHJJRFlee7ilvTiCAn+qSNrbAcSVRbySj+CeR
YH6R4nlw80S8otJlrNX5o20BMtuDKpK0yQ0o1j9mU3XZ+qHQpZwc6o6eMk0elhDF
sc9sZ2F4NqYoCL6/PawsEAmi2Dpr0jPBZSlCoTg13hZBg44IwShiMDjUmyyAjAfV
L7k2d7RRPoMLSswk98iuGCawG3xzq+zb7xQhblDuQ3pjWpvkpizhcD1RKIj1o9Al
/sHR6f99l4xWdYum8KpZql6k1XUKvjq/87oM/EBjo7a3M4J7TjG79Jn353v9QGyX
zmmWeJnK8Prt6M8O7W79uFD6J6AR6+lUzs0/BmX4naNnKvkH7AWNTfxsJeuwdDGG
tXesPsv4MA7pxaWJ/Kkv2saUkU/bZtaqPk8b8BCIKlpVP575ZQJA7wqK3Gx39IpW
S5xQ9N3j0TlpxOj1+/vaNDeCBSMuQJ86J4Gc+GA4JkDBziwBh1oxM8LzorMisDfj
Bpr21dcTcrsGQ9nIxixW/xOa5PNn96cPldnj94tE/yvHNETx2Nx7xlU2ZehJMN1o
jmYOqsDzfR38zMI+XwqA9wN1KwA5I4TR+Vl+jdfX3ebYqm02qRdhO7yeezJWLgOS
4m3wABDYWm2+gy5q4mPGzzhmyJi1IfQY25iJ5ezIXhsBNMQ+M7N5JnJSfReFqq4x
0geVm08y4fkXoCytn+RDM6hbHc18O+WKSl/EUAPBYzmOs2MIXRrFVWbutL14uo+/
Ve3xuxcvQZD7Zzgn/0IYLRL3sJkF8aZmHhBN2cPpiQvRfJD6yc0xqcqNrl1eSmur
0WDPAziJkspMlzig8ANeZnmNXiG+Mc9Fgs9JqRQ67b5IZaiVS33AJRYXkgnC06E0
02dLt+smCi8CUyVty3vZ6jsPoiXbn3H8O8Gci0/rdgt6DibwIJyqjsbvmKgW14Xp
moCBDIIgbGoM0GrYyl/rKWqVDAipE0MGFtlQhWLA0ZJ1QNxi4iiqnXkWXLjLwuPt
lYHo0z4QyNOmX2rs/uP2fBsnK+qdHSG73bSe7gvR/2YVesOSpKWRq+wr8d+4gohw
Yq44Sspdg3CKW6M+G4/j5lZa9Idb3BhJvwMs59o2plMh/i9mugebfui1xK/HN1wY
wB12647nkmV3S17Wu+1ckoGgg2XzbbqYjFvn6ZvAS7eGul3Q5tgx6CLHRLQs2wHZ
a6dppRIjmID758WvRgTjlcmOuu8IrW/4e8GdyJXTmTuygMkJGQVvOxknt56R+8i7
bLZCMBR/XG7rA6aBGQ3Q4uUYCKntsq7rjH5cTyN0bYofnatu1B7wa3B+7u3Osz6/
`protect END_PROTECTED
