`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F0JXZso8f1u7Z9EQvuLXdC5xwdhSrLEb9Y2z6F1KpkED+CX5spgmaoEKEA1rmxIz
Q7LL9pAgNlOenQEncu67VexsBiuIAZLtIdBnWFH/wsyo/Wq/Bu3LQe3qVEGqRz3R
M74+3h8zsa+rf0//0XgAUCEJNc4C5wS8dlvabe8s/MWXkqXycSQ2t3VimLGJyCXF
VwjhSjc1Ny2IWpESpAtGUJubD4Une0H8YimKK+IQ7yqZn0za/h6nsVwErA9YY/Fm
GAUhqGYxLuLcBRkXA45Lt6ZLJtE84Sx/HB7jBgQx63uQs8VDMzdSWZaJalZ3W0H5
r2NXNBjmRDuF+ZEHBStzJ6UVKRzj7k5bMKqv4BTMSLkBxytzp7MKxPNbDZ96dXxr
dBNXbReMHoF+17ChmB95AMdeYMMEDnMzq+ss+dOiCeNFkPfRg8KvuEoHWi7Z1n7g
u4B5vQ72NfxYyLUjoEBN+ol2YhnEvFTBRZhtlfNQ+y8jPHhj8378KS9Y+J1oii77
dozQdmye8y8wK9wO8+ooK1kXliTkVPD0alV+NhLHul3UJk7H1sWQQLom4O5XlrtS
KISHZJPFhjfRJic3KQxaxNF8WnbDhOVilinF7i+mLbXVc6QkVElxhvd0LY4NBSIY
WxGD8g1WdzIplzfmEG9B8Or5kWAVtvJOeLbc/iy/r685brQTxPN5Pd7hcHaXgsKY
3dP39m9R4XjTkHZWs/NYHlm6+R4eUz7Q5w3d+s87a27vgzGts2UrVUOMNdWPehlp
eGuY9bv3qqbyaX/tIunPwg==
`protect END_PROTECTED
