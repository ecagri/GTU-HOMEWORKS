`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rzh1HuKeH/EfsUVti+mq3+MHqv+bRsvCxCsUHX3im10o1AvHwZwjAAY4Hawy6vAj
UAMvX2Pcmkn1/SVqaC2xyy4SDh4BWltYa4xiAm4QS4eXU9ZvJvxnKMfnCeJc5X18
zK46/2UlS2HhY6fmRyd3x8PNw0aO7kje2QHqmY6/MlxiIArPacrQn2QI1qn9tSyY
9knIdT77fsFn+Lhn28nhoHgSktt1LdP3pVYI7+WUIW9tD1034eUg16sGDImqF5YI
ROkng7zVxmMwRbQEL8qJcrts2RbSqZNJOKe9Dm5oe1dcpgsDjxtz80agFWtYaPFC
ZqSI2m1yln4KszeYTcq6WBW9rgH5+5Jn+nwox3BVvf2hfu/tzxz3Z77dskaXsBHB
Xe4ZPyF+p8+W64NZevdkpUKs0q1Tr8goMREALDJWenOElQZRXkl7HiA+4fZ0sd/7
jD+HZD6ZzbCqyG5kBPpSm/H6s/7ZlVIekuhp8bepPBdKoYliuJ82Jy8OJygqo1zL
DX0JDMrEYOuYdAsUC2zwRwsdRhs+ENquTRkGBky/6I1DH6aD6u/ED2svlNDKriRa
gCp8760tfwRAM29XAXJ0dvHg47tqkobm86kyFcLzst3D0aPzIXoidU3Mj+fETxfH
Or0tTsEjLcmG/mNF5Oj8wkJVl9mhWBZZrMyRnXtgnEBd/yG1Eav4k7HMaq15Dp2v
PHq3rs90rQ1l4gPXQYswi8S1GKPlv/STH3PNs5QB36TClLgbhigLA2S/I23jKw5D
B1K3r3KH9u/CB3VK7rMQ442jIDasywpONr5RL2ktSlGl2jPwpAkYWdlH+rYg3QCp
U6HfERfxTx7M3iVEWa+XDToCx1AQDfdicD0jqxpSvop13AQ1qowVK3t4ZhhfMy4G
4a9rd1PwqMv8oHFiif4/19rEZ2Cxa5WzbJmuAV4VsOnXdWTYkCk7AmHls/Vfd7rV
D5OlPt/lHd4q1Y9jGWkOerE17xRig5h6a8pLZCiEexM7DC6TorpIqvEVH61BUeoX
kyCXEE6UgiNk0MN17r86o9PagCzXxofw6f0sf61qoLjLHBiy42PqjQThyuTWsSaP
6IKpkD1rt342Rqei+bMP+3poi41Yab9o268K96G5z1MuKxXTNd30HiigVx0uv7FO
O7EDZS9GGQLxG5f1r8QJWBdlM8LW+XAKJgR4j0M3LswLvFyhBXmOVs9XSVHLt4we
0sciDzzSu5713I0qFA1dEv7TgH5dGBuz9MU3T3eUO51dUx8yEag4R4R01NcyoWQy
VKYttmqtqj9nCPlJ1Bmmcm1ci+eaWi6YWb2l9hpd0tx/oX6nbhuE+BlQuHxF83sM
47EtqJPO9XtbVMC6zyHyM+7tP2lcjLIcbcvUgZocAdCS7SciMbFuVsuSqKk5FGWa
DLjOyVSXv+v/bFYsmdACwt1H7MVlQFZAczaFZE9EMtYP8Y2OifeBrVstcUAYEGQH
F39dVx5ZgAlRkxFpn76nYzCbkdEzfyi3Kpy+9AdZ5waWyXs/reBzhcsXflQsIAz5
tlMKyh3r5yp8gol/HXqgNfiaN6KT8DL6s/ek4E9yl0q2iYmnI+wCimKMWpMCj8En
TRgQSa/2OaXArLba9JlpNdm9fV2iomE/VkNsq+qLrU3iogZUCTuS8usXGgHuWn/v
Zw5M3qFwVrVN6rV8RHq/Tk+Qu14x/wOKQ71rPJFbLiqShHOmcm/9NBovkyCYxhYL
I4GsxKgljtyXRfOo3ibYHk+/Dld1jJNRMrUtUOFkiFnC8coY4b8U/Ki7g/J/Pzx5
s0sbXwLt74Elywfnbria9OJdKEWv01jr5JS7MoUsBpT6NV8urDS7ZZRQ3pLdB7JR
T3bboHx2oN3it/1hPXiAX88AU1j+1tO9y0PJviI4F1cBEM4msYlh3XwCw1UdZmt3
jGe6vbHsgo0IXGqEnBoe4h/60L+uirYViTVfvY1qXfYIniXtzSqHvwQUwIcp1f5g
9Bsvbu+NkmUsYlBskAun2PquZ3LbFIJXgj3RqLPx0aNkPQ1Csadhcn90aBvwwOLv
52rVNhyCYYBa1opqRjh7W4CHpr63GN0Ug3yOFuIkwQfGLo/uMnC07UVQlRqya53U
x2mawLOhA5VX+JvUnF7CxigXvrZoa1sIr7FOO9X4zX6GKSBWyzzrTwfokyzcRSWr
wlLRWTWmXdil769AUWIaP4yvsk/5YqPghB3cp5IBekVIEsF4UGBToXwZdjhB3Gnh
8UE7BrtGGpXR+nbO0Zqh2xxGHf0zZEhG/wVEAUl/IQb/3O9vfJNUC0C+86viUpiC
J4kWLsUwCiG6plOuf8kuRW/C2vOWGB2i5EEsF/oIzsEsGKRzkxmwBbXvpDr5N2vi
/9oUjven4BcXsn462H0iu96AbgaRRN2zi62FlW9e3Ey+VOmXjYRgBF82rIxo4GWf
feH6BqgZ7o409e/T8TGuHwv33pQt8bSrVdpdtSe2a16EktCvq8TgyjCgy8XyO5FM
P47zQBJ1Yr0HyPC1P5QPZXdSZ0XxpiVRRnFrDngOY9e++ehrTu4SokG2yDbs3oXz
+3rTkLO+Yca26Jv/z5XJzhHaZmzLAOnB79uC3yOXNlLz4WH8sxkyGHkSXUTnhQPQ
4lPJax8yWUAYm8i7p7RkgUbEy6u1dNipdK8osBX81ze406dSEVyzLsCjR3z3NqAp
PX5PhNk1ycqa9CcL1/nk6c/eKnlnPzZzAA0azPaoWoUQKKj86z1aFSPDdrNlT3dm
CKvmdxpBDYuLEl2Ww7FH73y62KLm22V7TGJ6BiZtyK9UXY2mOSdMmkXyZRhrAXdh
Ho7ox9gzdkcdvxKRcce51puKp+pe9B/aM60bwj2+FtWonIoYoa06jFIu+u1Y/Fle
oBu0xwOnz1U6Pvh3NBE/hwpIxBLkDvCjwiP0gW4xPAC/keRalwVEkaaijP7aW1HE
XC2UPI7+mz7iu5IPv6VmqqD8bbWV4WAmVLgj/Ns2mVDiJNmaffR2NZibplt1umSj
M6Fh9eZxnoiElU0dH/2fIvC1clLWQB5nI43PM9khi1vPY6w0O8XJtKaeoI0AE/fo
ZxClX78jshMkCYraIV860C644/5UovkzXrULVU+AT8bu+AvC4noLkTgUBm0NNhmi
mlLvsGSDQRM7OtNnJV1Zrs0M9ZR+LYw6BBshkCA23I/nH4MUzNH6EXh59xrtepdr
sZuSKxCydn/EOldlkG42V751AspgWnjWhPPV28+icx0neFrFbXRt7qiqrLzB88FV
67+xKHefxbgPw0QopSHbFDDDKv+phpj9sZeYF5TYtIbSnh8B3a8S0pKZNuJUpW6f
9mHkLal0LQN54wP0hgvTZhymM7XsAjpsSZlQft5AgEv+zJDHcimeR9v9/TW3IcD+
qoe9jruH9oAzA5UUM0NEcASus61BIVtNKZUzebyx8Z001sibr9Z7WcaEctsOqUfQ
MQOHA4iiHugGcPjuxiz/6UR6ZIMuAVZoxEA29A8bkJO7j7jScWBzEByteTLGW8I4
aGoCs5TkCr3we97Q3XDxijLHr8jEj+FArXNmMi5vICqn6deY+JG6tpy3m+YfASOB
DGBW72ElAldxvmn6Y0ePFzSYHCusCE4N1Wiy1R3+HCZS2suOI5mmnCVJcOH5icC2
HUirRhj/TNhe94foz7MUpKHWA204Ho1usVFQJ8XJz2P+5ZEdgsf4S9mTdBdJvyU8
CVAm4VedcBmWYA3TTBwCgRFdloXjRLf3ilSD8/1+AiOzAjJL/PHZ7vdDub8YZMoz
C9ytrlwZ5rz+hy8iC2qzEu9OO4xwM4SJMRNgDUV3Q0vRN1l0kXHlNM0QRuuLKOR0
OrHcsvZCYfZbBVp2Uwdwq9OmtXHz7/HhII7tcO8oEnC99DH1UWc5MENMmzNd8sEB
mUo2UNPQojqIFqn9kB7Q9ysuDjPIYOeQVQXpbnpn0Y0s5sCKKKuytPLNjvXSTZSz
PuQQ+IX/RXe37X+1I4uw+gPlx3ZtB11jUEoXIhtvoUy5TojL7zgqwkyINvZXmYT+
YZ/wP0BXGIZpw2Xe02XQZsJebFpVnirBOLBYQEFpMQ75O4ydvZBrnaKXUN9DADmp
FKLgrIZdw/23jd6Cig+S4J38mH8yH1IlLjfMarZroSGKL4Cy4ig7aWuRqm04Mtro
l6YnyctTNIAeNs8IPpAbHZerFk5xxa12YUnhJzwhSAVcM/hFJuoxho6I3jxz8est
xsOWCUQcj0QMz/SxB8MkP9c9lUswfvZhCgFTyjDrSB8h9RXug9aStQ0do5IBov9l
nEqmyvII6vS43u+1DAFmhPZeJm4WoVmQh4G5dQGhl8FIlEltfMG0CGkPLiXEoWDy
LGmHF9zkEemCJmPl7IO00DDiwQI9oiUVabOWVDNvyNiLHdeK4kw7L0+SVJUaPDcw
3ZxGNq/TDxVaofP5zVVwhER9Fy47Xs5t+XWIteWT5y2lwIrrr/AtpdPZ61VA5mWB
SnfYjgKBauHkffsoXQVklcFpOse2V1vq522+1HgZfme8iEMJp/G9WfR3u4ootX2H
paqThqqLNvKg1Tt40T63bw==
`protect END_PROTECTED
