`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wgk2zU2gdZx8GWt0jXbSE1/ezYK/qMgmvLLE1VvqEgiXsYetKz8SqfTcyhRoQkJJ
jPGbtyktj4ak7UjtFZkBkyEkLMigLto7ZeYxqvZb6hdBuRTNibhj3KXf3OxNMHgf
aAITVm1vTFjGqkbFCOu4PW/F6cWv5zLOHvHGmUSkcXNqhnOHxm/IaK3jxwF0ppop
ZjUqPN8vj0LDuB3fECgdYmhIF0Womyu6pynzq8SU1ZJkr/lwwDcoDhHrnDnfDiFb
7SVvHGWxuri95gxc1Vd77Eyvwmrnsd3rBUuv8b3f1seI2Lb8zx+VbkT0TNYIuzdx
7MshbmLzA/PH2qXwK54IZilx6u1aCwP+nwaRbLYKep9FlB4x1Pyf14eTWuwwIoLl
Uq53pKFnzO6BhsaR8lMIahFBVGCKi0TGOc0ZwygSt6Ad/AZV8Sz/70SUtU+SiHAi
zR7a74WBtvsZgSQD14B0s2B5DRZACW8PGVxjGf6KHa3cQAY0d0/7nNa1MONxOZME
jVR3s+GNqCCZ58HGlnFgPB8jQRiuZb2HeWp+DtPlvACNZ1jYd7njp6czRIngDQ7x
WtZ3eHtlV/KnOJP0NwVcGIMT3Fut4EuEO1PNv5p0PN2mdzEVKTwYrzjqNNSzjyor
elXoUG0HC1iinspeWXNHDdWl8SE0qnDdgof8ZKsHDNZ7kM73ugURQRH/nKeIjrQZ
ClKghSC+QLS3OFaN42aK8oHsgQfgoEoD7KwwpSBRUncNyIYu4lHpCmJLxrH1CFEF
sBY4sg/LFhk6tiyh2Wwi1g==
`protect END_PROTECTED
