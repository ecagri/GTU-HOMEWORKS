`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K00G5T4QLfLV9gBBEqV1rQCIkavMyRZogMaBCYEc6wG7W3CVIU17GLJ3KH5rPTQp
P2cAB5ve1byyC23O5APmcPFNcitncGT2SzGYK31E2bwi/1dy83K5NJLbWKqK8rtY
BTRQmboQapGWzNm20atAGyQHqJcE3Dltbj9gd6oUIQZLGtpG7hM5UiHVHAh/6RvU
a7lqdhDR2bGUkx8kv6PMCtc5DJQwnGugbNL/GMH6qbSQnAJ2W9TWqFGz8X4Ljn8X
c7BXE2Vptn/b8IOM67H1LqPYjZwidpWsJd+SueS/6dI/V86izp9foXCVhu/Xuv68
ILDzcFsKknOfWqJFLzltxij4BbhH7r3K+CaUm6DieaH7iGIFjaIJc8INxZverVzj
X2KKj5R9wBHZ7qOkawlp5DxrfoaTa8JvisrM3HItvmWQYvBw6yfK6ZPXweLZF2Re
BUiSJOQrpFTq2qf/SLXFfYs0vVsg/qvMauMGDQ3iCsEdrRwDFG0onnSmv708xRYi
2CWfo6hIpDTu756Nw+wYS2RTC2WkpXBXzz/5ULR/9qzNsaCTudNCgaUyam0EBMcH
gELrkN3ncy0adj9jTa2Si1/dM/GJdZcirID+SYtTshtDQIPSelmJW2hzDimHsrPv
VdnkVX6rJanWvHvjczHCh8TqSDlBnPuyFGbbBAwGn+TKqTM9XPXiaKB/7sf9imOA
wJblI3sHm3HibsIRLP/N1nRsZh/MTsLs5cjfETm5pvYpyq64wnejM6mCYMOshxeD
fNJb46WJfkPEcdv6O/W18uZ/Us/w/dXlJfPiRQF+Wj7pzQb/pg8PyZi7MFi7N02t
o2znRdT7S+UF2DpZhN2OJA==
`protect END_PROTECTED
