`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7QTCbZVGSy5vCwi8ktyxyfv63WELqsMy9N+PjvStMdiwrrHNJ2hT48hsBQuOBmbJ
WBnPHQarZ8f7GITSiZRAfbuIstM6qnJDvBvZd/AUrCihkSlj7jgQSd/si+nUXfvR
XQUtKxet4sFpvBWt7Uv8OhkMdTVOgWl2fo1SKRJBg2zupIlyXWT/LW4NOvolZ2Es
aYbB7ISaWUWXGYst7MnGlYVk8mro9/nep9aOroYATNo57oD+5U1xosKAVr+3IFPg
yEKz+4C/DpcOq21tbMTaBd1xu91rzdbm2r5diEPFgaXSbXcGwWSrhDC39EwQx92g
I7VyrlQKFBFTplRd3uYr/ryY2srVE1PmmhN3Uz0kI3qfwkzrpfnuEjm55rcXcdy3
daan3dlcTTu8JT2HWPK0iO05n26KJrq95GZ9tqxr3/TUFi32sXWLZSwPG5WuwS+l
UWaMyZ9XwFMk3uzpm3R5mItqkkF4qhO1aE5Ofi+esdXLY8rF4cUv22QN1D4yxVyX
85V5RnLZZpFncTcK7KyfmODJFH4caAuubg/v8MmwSkpeUzqlvCU9+oicZDBU9unc
6mfXZSuaqEjz1CjPwxCK0Nmd6j+J8JO4dKzqaQi/Vg/9pnp+qsxXFoXcJCwZp7TG
Ewkm2k+dzIKyH8TwyrRkXKq/GwuQ5zQIijTSnPzLE2cqDv4Ic2403fXIKaIlU4Ae
GC4uDCA9sgVBafafyxvNLC1Z00aq2ov7BzWJjv3+JOt6Z9h8ZY9mFk9PjwZ/+t46
vC6TRweI70cqS/SI0nnD9XgFiVlPMd0ginvPTxFclQ7ljIIoZ3KmF6FKVxEvCScU
q0/XVkuHvCFbmktiAs8VJxoK3EAks/cLtL11sn2v0MMwhnqYXyiwL/YjceoyFy5n
yER08Z4o5AiqtTSL62nImzRRK052NP10BGDrLhUo9FsaJcZaLnQjgUj3tGvXMooR
0+cHT3aSeQ+UYp0daEp7kPNEtaDsUJ8FMCY/36p2Taop7AR0FGNCPTb7dGxxWtA1
ecZsmeW9f1uUbmfdfpoWaEULsRZBkQVIDx098vVQJbbDoHc3Wi5ypzbQ2Ff+4IcY
Me+w+2agB8YqIySTbXDeahZylkk+ArcBwPZEX3VM/bmzQOYspr8OgGplopZP+e+I
yH+MM+Ijqg+RniNeI8DUs6DujFOfIKXXkd4pr09Z6Fzm+ucZXqKh8U+mnpi5IgNw
EQSDCBMYLb0t9xy7uezAfWybb2F0uQwqjLnN0WeDRuUBQqleBky7fekwPsjVKEu/
u1E8V+5wmatxkSuXIWc4dhB3sAiKxR0D8zmIczfUsU8k/8P7U8lq0bcJAy5lZg99
jxAyzfZ9YYkZejUukDVvNLnSRSsFGJneOVxyEf4Xj2lfL7cWvKGWaAZNVB7/AUsk
3zgW4evNwdArT/6y3pDEZO1Ut8xO6zkbv5aFQrPAesPsR7QXdpmuc+ewcu+RdyD7
LT7E2aJmHmOELP1tXuNEZmS6QRncod8rOOmYfxg8JGe51fMGsguneE0tXFQbIMQo
KPBk6/Rhjh2KLs/SNdC+s7UNrYiY7Xmwx062egmhufLzXTsi3orJBGMhMcZDvZtP
M4af3JicgzkBdGTH9nyMptl3Je6dcjQLJviYlijpZXcGHzEVDmYfHiWoYFL0l1oc
SjEvTTP1XFseglPCZ/1geTPLomLYd2zmCDG/BIxpgPpNaHUPekSz41FRO8hub8zf
35FxnIBhQYx1U3HU4N87QUnuJabe7Syu2zQI/Rw+ShCdZP30EWts0EsIK/+6S/iO
Hcfyk0CEjUwV9iMSVnc+q8WPgF5LCavvYce+SBOoWtNKKTvjVBiZ9xlxvHThc0+B
7zJZjBrqFAOpYm2KXuOmz4IJiPQx5M1fGOEOhiAW6Z+ZoLNvC/WIqEnDmQARWjyJ
WnzZofgPaXbpA0mcZDGyzLIcGiYUw1GPzkNEw53+wL/KuVrmHZxcjdpJXhPPopeS
k22rDQi5lWU338QAhx1NiQefIQgjgQiGzZe44SnxupPI72VfXGAPkUIysg7OBw6n
M8gllguBu7LH/Q+p7h8We5/efyuX2anKmmgJOnpOFuJRBUMO3BD+Jdap/WG2bJod
X0U1eQ5edP/keSxLAA94k6qt58zdS4Xv7V+E7ijst1DJVSqK3wcITlYE+wrMUwRW
fqZuKSn0y2EULbuw2gGy7qMzyjJU4L5edJbm2+MHsKzXg68xrVJK7GPnXJomu9kH
rY0dNjfvqQ6yfbDyfOaQV5AisNqraXYwKLtX7Tb1C9MDq9nIqDtC4zZjCuTJtCsH
7xf39WrhoFhkAJKaUOCe2hPzKhknj3iDq6bkf3Omc/6V/jgRWkSnJoIcst0MrMpa
xu0pV3GQvJrmuBn+/b+oUqd+kUkDRqWEvgBUetl7MHQIx5MYwLcIxVJpIyaBtcNP
adCha8x8ihCoRIuerb4PYXhcLFqG8cews5PdE8pJaqY8TzLRSfGMYwbFJ92GHa9i
yGNBVoTJnJoZmsquJHiR2FVdgKMQz+IKSXquqK/c9tKEQMhFnzNXtJ/ZzwST97EC
y0vDSAYOJHPoxcNaJCq3k+As9l59SsNXpucqv8u9CNuyFOWqhaNXMQImQhGUNwiJ
PWHOipVQVYdbObbobU91oeWmDxvvcgrmHFDM0t4Sw+jN23j5rQKnpCNWqPaoKMVq
UTnq/p99frRTxqVLybqLABvjIWbkLVJQEGULp1oRwXo43MqRfS1t7R1/DQp/Nptn
dhpeGRt2h2Wx+a+YJuV1ccHxEOENljCp1lqTBTIRF804fw4G9c24qx0HQPKhxdpY
bYxbxVJ54DpJfqmnjHhnIH7vnL2jhjLehsx91k6g9bAouvtpx8thiqjzsRr7Jwzn
skn9iclu8nwrn5l9cOsraCBqNLbSvbsr92KHys0CzskjCA+mTvGK+YWgYuXUwtlM
FujC2MFoP+Zn32ZQsBib1Z+rUAIMU+PxWFGw7aiD9Ma8YZCvBu+HKB30jisktayk
iPHTcndH9bApoLwBjT8zaLfZRBR6tJumTEBW0bcUsVyRS6tfk9jRPxXhu9EH4Icy
CL+8Sau78vcpRVWzO9YbYLJVM7sRMKcZn02BejQO6oq8kgYNPBHL2GMgarNJii0Z
kn8UQbEMERKMN5+WtZgXH90oy09aMBqyn34rILCEbGcVdMElePjv4lNC/ts0Lb4F
ohcu02S+v2JlvrA3SuWk2d0k4bTnp+Qxj+Y6bjuki6xb+nsgJuhbk6OXqwJZAFV3
JhLy4smtC4BBOze+gFKA2uWMNP7ief8Dn1ZBATvNu7qIbZLtFnkt6UOv8IeErp8+
qkDozT7yVKk0ongPYqV5MrvqJtTDCzkoVM/MICf8CansQD7Sw883nB4xmexh7WNs
RGah7i8I3pb4Wu7kVydnyNO1zD2coV4t9reWg/zgwV/KShiC/Ani5BqjdQwLFjzL
FLN1K7wlihm8FBHjvnmZSEUP21Q5ZOnP/zevYp1RztPnappxafwQ4dGAV/jsUC9M
w9h0dtOMYWkbBL1UxDHlsFDZCaURZw6iJf930qF6wUbtCp1NvbrKC8BxycKP1PFt
a1Zx0f1TuUfNkkD1oJRJ678Eprz7dCzj3KwHhLGQwBcXlfBZ/ViBKpzhdO4IOpA7
RiOq1LCxM+Yae6pcvG8/q/lMzBh5xaDyqFP4BZL/asOSCQJ7kTDzGY+TAlw6CjEv
fiLtoqOX+1XsnGjmFRkZT0TBtzW7flY9ItZx9u05wTcvNLoZhoB14He1YsZeUNZo
XJfeoRBZt9gjcvENgZzyCti1iTlBw/q1H7qVECrG7BOwG+30gxaLtJ85tlckuD0S
i5mHpe0dxUD5c473mjeREXezBdlfuBjnHV16KeJlunxsFkTlbRPhc8ntKz93Bpif
8OJdcwBJdhNYwFUrL+/i/TW4pgX/INU71J1CV7ALYmrN9xa2IFYmFUJ2l1SvFp94
y0GWC5CvAyVdtmHc8095EnUbM8Mnwtb0jMlV7VhKnL80WadOMYzT7SVirvUsTRI9
ggxlaf3Qfq0O2NDwrXRjk2l/YaFYctvRVZ8kvhiWAJP4eJ0qi9xz3C//LofZcmU6
lF87XN+MKZ48BvaFpmdxAwiSihkkLz6vX1Kg5Sb6kd1o9t1PnBN5vwlBiGhkT8d0
FQqa3Nq68P9k217JnICT6j15/sAKz65THrKbPm2RQcFt/XC3cDJ2F4qMSr7SnWtT
yTy5BIrVTvMca9cnE41CCSyK/bHF+YmyIZQOUMYnxZLvD00xcJSHTX72kV9zld7n
`protect END_PROTECTED
