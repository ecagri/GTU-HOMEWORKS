`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RPdbtF/RiQXzCcLunD37i+2ldrhnAOWX9oMcw+0/G1VduGOjlqiaFoEbW4xupmNR
eLqVwmb4fZlFip2j+WUK28qzl+onx3aAM1HqwR2OsSZR2KgI1mOLTnw/aErwPF9Y
SzVWejw7e+idQ3LuqzWvmOPBzQ3NSj3I9im4aGb4vvEI9gZT0osxa8H6KS+qBIoT
/EokGnJRg48KTNBx4HEy3HrHXJkHOoQav41I24J8orWcQnuDBrbbzC4MyeK8JC3k
B1hRCxo6NHnOLdwa/cW9jFPOlLwWhyPAMrIofuVZgZDtQAp+4CxPKUeIQPwS2kH+
flIS97Hq6HIOwYa/7aGLBAKL8PItUn67kjLK77Ue0Pm/hXrmFWsrWqK4s8ygCtSZ
n4/8/5pugj4pXuJLyP81OrP4IbHMKJIopkRPl5q3qJa13SZIE2Jle9WgNk2GMbHl
HjhXQbypgl0OplqN53NhNSHIOVLxYV2teHJ6f31WPo+tII2rihakFNkDUSikCCpX
rrIqUzI+keIEAUOWaaj/g56k0bXlnvmw4rxmGAwnMQKxNeeJ4u5mvlxOqUGAQV2b
+aUiLilZ03w5mLAUyya4uaKlpkRbP2xq7c78BoelFUEj1Q9qtH7vizKi05QWvl6q
bSWvCxFSvXCSzM+5XR+xmU9Hq335XwrWqzRpx3H8CT89/WGp+76nFO6WMZx8EyNM
ACEA/gSCYWXfQGfz4gZgur/B5jirZU03nPLOWVMjJjBozDBI+3kOADIK5+J1gfIX
SqWEkrCns8kIRnwNfxBaWAgKBDMHyMNVj0KE5IFrwd8pt5Lpv4LWwzRvmWGQbJMK
`protect END_PROTECTED
