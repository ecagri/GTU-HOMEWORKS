`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OD+s2J/OlfrpH25t4hY9XvLGGsxteKDgixQeZ+A7aXKJ+yK1UASOJFgFrz064J4A
G1F3RBSzfQZfbI4q2FYx5A+2VvQ8g95eDTwdLZfSxpsL4+38JCw/RrR0Cn4QPFC1
mbzzQt+wrTMfwXx5d4g724sm5ThfN5tTqz8Zx1/G0nkdIA9APO69gJ4Yv5qGrBRW
nr0amgQNcH3iYkCifniJ6MtUYMj2ceF0uk7cou7MbBbY9xF1nAkOC7JPqmX+w2qY
/qf/J7ORV1ctj1ff5bczet9hmiiSPMsC5P4EVhzCLqxDnjaCmJDvBjYgIEbb/W3t
H7fiJflZjMYXeB8r44N1FsDRVwZd3eB094gP9h5Y6Tyzo6+qIKAWuLomldt8WS6T
s0mY2/gZy6j36xoV3arvKn1pzEj8x3d00LG7Le7038k=
`protect END_PROTECTED
