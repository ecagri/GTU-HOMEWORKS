`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CT+YhPIMLUBm8Lku/UA+6/swb5Ig0/S7zoPMY2Q3bHIyxusrBWJ977T8iJAns+As
YxSnf6PTlicj7+GUv9c3l5148vYHCEbfFQ9vUMS5LF1xtgFBQCgnd4XOEpgcjA5k
dg3sRAlQZW4Ajt4jHMGL82YSxVvkJcvZNxcCifpDYXCvsgYcjSYEURFoRyySTPq6
J458boBhGBWglLVYBohVs0tdZbmpPBF9Z6yxXA+HJYqOwZAx9Hg7ClIbkhyvzTv0
+wYWc9fPeyU3W8lxaqh8Y9E75in5ctcDfKTDjahwwWO5gqh6wacFfdiLzCuWfLIx
Ok7SFNkO/rNBey5A3Hoh3McZKZ18vLBr7wLppKSD9ect8ZYrrDTOJY5DubUb//vG
RAYPFba30OSitTAGHAzJYLUftydOSR4kJlgxJQQDzEEdUsd8kP3HLYSiwNGaCCs5
cOWlDIvtgxo2JFR8KFq3zT8E6rJU694gkRFiqX+XD7A=
`protect END_PROTECTED
