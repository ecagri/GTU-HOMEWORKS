`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o/QLdMkwZ4M1YrDof8fr4rox0X4Yi3tYfDPOWqpaG/joba8RA5WAyD6kMJMDKkoG
zVL+1W2YxwI9Tx7f1j3qcqiAvUaYxzKnmv+uFK1fyg5xDMPhXvQqIduFDLfzsB7G
woli87ezOeaqOE/G7AnkoQH/TnUr6l+nrH5A3cofhcIWoaNvJjx7ttqsRt+Fssxc
SP4og/chI9UFNMNHZH+PG/+fSMOtGtWkQUJr+DOr2dZgRohMT//Z4P4EG28i0kFw
bnhyaRzynlnKuQzxeuY7sdARFkaxgn6EK0GsqHYtmU5PYVH0lPKKEuuladE612+F
LGoPoD9hjvg3dcfsgW8F4MVyB/M3JGKA8UOSpEVRTDGbhlXbWjJHOiwVj/WK5Q6F
rHukBsYNN7vczT8IRZPofhtWZb4Hu+ix0h+DJJzZdBRlU4FWaLNWRyrjcWwlEpiz
n/GuxXm8i6jdGU2LEjeZB+AJiQ37U0qMtug0u+E8bQehUz/CmknBebnnUnHmYCxx
puI4B4CX2dO73i18kGY0OSnvW3K2pPJFN8hWqiRaOwGqNTcck1P13XkIO+KOE3SN
9+s/Qi/CCwvh+eD2PB47lnw0JYn00f05IbM/ACFVnOW3Mrng8JyIPX++ZIvKdMJ9
T/h3Sc2pKokLZORzBQ84rI63DziCpcWQe/NHm2MtK2NEETSV/1/gUJenOPF2U5Ka
psu5JFXlwDJpBd3kX81eQ4jNkLE72Ha92hCvAezHNyK/qiDjJ9myCvFJSVGho3Uz
rHiZ/wE3kIz7eqUuvo1UzKQ6/pTcmcWQqLSHR0gPF7tnKO3m6tyTzWsjoVk1M/S/
Sb4va1G8Tz2g8s9CS0BCodM6XEZ8LPrnjF0Q/6Ti8vXLMUKrn4xnYAf6KjmqAKwF
MoltBgSBD507NX90+YKYv9Xe4OgxXErxpmm9rh2ILkDGGLJ/fj9KKn74R9qEdjPB
c1n6n95FkgTgVBX9lw5Nh2NzoJXkpf0bH4Q/xe4t2kUZwDUbGh0bKKli5rsEmOtq
EOc0yfZTy26E3KxjsX5M5HhdZqm23kygIk1kJ6B20l4PoabzdrSx8jltzHtDP3GS
hgrXNlL6raCwOjnWf2rt5pRKNKptL+du5hCTCKYi+gWS9Gg97dftvE+RkPLNYrmk
V1l+zO910Z8aFsQFYlq+JvAa9p8l14FsDEswANNBInXiDT5lT9b1W/uccwI7/e9f
p9Bl4UyEzt0TG3bpJ79dylKOthKeONuBP6H06WI6mBz5UeB3MoT7/0m0WfBkA3qE
NpKy9rq3L7Hk1G8axAhCHsmQmTxjWhVstSyNUkQHEYwq+Oo50090RnPKEuVby3Ms
nWSNfXn7zagDZ2WIRI8j9JgssL8i/f+M4UXaVbx8cY9BvnclQMQ1cNTdPifaIi2g
WAsH0iEyfqGvSbkw2B1+DcLgQ+jzHzUKh00U+mliuRsGejk3g4xpCWvUyRxJ3H1B
J11nUGDU2llFaSn0MvvlogpDB/15teUDIT4MaCEebIrpPPL8nF9Wx7LTONHCui6R
t41WQij4hX+Hv7SQmvA3xoCmMkg2pcy7uDv1rku+q4Fn7QLBtwT1C4lBIruMmOa9
ldp7FjblCcDMqlhZLlfz2yfosFuvEnaj1pzwc9Tu676YXgSr9wJSfh7lgehjfEuV
7FrrSt/ovc3DmeXSIj298KXt5WM3+gw6ctbfFYXShlegk+wRUqhzB7BpTtzxx41G
GHPz9dLzxDHyqgm3ALREqEuKcyBrKQYxReyP0zWkkY0WHm9Mk0o7RlZV23O45viv
AP0tKrdIBae8QjD3dYAdvsX34UIA/N0OaymcFnKUQl7rwBxBE037zVgzuikGwVPL
6vdfhFjeL/xfTrwUUeJjAqgYJUlzNcyq+UERw7ud5To5FrTca5uqq1/E/nqFz9C7
hmczJhd68ra/jpa7/cLBeSvbYPw6eUylPZYOxjSw1lMlPwOvkE0tiwG9Vx1S+aVF
qTwi829eRobwdXVWnoTncM+ZtRQCfa8B1U+Ghn/S/1t46lFHoCeNO30Aivv2mthV
9ZpPElOqjiDiW4u2MA+deKjk9iNLNyIJflK6h/c7x81G22NsCVs2wPawEXpXFN9O
anL+KGzD/IIkmFSkkhRhaMhEf80C8mE1Ra4QowH0fBX0vWPhJMlmDa2p//6XA6Dy
MPpFmLeJunkdaNOtbCcEiOH7lsWPBeTE+NwX2EGMJJFMhmglS++ilvra9drNbIl+
f6RmxY1nXe7CpZ4PINvthFBjS0cKoPIBjKa5pno1BFc+0d2FWHr38y1dG3joftUJ
6zA5QU+at19O2KLSErHUvgXrE72uz2ouPsH55XAueMOhrkFNGo/rujtRakDFTtQq
Ekv0/UmdFCd8o7Lv9qhOaeN2ELuy50FcjM7syvyNPShmnstoxu8o99y53A5IAslM
DUWBBAdy8KdvQw2KCIB4zT8Qpfnu6Gtm5JAB04KmBYcmwQX8jzK4EbH6UB6jD4O+
38okkQecPUsrLIKrBPVDK59HsUqFKtKaGVKaODeKBNCCKhLz0wRzyLGsy0BRaLVE
g6Zd4ZoityeBuQZt8jg2bgnnq/8J2WpNtQonQtN329ZRif2gvi1+kQRnN/MCP1G0
nFYQ387Fgf6u9haKOtaP2IegdMybimT68jrQDioWkaUx2Gb36gGVVViHt91uVvjb
isSB69DYXRj8HxMkW8rCZxadxnSm8yp0tCciUJom7MUD9hF+HmQQdKyrQHlh2mIw
YbRkG8aWj/C0d884A7npJ8zI/8WH3YK+vhO/M2V4usV1KubHqKDDuFPSZTNmhqBd
EvFtOoP0T2IbMTxbrtj6fStszT0ESHR+Zj0bfrXmTag1sLP04BcNH+yyp3KtiTNG
LqTXPT2QKRLIGeZIow+XL35WY57pB3MP4SvNK6VvQ/BQR1mIvRy9FpM9PPnFYZ6v
PROpCoESyQCgkftqupISLQ==
`protect END_PROTECTED
