`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ycuCzFi2pRqBOlmeEtuqZlecw/LPXe3DPG/DVvYTsgtTZ/EZexhsYECp+qIBYrkj
NIZ8ZQQam8GV3JBfJIOokJ9U7mPnclBmMGwlRuNg8QgcPTFWJaLLIKdOjOxELvz1
3OJfIy6FZZEEaObos9kB+EOjr0d/X1UMD4CSjuB8zQHuCSG45SAU5+/9VGpd2AsC
OqdoNsjCbrZK7s09T9HwcuFsAeP3KFeSw3jnnz9Mik4ByPebn72PKJEBNBnrdKEh
6VdQRGzQFuNuGiL5PHh8R+AQk4kWYYRteQ6jIx5p0vJqa7krtfEQ//HxyUR0WTSU
GpcUY9Da74WBZYV1kJu8zPaoc4hKuJrUUyHyXIJq8UVsgbkIPaKbktMonGrjs6VR
FsLOm2G/DEsuFpTuzhfsx4E/CzrCc7lUfctA60Jsad+1mD+h2RK3MFrC+k2n7nju
zSCBAQ+IiiKt1MYEKVSWpeXQ4GF2CbIksNRMZutaX7YEF3ebpCRuFTSAtc+vOUN9
BwcRQRDmH7ced6HzILOphRon/2+9QuFtlBnUfiYPao5VEXzRtW8akcS/wa4hQbN1
b8dGPbKs0sEOpZcdb+bTaxO6czXvpaaIR0TLCUPktjqJxdOjLGV4NRWa/PHM9pKO
a2xaIWBiUZnUTFux8rnFczvhtd9nBI5B/VTE1gxydkB2IOwsNsocTUo0ARxtZIGa
7f7fNMs5DCn0C1R7kSs+nIBy0nI4c+RrO8MVM15FNoUgbyViuPHCghVod6vml0sa
4sjLYBSPHFXxJqXTfcS6uXA7kkvIZdMJbS7cspXGaA2rnH2z602JpJBQiJmqbMky
cVqGHvJQ8+SRIUb7DJ95Wvz8mu/BTfCJDQi9p/Pb1MR3W3vDeRsq4VNOpd1X6FGu
Z18FQdvZr2qZbS01xbq1a+4amyccdS/SStMj3qtrw17Y0x331XgKSe56hwKlAQ99
cr38JxgjpYjwny3VT/+DXwA/p+f0gZNer8eSwjoHpAINnbVA9byUh5fZ4rCYFGnC
GuLGtraKU8rR0p+bfC9XNHcE8fGhQ2O0kb3rQTJvcmigHytzKjQpgWTv378vhe0r
PL0eHG5RTMSj7Asvc74hKeBKvwAQXPE3QmNzHyjuj5Rtuj1Twqt5Vut/+VM9+v6R
GaYMGQx1kOIlh0MIUiOt2msRnWxHhr9j/AzFsFmFnTWnxuTPBJj2eRwlc9LgLUJq
m8emH4UpaYeI9sK+b7o+G/5FJGk7ikVfvT76aE6298f3V9ulDj9zP/MoR5NT6Tey
hlQ/RUda3Wzufj6HfjQWKwRk8S3zQw9AR/kXHP+KXH+X+0FhRqeS6pft9WaV19+8
4ZzZfKxPRDOmKGWPFOFED1ej8PoQXalH/0G9b/YiQXNQ6iEUjITD7A7ertqRqOo2
Z0Ri49RI7sXEeK4RuR4fgeY7yRJIdlNzNz0NqRuf7xkEvvqjkhOrdn4ZLecwGYwb
uUFd+zAFcg33BZygBKXzw508CxOH6oYQ4YbTU/Q6q3at2ND4FCtYmpmhSsbiuKVA
w2mt2zLnOaoNCpuu9Gdn8a9krmw7ogXf8pYeXQScm8upNKyokklUgztcSBPNNWE/
6q4yJ86t+Fz/r2xOns1qTdYn4q/1yQXjQNflJiRNvTRyauupANqIIqnJqBP08Ep/
5GMs8iUnboSgvdCyWx04V+lhwHqxLSNp6lIDq3r51QumnCYRfFMu/EoNXteY4+87
LGl1IuyvSJ7ovDkc9J78GejZccTjCeN/1TnbJdz/XKwBUEIJWj/GGd+F5E1cab5+
WVrMEsvsIYkBKV7njzjpMDaPxnPmkDD7s9uRV4Shpj1UoflP4/KYLKQOWmEGE6fW
zk0+4XMeBKZU4sqIoK6Ruo17trnqfrCbPNvhhDrcA33JqtOOa/1OIAQrTRNZre66
r9gIbqBp3uauOMw9LM3Nw84fAF5TxvbExOPqsNSclafIb8zUkDALiIQc7UlUIQN4
tJK0/9aU0nfBPPFYlgsamyn+NKEE/NYKpSbIFxSuvF1fJfhKAWMIzp7/InHyjvIa
42tJbPesE9cknv4ZgvhWG417ywRxLbTniIIMtNQr+7yI/oqU396wbgvIyqk43Lys
Td6o5UbytFLNIEZkmrNgHPAK9pXQN7NvzSWixR6m4nBbPOo7qxigQm7jsGDzMUZk
T6hZBnKeo6fY6eebbqyFAET3BysSO20YcKqeZ4zOGTaSGA7RtQr8g7WE/bWDTaik
U38Ney9J4c4Vqz7/dq+f5tiS3iHB54vOJESaBUSxwyrZnpy8W35+bVAqF6+S5dfj
oLqUT7EcrCZs1fm8fF3MPwVYkRvVIaFk/K952ZH4KXDcoJ3SzEqDWLM8D3hKNSft
0XaU2wY2bzRDKtCf2G5Yn/AvOb+DN6CqZvZue06R5BnMTZ/uec6DNmD2nSkB3w0m
Kmt8cLO9Dt9ezgp5ZK/n2n32Zbvpo81p1o0k2WfK12NZKsKSS8Mx3sZYkeW6Xp31
Gx+FedcHg6hE/HfjWCFxrSeF9T+7v08KGhDG4lm45c4Anw6ztWX0t1jApXBNzZsc
/pl6ni99yPY5QvqWMM9Rifik4WtRp/NvYvnp20MyaLl0sO9vsFQVPmlzozoat8cD
X8Y1ADrC0djiT8SP0TKLKVRTKKKhrGJ7OjmKtPqRohX69ag/trdG2Gtn43EG4aQb
nisLeCjHwX3ycjPCUISe1v37tvaf2PuGsLlGWsojvcWHNDBbYiXw+gCPR4R7kTRK
TeT1UOZyxLQrQNOdpSjq4yRSSD/EElHMcYTTZM99UbTCVyIYWuoZMjLLmufrabnw
MURi1Y0KNSDygDyTmfTwDJOAuYknCUG9z+MjkMduImYFfCl9IJBeOYHCzxT65TWU
umwjWH9Fj/TaVTagzPHsiPgv9jMlfvlEawsKIPDrRq8I9YkF7Jr/B+hsyWzT/F4x
ckfclrSEFUx/6kL62bKMMlj5UGOtCyzN/argy4Z6HafZrWFu2chdxWVYacE54JtS
G8a+xN+DuhlsdR2Fh0yj3JL0cBpFuhxjRuz57ms//aNRRSvbB2LNn7o182+rf9Ba
/IlFcq+PO2VvX+7Tc1Zgn/34SIV94rcyQ1QbPm4mLFvQWQtOl3OsFao6iKRkIzTJ
bnRrGLVasEpb1Zt6B87ygD6yTRnc2qW6+NwzY+enofRkwCFGQvvgIQiv3KxlQTic
i1BH9EwykgAVfC46uLXEJm7XrbhlGDPxo/28h7mzjFYnHA5nhm8LMr+VyakGp5T2
lAsZTI4h4sjBzF7vIB3dyA8FGnGPsOXlq1sJH/Pque0iZ+Ifkx+Oj53zqF2kQjK7
mLwArfZcZXZZgQhNxrzvY2CAK2qxVPY4yzRepyyh95E9kxxe1ECcMTBhRd8KqlZd
hv5ph0G2Of7bATHWqfQ+L05hn9bqafG0jogdgLxiGE5OOUgHh6Ctc8Qwk4ppQuAP
vkxKLXfYdPPbcvqizp7XKvBiOIdnWPJw/RPRPgn24F5FhGI3JzFVx9Ci4kWVuBAp
dphijxKv5JPdUOwUT1xZPlx99XeDIUe2Ob0mFfTkhYhK2lIUeggpvzEJtwssb/Un
ONX5S5B8Gnt69NGeJ2Cs3u1vTNQKpbzOJG/HVTQJEFplSGIqbI1x23XX9jMrQYhY
78Ef+RznrxX5uW8r564Suo0RnzcIsN9E+c42HJ7DcIA=
`protect END_PROTECTED
