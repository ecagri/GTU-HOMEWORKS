`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CRkd8KjqO5UvxY5gWr6oSOlnIN3rUGl0DK7NdZ4MNIqIeKs4U6UwRXo9TcUe09fI
aPVaJNVtApjrFrzanOB0AU9ukNUJblXwD1s74TfrWGwkC2SyvhbN0ZVAg4O2TrTb
Q2Cf8r9mztuMLYx8v3/tEhdIJpsftSB+kM9DZ+b/ALKxXULjfYPUPN4wP6QP3Xy2
DqK8sg+15UudIvar0mlpools0oIQXz++Qja50h3IimghRNgxmNz3ONU7z0W1rUoR
JfiZ+xFzAwFco/MxfzOtXs+UgrDs1VecgRJ0Y87A/lZDmuqq2o/AxVVDgrDaXKge
YWsU5ZUj/ZwPiViRroxO6tdVaqzkXjGJd0+Uh8PFc4WUGVNZoTBu1bOguG7UL4X8
K0Apk7dsREsIvO4GGQXn48OuG8dtGCcRlmOVTXmNDuH7TJF99tHz4TDLxXp79cMj
/r9YKFqNlRiEPLxUHTQr3ixoyKuENb29tJ2ggmfUQ3VktApj96qs7/ig1AXbw3Y8
fAxSycjsG2DsWjY7B0FZoho1/6ui47/w3VPtT5GEaTvFYO7bOnen79lvabo1GvGI
O+eqQZg+nqa3rPY1W/lug6fFoGI4ZEo6JI7H3Ex2/ucGb8mZGf+nJpfmR80Kg5UB
xzjJrD6ABf5SsWwWfxR2s021LXDsTbSQqIuAk+ZMLdTwncTUNYHSTcq7CERKp1C2
+U0sVwtGJkqXQVBViW8BVFWqTAj+yILNdyl5vri1Ly/oJSxeBd0f8uPm35koKdQu
nlOWwgi9ohklPueYdIXy2NyMfnPX1tNX+La+86CTfvqlvLWl4coVvJOJFHHoec6D
A/FILzKVgiPEcJj5WFJWnsL8m3pmEKkeA8tREtFEgCYGMac+8M3hpMWpVuNOwFIa
1zH6lNKoqqI6VdwMk+XAjF7rqjVnOahuQe7VG1IxV9RCOCdVZu/K8x9jY4t4lkVe
CLI4a4inoUkrQfFDI0xm4acunLOKXBPbgZGY88Bg4yjvH3W7N7g9109RnRP5nJ9H
x49oafih7VenY0rnvs4MAv9W4N9JrTOkG8bQI0NJdvb7bFWx3s838UuZ5wpXUiP6
Vi/0j4wQIbI/m2EC2NyOnNXwmxBXssKSrkvFR0OEUwIt1X/Ez3cgO4Drter2pZDz
kIY21C8XBZUmfTIdQkS05Lhb8+LyahskxEiMUwaIT2ZqSb8KtyehAvRxPcEDxO7u
1JoKtO1K1B1DV0Yh9mJQtH5Nqim2gaQLceY5ZnzXmOmS06XWTdN/DZ18JOpjGXw6
JjfieScT4WZwY2lZsmjoTEVS+gb5AFI1H10Pr8lQ7m13v3lAWkAbGpu4sMqXmmSp
RmfYVv/p2vsw1qHLAVCBAbcfyfWwS8ATAO5kVksFh9jqXBmPQMXqWydHfTVfiIfb
0i6//ZRNVxcc5xYPMCOBo/JRMv+lqeiMOnTosoVflpOhTFTwPdUZgprJATA/cy6K
bWInA6U1KyE1+CDthEyb0SgPcJwREVn7NiBis5XBnFDzv/xub3aRaFvgtuf91pOS
bP+sgdJiAP52QIo8sIuoi85rVxp2+Y9H9v2oyQUrVO4JhWahBZ6jE8HWqC9WgKJy
udC3xPCYm0rhSvcxw5tZcAjdyHttm5fbjjrlmKk0ubGE6j8HbBof98CvRGPhEaC+
ub5Eq+gxk0W2HD+rLJxfOTMcJYPvaasmu32Gj88uOswmhE9eVWReW9Xt+R6P4hO0
bk9HfmTjCY6MC4S3Ex/EVtsGUcA5v5hXAlsXP08AmGofQz/I0mYZkRb++UQ2Qmfk
DNQYhDdP/jwl9HV9l18l6YDzrbwQOyDvYwaCvsH8hcn0ozxW6Pw1d/9K8iyMq4JZ
ew0efd/R/RB5TQKvu3LQt4z9pR3L3KiJxmrGwGq3Blz3WrAEuXr0W1sa0zfaWzk0
1dnB8DclFNZlXGlH6bA8KEIXJHWqQqEdXwBAyHJTDATSK5JlNjY7kjfXmG0WePHp
zbairXIYHmHk60DRZ0jY2+ybDN//+hfuGuARIBv9/1zkQ7nC3yIX6pBBuzCW6lRm
AnmIGosKzdtANMMM1p40lTLfGlHBq5XbZcUFVQv16sidCmSqcJBqNCkVAS6/xxzw
xtc/637WiHfR/foDv6uewCMcUhKTZHTrwT3EXG3pvD1vwoN1NYrA0ObrxjGU4FiL
x4XEu6fwYvylHfFPfRk09WsgoernMHC5jfltR2AWgnrOIiB55C5cRLdVHRWpRuOx
C1IcSY+R1PeHIrJm5YIow3nSROOqKNL5PRC8FIbQ46gdRIlrWKOveTINYtLFEYAz
t5QuWm6JcfWTXIwnHmxtyHOiMvBlrtNoNW3F3rvGlW73gq+4FjzTpsoHxQZ3L/7W
LXn2Iwc68//Etdra0WcYlDIMfukzH4VVa3adLuOygO11n1QDVSJP5b4JFnhKUS5W
aYNUEpaPXvsy9LYrfOvQhw/AWre8UA+gYsLFDRICpdCK/M+nxf5A6VphhcF2uNYt
iYYYdckP8HPVD8bB2Ami2BljlASoQ2eY9lPKAp6qWnTDM3THoAbeu9L3MvPEahRG
BNSYDWpCBPIzQ3ioVWM5NlEbhbW0MWcsORWtUVr7GCSC376Fzu/9SdYzXsACbrSx
uw5ps8YimhbyhYVNa4Ds0B+oEDPKHJ/RPh8jDs61qJy7DeKIy9ZIibBrrRhLnxCk
jQCGYYTz+YD6W66SAlFvOahC0SsGKT8n56j4szZW5OmWWrsMUrZU3jP2HT95+xq5
4SLRjp6ZjGQryzZCu5yQ+g8CfFsc7YglmsoI9QLtYBWruBf6G7K89sRmGPNnGHc6
Zgq8FUktO6bEkagLwfPKz1JEOmJq7yRF4BsrKY3FgGgli1e0vOU+Es0xXLNzS/mg
01c+qARnwOLBmi47K0PvslzXlL1iet52vKl3oMYB1U9I5A7ntnAlt4mHx9qzESHc
YoCJ1wdSZyv6utQcbssAD+jTyrtqg8nQC5KbtoFbPky18icRbaf6uylx9cGyc7Be
1t3BTZvhGsnjetty6xdl1hNLCDBLPcGrvpHnrLWi9/fUY4M2x9pHTe3Ze/UVDEAA
hdstA320FWdt9F1Mcd2MOf3jG42Wk89YVxn9ngZJt2xA+ukvkmRLfXrkT24tUmLi
73jp4DnPzyc4nqdnNVxs+pwBQVtkQC1OqXIeUG7kwhdrN0DqGenXuawBuQlfRC46
nSG+SS3W9p7V1L6LN/rYsksFyyPvMnXhWEnBU09VtcSMZEGAoVyy+yMYtNYSIMVW
ENACtM8veKOjJfwYizJ92KmA299pEaYm2P/tm78kdgNewM91c9lyzN7uOIZ6+OKX
v8x0J3RcAeBV/owRoIX69dJQzqTuxEOoI/7IEoxj87PRqjkv/cE47pG+clZE/joY
brGJeEx611P0ZSxIkstWDbn6Yjmwky2/SAvHa3QSEjnEH5zrJ0e7THG3oHfd6y9N
QOqN45rII6bnzNYZ0dlg+wyEX/oGbqm3P4zcdU4+qbGdY7EQqKZQDoKXjRp/Ov7/
V6mOV9QdKBfmWvgqoKzdQSe0wi0BUFKmrHAGzsuWGHD56wBm3kM7nME4P3ZbkTez
3JHEGK20v6ZDHEizoWuVDXqiB4dNzvX34OBRQi3juENtP7S9l6kGcxrro0NOcEV7
UzNWUY1QkRASU6v+QegoPqI8mMPVHEmOAUfSc/Xv3XZ1QBHe44JWp8h5SRA0Q/xv
iXfY4VOC/zOyFgrEkNG7QbZDt9tUtpLjAj6fnD4z2P47jztLYdRnYsMXRSNN0PPV
xLd0WoTJ1sT4HJby3bkFScNzd8Y81APnYkYQqYLgd2QMGRdKI9Q24nw6r60/IbJ+
f0LqVCsKwr5FrFar/cEgeNnjSdJaZjpdXzPReF6BdItDBbAoBCR9awnGmUCenwYy
BTuQrd2FlBWx50lwvuMBeXkv1pirxsg35k0D95zAUvXDsmNjNpWp/CAoBkhG6N4b
iJvlqVwX0+Fk0uUtFH09RVZ8EvbUVWE2WBXa80VsaVRt3OvOSd3hbBch/3qX0w8Y
cnTNh24BDlJbZBhd3B//TS5DKQE3AOFGrNeulicSpcBbYDW5rwdXyr9oveuLAVUl
J1fr7ECMuq5iGZxYcUwZPIa1T1CkLj6z8fc5MneQTy7QG+pktRy4Yw5TVaAnjaLw
fl04Jx7ofN9BNWg5hFbcLcITWEUpDoHe0nC7QDfV8RX+oqyUPn2Lb8NSWmc1JhMr
NFQ1vjs3NeifFrgw70MWwM0dmqqYHv41IetSBcUdycZvOwP2jqMheZxzAwu4UlPT
YahrWZl5bLgs82YlRmddwbJ7sM1AhGJ3BDBW9tdVuJLy506bdNsBCV3N8/9efaFN
xgztNStKYQcP2uvmInpaKq7DfdgVZAAwlE6kzXVYcALuneslcQjFcHfPDezGF17e
rfXYgyHHcuc/Td3a46c772dw0dyWdR5/OKcHOtNCXlhV36wbTaSxj4TpoeSslvLb
hOXrF/MssX47nFktgywQVP6Eiif7PluuuI0O+5fgS4NLuysCBwd2HBXVeueJ4XoC
GwxBSC9dITOieCJsVkRT8YXpa7RNuOoc/WVHyJuYlvxOSbT/pWY4Pf3Vis5HBqN6
VPat0T9rMfVL2hehDw13gB47S/k3r2nUq2uLz/R8DTu+iINDqbBocFmDg0AlKnSX
Dd9XGddKRiV8cF3mPrC3QDhJdL0tscZoLx6K+xK/wW1Jva7oufL3qo3s1J29yFsV
pqazkBGyXlhFXE5NBr/ayi72FZBrliIIHASGBUEUkZS/eRYzsA5IfYITszWvwUQB
bzTYAFWApYXc+xZysNJ60w08MQy2UF2RAORGTqhUtLhD1/kFPyfDodNp9drCbIcW
6goeyC7ZahaZ86UJn08crwlArt2puX2WrJeWI9pGzjK3M/cs6cgi4loAwkQSxzIX
`protect END_PROTECTED
