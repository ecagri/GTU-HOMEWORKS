`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MMxNJSX3WP+01A52qCuYO2WtjKK28Ojxue8WMQabNI7+FUVKH76eFD9bXmMQ4sQV
VHrSELxvxzawGPZFo0Jt0b8bsy9rHAyRlsViFnaVie/KKkj4wyHtb34ZWtd0tCp4
yjlM7xbcJghjS9VpNpPe4dcQUcxUkzr+4oXr7u4jyFbtOQMIvGsTnSvJrvx5KBGq
OyB3ufFPa+iD+qcOHOojeplDhOebeHINFcr4+HgJor6eHXiG6v/2L9AMmDzyAMY7
EH+/Jl2lSnHP2H8MjW/2J5kzlmUB/tC7O7E4iVSUj5f2zZOV800fyxF05vXOsydl
SZqUWDNyEwyXvcmIDFM2puLMhQyFXLdhBCuDntSe5J+IuwFXS5f1CRxLApX4OaRz
wa7EKe2lhK0QTHOHlwFzYz0uaxZlpQMJxiiAKE5t6wVEZLYBAFPcDTnE69TB5Bw3
CvPbtin48MV3DLTWqt7i1dKsZf60Wh3AJIjnEVrwiZc1fbToHxFyb+Ynhti8cBVB
1eO3+vByjP8V+tX2R07XUT3F9bpDnhjDAoOf80DiQ1/9L6VcQ7zYpmzzGptiHIbj
xHiozdGmNFReryCh1Zej2CblGGGKRSa/oSd+7uNomBk6NTQNGmtdZnzM1rx8Ers/
bdtkHGnIRpbT7+1ZkDnrOhOtJ+cD/wG3leQi9341q+bpPxPglKwDeLprFzu2zRl0
YObY5msH5smslv2PUPDRW16MSEI8DY3TwopYK9BCOJynJEwyEiqcss7A5HJsS0jk
MyE9qPcnENE7RPHdIiQ2lSh2IEh3vK90HLpXe41w0E0Lt3O8uTzR8Urf7JWrQKTh
hSZBd2Ht9WfdVd3x9FuJJ5eWNsfZHTHlr/ZuYIOAoJ9h/JQwwKNixeRiTN0QgqXk
esc5D9Vm0xnuBZIG0s0QZRvjhqBsQ/C7igDupYI3drnJYIs6kJusbE/pKMLdtjVQ
Hvd/wJkrt99NmsxnDg2Ep+NtKmHsYrz8eJd94kv4GMF/DqFXKiCHD88kJOIOVk+I
BJQRAsY6LkEVWQulaNIIz0jKcbcESw815XCrmB8SEhR6ymkyQ5EBf6gr/OUz+Kvf
VgQ+ud2/A8Q/9JLNH87lVqU+966tqPbpn09D31pfOWHVHS+b84C0lURYWRpNWXkM
++zRcqDoTVwI6anoO7u6txRxSUTibpweYG/0J57rj7EoLMXLKUtKg7V9HUS4YJ+i
il1YfvnXgfvZVszudPAPzL/YsVYcy9m0AYwrn1oSV+KW/wdxvuQqSg9wM5nO+1YC
nBPYg7pGPgNTeJV6h4Foq+4w9McA9y0And+QnXItnhHhdW6yvPbVSPNaMRtHO76P
cRrLHjR1wE8M+bvX8BZQOYsueSLYSNaxV4yLwqrb2V7uEXyeH6ed4i6T7+szGbpe
XQkizTPCnF08QAGDWzUZkGAFpVGhidR8nhnauvfEzKsMK8MoSAzTD1r/A4fuASaP
B055cVWOyN5ZyCFnxKK5Djr0nopv5SltAvDhKQQXK296xVVMx6BczMQNxzO6zrhk
H/vX5s1g+tQdmqPRsq29gxXaEtIPjcAmLqChW02bGiZxwhT6QYnrjI9bzrDJ56RV
jTprtk4hQMoIwe7aMf8Q0QDg3hoQg/28giGEmmIxPJ9z4sVrl6mXQssJdXxcu8u3
edSO6uGvBcSzRCR9Fx/LHkab+ZAm0JYvMTYCwuzrbj5SntYYip1JfjLVymmuuVnS
mb4Oq4H7IMX2wJRJ7YCtiJuQgICN0falykAF2+4wyTMSgIqCcMHIYcG+SRB6L1CP
5351OU3EyKF0z+aYV574xj1nbnipeZ+kl2bcSJvfM0fKfcCUe9nGOW83JTDKrXVc
/ukdwL+O95mXCH+ii+61Emi6lTG+ZzW+Az66+15XcBKMNtErsT6mycjnNS2qwgyl
Ahx/c9u6cFUoyKYwTKUYlJ935TTDWUx9lJZtvTP8i0I4WLwuJiwzR4jH6QZKvs/Q
UnxnlMkgv9+oCuEWTT53vsdMzPWrkd7mLQnCgzVQmm6FrxNpvE1aCI6XIdHnQmRe
tWq2v8xTjw4s1ZbqYvQZ1PErX3x4JF60EuFBsApcAIG2Hz7eTacDCMCKBdTp1Nm0
AV8LnfLZHihlKwknyb20ObKEimzWrcjAt5t/eDUI1OLts6cpcUDOKOHhUlDeMUWm
zogMS3oaeTZ2kSz5Wx+uSGheGRbv55f8CuIRDOtg8IMH+cUfNSPBhZEPhPzF4hN8
WLYCRaRe9ATWo4kw0dWGWoG2r3LRnmej5NtiOw/XOnFRIDzXc1R1BPBe0HhueoEd
F/7gVAweIy2Z13pxXmXgWA==
`protect END_PROTECTED
