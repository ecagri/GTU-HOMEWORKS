`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ItC8mOi8wQLdXyDTa8JFiWmMqcaRgp62TFoqTXxFH/4L7GkUftP/BwYqEi6++6HL
KNCJfuuPMQhgWF66Fo/rcfnvVoQV4ueLBjLp2uqfCYsbrhrpV++n9LmvRJ04G5cH
/cWKgQOCT+BWfHge0pgV3JtOI0BSLfblUQX0+5iBXrkg8U6h/zE2jKg+yCp0/c++
E/oV7RstMLiEASfsh5kl04rKLywyQwIzGo/CUTiIDbUAFQkgs5nz5JveS/oTntt/
Np80bgvWwrYspQURlsopP+CZQ7DPwwvl5Dvc9GJ3z8VTnm0oj4K6wtw8N21f6a4U
gXv0Jl5HgtgToh75bqxr5KDJBkUhWVz8jPNGM8RJ39apyLZcvOdCXapKKywa4s/B
PR4kmzhAFm5ekpoKuuIUAz9eS0T3drZ+MVJVvTaaLN7nho++hCvUpx2eiaPsYaT1
eQzL7b8nIPfLyhIC7twvrDS7r7pSQiKtC5n3Zrl8KAdJNLj5Hp6ZJAcJ9yNsa9yG
e0X5QZzC2sVduoEJSI6gLr/wsSRaYuEbfVM0XVAEri1pROD5LnastcCiY1y6vyLX
5Dw8HvKmFU1N+XzD5fDcmaaymBFKtdX/u2sMNiFlvsSoUclI6oZRmDiI9YjtkBp7
k1o3TNPQBKPETTt9b9VtWSUXjGgNH+yx6byrx84PYbpOuJJ0xuVVm8Q6C63fMtXB
CMNiBaYlMha2YatpWuyuZs8veDg2s2h8Q86FqK/Jv71Q+0pcZDs2zBYOt+/0i0eh
PlhopthSwp6woyLdjS9MoIDhMPCiHCUDAC/jSVRfPCKaX9G2bHb1uJwcSr4vPpYr
8XReEA2WtE7wxlf9ddA8P81GuZuwAVZ2Y7PB+GkQZajGl4MMRQ3eLUOX7Lh0rhlt
6tFm1vTySke2NXL5gn1vwNhNFYO/edhjyaYJOK52Vn2PgS18ji0czwzf+1NwVx2W
ivC90AMRZGsAKkxKmdLCAeYA9DVaCxqgBSLEq3eLGkvkgaMqNTwXpdCy3qWcdRyM
7INgPsLtXK6WQOY5q1sbHbtL06qLFb/ahYmill47DszPe1nEVkERELRt0en9c5dl
OIet/AdARo1DIPyMGkCID375rX1yEFX0Jgoic+AhlWmtt9DnoNUpFaVid9Lo7tKF
TtoLQ5fsfUePXCxGrHTABIKOJPW6HqCSR7k60TQ9iO8ZAm/ti+LwhuJPHvYGu2L6
AeiF0Eq6Vqld0qY05wV72Lr/PdlQk55L/Hop3H9+kkvM2BJXE1HyZUrskgjP/fzQ
/W2CiC8eE9X9cxKI5MveUAl+FrL07eaLXJmAYAVU9054CHcAvKJo6nyCWbr+1It4
21/7UQADYFoo0RgA8YMn6Fj+ds4WGc3LXWrgYkc8waw5ty78wjjt2he+jaKFF8LE
Dh7KXVWzUeVf2VqdywvVt28IOZ+H8TF5bSdBmkhfXqg2KGuGoWoJ7Hbe7+zCMHOy
+D+de0t9s1NPPFjbdvHEVbejy+kguJjomcgMqPnc4Qxk5ye3NmTkdRoHJlMUZzdv
RsTmOs5aGfsq26O5+KjR4B6elZCY6j5t0N6lZiJ0vEszTOcYBEI6MeiLnbs+2Z9A
1eKJhRECJnqbxR7ebI3+20w3Br23k8ZDMaw1p8kgaX0g8GE4aTWThLQkHqbI2fqx
gHMBA9X/nRjYCwqXI7S/xX3vQhrb/KSKPQaD7jXLEPW9EPeabRTIsZJW8MQnJAHS
uQfmCQ8Wp/bCzPu0TVm0p14r0TxuTidjOezAxtAtlDaJjr/sxCrbcSC15rGvao9X
QvD7WgPEaQzSB3u+Eg44Erc5uqlWjko5C6hVeNbrH6pJ0iyrbD+f6ytNOdSdQa40
hDIcTkyGG0BtCQDwts1CYAJfMCpQ4bDsK/s5rl8MadJryTu4cGwqNgH/0nL/YtDR
7Dv1JD9D9epbKJ6PbzxpWpefL0l5m7BvKQJ/G2lRCirGN0Kc+o+od1bRudaoG471
+Jy2fYV9yMfAv3zzQxMtsEU0Z9npDqLa56qiJ32no0zWo/owr4w9e+8ukxqT8Dvf
aQnaWE3GpG0noBhwLQWoBcF2A/NCSunfOxpWkTV6AV7KHU+zaOKsr7Quql/KSa8p
DhAyw/DK8SdWyH/B4MDF4LOEUr0lU4P7yZhVXLWBRFIDpJGVnGgf5QG9zCPYrX6K
tEcllb5OrduMOkE4DzhY/8nboQauwM12qDUyMpHXclZbO+4wY/AAgfsiDezK2/H8
N8sblxdymezUky1dD6p1OxVKpmxC7GsjnPHNefoHk0t508BTUUXR+J2Tyhy5yn0J
RCqze6JCsXDmPf8bUp1FzaTJ2YklZjk8RvYLLixEWwOFPk3Ln2Sd3Y/7aA3PoxPT
HCDRv9Z02bb/zOyG9XGCXaOV2sVg4JL/O8UW9Qho2mWIqNGdtp737mOaa1yrfnzS
qROSbjbX5VaiDhUzbGuHt8R3ooEDxzsUvnKsfQaA2WmfhbTKqaMRaWqw//2fC869
XqpTa6ui2kIdTUL5UCsDjnPKXAqnF0CSB5OGXjVlMsWsUE010seSbVnOj+pu7o3v
ObNMCYS28XznLeaM9MCvHF7XRrnjHBs3GgqsA0hNnvGSdbBlwbgUH/bSaMTfk1J2
CPIvU+eg1cBzRrrLH8rxaQ00TT2LeUIApIVxCneBN9ENdgXjUMxGw/iIw+0/mPiN
T6AH5QPHrRZJRsDSVeymNB1kD/qYgAWuX0YUWO7Ck66YF2UxKSf1UcV2fal/iueJ
rxCqk8VzxK7FGX/qaAxTv8xP55i0OcPjIGTbFyFmCCPbzmjg+FZrQkEua0TFB0yz
hiql08qoM+YT769OcktRcNX3EL3zWkrfvhfb0SvYKMmm74Sw9v9uOgHatTm9TwCH
Q++beHekgH9FHOkrYJOSOlU7QcuRTBE7i0+d/2/rnCE4ndnI6vt370sZ40oiQk6m
U7HuErN9tFkpX8deJPP3MgmjalqZLuTfByWMP3OnrtQ2GQ2CnEBlKUQTzwicjOyD
PnvFlmLJXOQvW3iuCnsAsRQ6Jyb9c6HecXzdoNc2ZwH2HwKoIMZMl/rA7VzA1V1k
MZtY73MbyTz45aFGF9UXemljgu/B54qhlU0HXuM9xTQGNiBidq1MEhDJfgkWJ28H
PWw/LtQJn9ueBF2LthlIuFyU4jmZUT/rB058opU6MN5sqY7PkeADS3s3WdbrYEXz
AMeYValmZfOFwIjcu949lIbF1URm9yy1MsNLTd6+EZuu+YHfqzPeo+qZxftZYJUR
8tgXaLXeBPDdBtED2Pn7x7RBCQ/MFeC9a8g7m2nKOhqcEQICbOvj3Ja4TgT5+k8O
65PHh1g6q0x+Hbr5nt3Opc+a0VU2xA+JuyIezSHhrpK6yPD3QcP6tEAFYKl7qFdB
YjqyaPkqLiIgKNmpNJMeeoLy7UIOP8el+TwqCNWwjQGLuZLPfF1xL+ntWhN3QpNr
GBcENd3QvlXDlejL/xeJ/kt9ZAgsRozHrfLcgBge93Ke/42sYqjZR2gFKUW9Wwxb
/C8TQTsGyIh8/Cp4vjYWI5Xqq3u2T5xvkss9p6zQ+UBuUs5Wa3iareKZPcZ5PtDT
XJm8m7MwAWUSUFjbJvGLEJszFsGZUXRVLxbkxYNBnGdVgm+qreCr4ZzFHC6W1hPp
iqnvu59uryCtqnpRh1AMZUzsHaV7zwE3TlFENqMg/KuHIT5Xtd0DY6lM3ngqUH1r
GglHM8beSqQQdRLWViShMiXdhcqKH2kN9Ews7RGZ3n4LSeS23Famiuu/OHM17Qsq
z9DaS92E8h9Ual84X+C0GnbnFT+UFp57XyTXi+/xWNFq6aoZHzSgpFxxOHZVxWh/
npUW4h+mQcIFTXxTkj8Oyio6Sw6c8ILBhcJ961wW1UzmeE5ivhxmJkKAvQ+Bo6UB
kknq/oa0u6hYfBaodYVk03ltuv+5gJkm0GKXJxFmdFIyT0YKcIgtlrb0z+ghriEr
2wovV56BVlC5NXccCpPKEMl/BTsywSrEs7s/mo/o7v3/MFirTtr/koneDIRB/DNn
CPtiiZnFZWJTxrTOAghv6z61TY8EThbbq96cy752oSRz6cLJtOg4llwVx7naGo4k
vqEvsqPorybjfVnxg85RPACTH5dQ6ZhmO1X0T2G7rc1c6pomA8tXb2htZ79xL/lQ
/dAEBq9NsZIXh2DRa5fMQymLgRF2xfCYc/1AarE18/+pit3zvTYUyyXUlBbhy8tR
k/YYnFd81g0lLYdg0JYT84AmuLO2A5Wj0fkEHFpc2JpqAhSaKRnx2kjAcD9reSnD
1Rnc9XJrURynQyOOywzVMfhNORGy8fr13w79P88nVd/gbvivCiw8b++P8aaznsPp
ZvNB/PTXt3zZX7B/XGyrmsJlrS1ZLxBHEdMiXqO81frRA0sNQyDnP478zOr+My0x
izOzBbSPdDgKdVp1sXBqjitsHsEaf2sbcV1vymVbsyp+y9WNhSv83IkdDb5fcA6U
hdJGjNFFF0G5IaM19aEggUm8KQ3J+tbgjDchSjMnxe/TjUapjLl5WDuMBS3Bd7IR
G0FEc84qCH6ILMOr98x9T+1j1INcD+rYW562ZRW0xyVBIQN47HIc5CjUGoCoBmnY
y/uvMcAlCbWodNbcHmDdlydW8p8q4oSFRZ1PzrBVye8uqeH882IoXqJV3r9k+Dv8
mQrfJ9nYQ1xZiIpDU/NrUpgGJmdD+4uWyL+6jZjrKIS3ucReC5ZZF4LRqBZj13A7
2++0TiY1lHS4sIItvA+0eUeQ6r2FoJihEVqcZx8zYBPYmuaZnHQPwtHH4f48lq6U
tsP7ZtnBKeFbRaKJi0Tgmhd60TcKvZw3tRJ+gf6uxq2j+sjoPjtWFy147Mlqvjzc
dJIRXH0cCUdRG2EMoAA0s63pV0CEZx4fTZhAkMBSsQ/Lx3l96QAPPavZZpoIAQpc
m034iGypOr8qTdNJ8YRJAJUdGJtyMUD+6NIIcdX0/cPLDq8N/zhrSwHflKFj+Hpw
0OncoOt0wq3u6cuOJ5Z1PmirkpI5dfxMRvWCs8c4Ynch5G96ikRER6puN1T+rewi
zl1+mGW3ylfShxgIkUEehFhm1cHYYDlfttmgd5UdVVigtJTZkiwgaxkmh3XxABEr
rwSFXMXEEiMgPAQjyHjy0ErwacGGxx+/Xwy89a1xpR79MPHJ8cRziGDHA5xDXFzD
xk3tMkt7vtZvy6NTABrcslVEKyLoGZKyR0eY78Fsh9OK7dPYb51BGHtRumWk4htN
C+/mWB0Q/+aBnz6PaADrhXDEDgzmoYUfetCUCcelxTEevMP3BQf9TKba+V9Kt8BE
LmBkUuemfH7aGJbq1YEXkJfhEcMXg6bGXEoAN5M4EZYpIjkFapZLr0Ml6V5OL4Zl
RMZsnVipyuSdBavE6WTfXOQHGgAC3DhePlUwDPmvqhLVHXKWl6H6aR7+h8R6LZb2
xkKNFoj2f4gFcTmLeRMgWvf4jyAPX+Z+y6TigPlmFBUv5rXhpjamg7WIIDBLZzhk
XDOPMcpzc7jxudhhl5A/FuRzIJqyKo7XqO4OLnf8rrDHSNzIbUuRimeYr+MWqDSl
c1XKLU8CpvsZWiKx6rXVWvVOZs+V+UJ2a4yNZgkjSvEdui5b8wtLWkHXNbTB4C8T
vd3epkg9kxBTuvdB3HymkGOwsOWLPoWzXuR2UqSPhCwbtw/tJEaovOblCQD7Lh8L
Dn2+O9LpNm3vqFKA+pCiJXqPEP90wAVDYIsCYhYkQ34Wliam7oNh2b/HrzHT0Tzf
RpwpCVyBjXVw8J++ZXDz8CYC/fF/Rk8PZa0Ra2OQAM3q0jW/gSavvKGC77Wgxco2
UaBsawDDf2UVLx32Np2JkcFHzzlJiJPRf/3micUMsYVbRPhHlpPIGCC70hbu+3CW
8xroeOWbhPxPucvStkU3+yAQvmU/ZbT1POOAdFfNuC+IZmexSRwwMPRIrq4WE0VA
By/ijXNef/PrF0VdAjCtI1Ufro2rvsGwR+Vgg4UNBnkd2QgYa3tQVbYtqSgik2ZA
va8NLMMYN5jUYq2prPF6nQ7t12WtVR+4rPxLKp3UD65dM7rXxVAOBaXMRYRkezGj
3hznPibwlvhqM5GG4jNXguGpWDQFjtrqJmjknWV53IDeiARLnMo8KhyhULtAYqgX
YACT0YJgzHxJt7Rf7VuTKfpkYm6GkmMC7uQ6c4oJG/DJzHyXExfZjoDJfxlbWLc1
saRXpTKrxyZrmEmR4Qg+Vd8v6Mk5znVi7ggT0/wZq/wr2d6HVhIug8Z4Wu6W1XX9
MV31Hxa6yC3wi/+S833fjPR/2F/awHr6mFJ6F34eFkVpS+yF+Ye4ftVd6DQBqlL2
lKGT264Y6tt1hoisUzH43LnvSXQWWGzbEHV/alKHiOp8AoiAUSepjqrtWOU/qxqw
sGogLqwjM3UIy8z5YuV3D9cVsqFLCXNaNlnIPF7QWwDSSKfDtzsmq8YP5v9Kti6k
8hJl8qzwMopGHvw1YzQbQo5qd5aT+A+xx6wx4haEXIz6o6qApfLtbW6gUPNJ9S/1
x0LN8y/LNAwxNckpBOC/mbGikAcKOfs6hMG2hBxo6rxymZKu/y65hkETK0TvXEcl
XBDUrh7sVU+IA8A6+IuVMGGna7kSKdQGBItUCK4amRjShhix5gkfY8xlNwCZl6QS
150bcPHXVfx64lJzodXqwG/hT9ohBY8C/o63ueciyb/nT6VCQjVhAEgiDOySNkbf
77o3oLRy9vURuxSdgTr4pnAb0EQpDavKL5YFm2X8PDORs/ShSWiMyG0vJunP99b+
ZzlxGTJT7ryqZfTjORbvYzyA9AMrKqZUvkmy1aT6uMu34dSBGxtvCD91PaSIT091
gf7Q0B33uzaB1RaWmQPE1gUZAg4It9bw1Qh6wjecmDuQOeV8j3pZsN654e4qopXR
aXjnEqGPc0f7gcJ7zhIUK05jig+4ScXhKdl6yIBdP1af+vsjM9kdUUAXOL3RtJfJ
/zVG5bFc3arOhgh35q9c74VR3puB1DnBe/2BGRAQBlbOLQfS5IlhwO+JgvlcAbgq
6oGz/KJFe1SeWAJRuM+hbdr7/pLfl3TDiBczeNTS6mLtzA2AZq71hWJq2KO22bFO
C2mZ9A6JbDKSQKijlayFbO7bdNTw10t+W3uz76/8h/XrLiPBnLWc7kx1Kn0HVClc
I2tBEEVTskmZ247P5mhl3uwm67Cg8MpixTshEgi/bH3qbhKhv1xqubG2sV6uZaeY
6mjw1mlw/WbL8JljfzJ3/3+Et6H1t4Sih3lgDtGVAa+p6gkAzDQblLF8De8pH4xK
JOz80AHB9d4VCSQf0YKhsdBIYdEhCSlXTPh/LbwIFBfgInEQN1wwdHzsjP9MT9H6
gBIR7VWiniRrbSD9C1jcm6IlPmpwZMh2QdsRA+B17ZyM0fL98ON0PVA1j8+KzYIW
88xDI7YylrOqC8d5dZQmsAPm0S8XWN/1s6IbsHjn/qoOOP2mPtlb427DDO4scKNd
DEOVS8vvLtZLQGAbZyY2waOo7lpyv7X2f42uH3Fan+KExSpmeu4m89CCjPjpvgsK
ul7Cpp/bQpc6DV4zOHehu4gH6xyRA+lJ4mevGTEEdyN1hxjLGpNNhRS38GlrVtA6
p/HMok/xroyG9Kg2b5su7Kb5Xhs6ex1eHJu+lawOvLHi4dGNAy5rounsIEJrv6Yb
vpnJGV4CxPpb0Fx0PMNbbGfboUPfjj0q80iC/dg0FUC/H++XfWEd+D42Z1MK1G8T
gnFzQtb44eT9ZmUdly2jvzzxlIPa8/m8hL2zEOMnszA37MN/yMJAzYksLjcJhXrJ
sLqxjuPhXBXp2EGcEGV6MuUR096zJcnGREXxBIwy3pBy4i7EKTda0QLIRlM8YM3P
5ok35I/Z+efauQfra5ortlxpkmYdQuSfh6D8bEr2IrI72VEVrPo/b1D+396NMFeY
jgrDvDe1mlv+HPrZiQiAoWyeothUU69Ffrew84A22QuxV4llnkRCEbrQMs+xJQbd
dyIx7R+ccbzCJ23rnUrbYlHHzmFcjtUqyJYbudJSTCwTmnWlKvEkX0MhqMGxTTgn
ot9yGhXvTqQfjmzR2a/qKITni5/k5zo/+Z/0SETjLFou4iQQXV0iC3U9c96XgT6u
`protect END_PROTECTED
