`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/ErzbgnGdbNWHzxroRS3yC368qbSmah4nUs679R33fCBaPGLUbeo0/AZGiS++WuL
lov1wKUn4k8BwmCaORh5FVYDDPc/jpkfNfH/TFnpGLwA1mGm2UR337FfWQtQMoSQ
5qvor2sweG1vsYXLsBMLZ4TvZEYj3PQf57Lm3nDFy4rys8DmTM9jlnxwvwTU+xFr
x535k1ZbYLAdo4vgARGJngA8klaFIV5BYNHUP3ALAmRiw+5m3nti88SCmH5wGo6P
JXlRWrF76Me5uGbOGv+WZCxQZPYoBb26TaihqKnu5oZlw9G5Zz9gUeZWRmY5xAlG
G5JewmrJPdAR7jaJxViuOxfSRuaQej2JBIHagHyS/gkDxLpIFIEo/6oWjfJCPLFR
rGHRVqBtfPqScpHriK+Xp95/w27A5LS1EZ4JgkRI33wpM7Ej+Z8h34PLhBTWOW6O
rLIflqaL9m2oFL54HDqS0rCkWBAN+T429kHTankKPdqiCRAi+lkEykQ0OKs6y+sq
cAGQicKdwxYgaKEqP2YKrNHaulXE6g7q+TgRB0Oi/Oi0BvIBLpGHFv2lXNXbppNZ
ZxZ8r0s+SnJOhYn8Snhi+Ceeg6hNPu6nYk+IVE4sGQ30DSUagPzfV0SAZMNWUbJ/
XyUxEftv3XVHzHHXbNrnPFs6YvC9ULNztJFif7rmCT7f6MYR94F7P4b5/NcGZ0hb
Y+mfGzgH93DhVzdPCKsjmk6pDdDNAUubQU8daxediQMz3s5ohBbzlb3aSUGuS/lJ
8moFvu9iJKHlBiHD40VZmJ6RQ9U4Y0wQ116fIFXLX851Zy+sFZIGrs7FVo8fL5TF
snVq3p6ft7qWcbyd0JU8qYnV02IKw8LFf4kRvMLIV7UlpWXSAyZ9y0pORw3HUF/y
CewEBoAXtfVP00anYxZ0W1ZpVw6ZG49qfeLSphQ7mE5xSSPJ9NzOTxhfxsZEvtFq
DLCdrkLjB8mUy8Dox63PNSge64k9qb6OEgADU1L2fR53gvG/WjD19GtN0UtxyzbD
O++spN+JE89O1pE89SUgmuWc0rhqF/Klj7oXRWoITaMqudTI/qFA34r4lR4l6A6S
PvLNtnZkTbee6LivGa8UuL99Koa0MGqIRvedUFM3VUlMLEPTK/4Dh1UJqfhWXmKD
SNpDgsMZ+klC8VgW5022irzLrF5oyTdSFzxwO8glC8X4UQvOrq8YlkMm2zy+UFLQ
Y2cEg6izPnmdqfmMn/lZeebq8ae591VnlEsUBnMMFazhGOFOFg5eMrWrmBKiLnxi
oz0PlbTAowPttTEw2eGVWVqvZenquxYic1BfUCRyoTjhLT2MVIo7aqXFI7RTdwRs
A+fZ/ak0RLOhSrdutv6cEm5RF7TZAQx8+zBQ0CucKkHbJiVCap0N/IGymMEig847
IkcxNm+V8bgTgJ07hz2MPtIF/tb9qWTuCRYrMLLTCMxh6z77K/it/4RwyYJcymv5
d78CGYHh/PY36K3QtOgAQNS8hEUHy4HCziBzODSUtNuRfBHvDzb51tU1sNpRQ5HP
kjOjXPrLfpyQwUpfn5/Msv1Ubg84dlTd8pGq3ygMO3LXf4HjYZCwqcV/fxeASK3k
v+Ky9S8N170vB/XubIjT+MP3sz0GT1i6VmYYiigkS7C126gvoyOFYSTMONzRGd8S
bYUqTNgVFJhv31JEZzu9la2ln5UyPiM3jzA6WbojYZKH9T+tGT1mu+MQzyljzrLg
FaQKpASyMb086lpBGe0uCa2jSQiPJ8QskTmGGDqQIGHJsMYuP1p2LGPBiKCYEU2q
iep+KDNr6AMDZP9hVWhnZcrxuByJ72t9WRUSvrY3AFblSM7nROR9rObxv1lfCaPZ
P+t0ma2h6LsvZLdAgx84Uex/s4OZn1pP+7TjVGUI2OzLvuAKa5WxqslGLr10xM3h
BDv6sqrR7aSS/h7lJ/RvFNQ+2LbBCz1o41ANSd5pSTz/CAmlP7EfjfIVtbM13/sk
yKPEVRY1jSTKV4ZdAnKQSMERafTXpkXofWmah+9M+FNhw+F0E+WrsyHxbeHipepz
HaTLmumgLJBwJPbCs1a8G6udS1QVWlfNTqy2k9OFXkiq7HD3tH9rWwIn3oJkpC0E
Irpr0ws96oG79zvXEmqGSEA5z9tU3//68Kmcrn5YnWE88oBaV4iSy1a1PRE9QReT
rbPMpkvP2DSnCA/OcjusyBeCWUUrMNCizeuBUaxLNiZNWf36SJemNvtJR3NZCe5p
tphpfsOAX1fEDtYtn6JRW6nSLHS0JywWPF9xkfoCoH1nqHd8HrcwEFg63EDEMdfI
hPBdjLhnxjG7s2aXe7d3UfnImpzW/czf4Z80VEo/Vmmt1rpvVmYDKrqZuBVSqN0k
MUUPIa5dl/cSO2gH6h9yFQnHTM5ydb0EVCdBcpftGs3cSjEOpYeMcH60bo3J8XBM
r47PV8pskzwqILj489eWKGiysnUoHjJDFeRAoDMBmFXJHYg2LE1qL4jt5tJ8hxZb
y+ydU8CJbfvNEGWdUGsdcrUAp63ko9RqL5md5qMVIrDhVExDPGE+7nR7fAwcNfU3
LgUTxE0LVU1razIodWjBjMPe2yfayD99bTFoE+vGMNSBiYwfs5MI2FYDJ4Bn10xC
q4mvwbUkdU0ILn8S5KrcsGg1Tohi8CIYj9ZKlPR4uDMfpVxxHp7h1NfD+9/JjesJ
`protect END_PROTECTED
