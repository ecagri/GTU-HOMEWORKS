`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
degBmBTzmu0gq3CaRu4nNY7ImIn3FMTzZqA3SxQoAG/a9WXCAV88/9DtzX86QRz1
OIN+vxzBLlmIm4c4PAadAxSJd4WjNeeN0UBur78q6ijo0hvdjpxvfcsfq7tSG+6p
2uvCpsMsW4hrNbYM6Y3YeuoPYXwfMl1yk8KGvh2tL3UCOKpsa+JKetCWw5s4yZov
w0Weow9Mppr4j7u5ANjHX/WC22xshuk3xRmotHuTPjopwrElzvUP1vmQKBXTkGWN
ouRXPK7ziLl4uToxY8v7yGVqnokhw2g6+IL3CxgNO0tptgS3xRxfMCbI4Qngmu8p
pz/Clg3FI+gFH4Xh9QfRlydM2mbdQIr81JAPVcbQwGExvGglO76AlZ/JYY6mDDSG
2pwrPq4NGik6iBgJ7ebdttdromz7flwMXr5FGLb5IKoLBNTtViqfFBcwi74oUAXZ
qiGEQfAqrYb/5AfqEWQh+XItPrOwUv8gULcb7f3VcmDVK0ciXQKTGhH+FzIcKuuZ
mZOvP5XoC2pNwySOtMDP+2p/OVErTgOyR8PQS9YVcFkXVxUJel8Q195xZClW0v6i
1O1eEWK1LK5/mW4U8AG0jdUjJ205mEvdpMXC81TE84Vx982WImbOzP0p31QryNx2
up/QzHpSCqZl4Qxi82PdgT3CyaAOQy21Y6Y2s/IMhuIGI7S6RvhoENeBdJ4kfAvQ
/jHGX9zoxT7nfuPKiltzlEr9tjnyBMHui+5PMgYbVR2VLd1aZTEUjoj62GonPTcm
0Pm7g1z3DRZwZc/CbdHD+lZkaLAyS9WNU8AkfDzvdV28yci6FXlgCF3bxexVOEP8
chfaHUUPpZme4cEq/wllV5PE3JiNmgCT8C2IYhYUYwX4tb12aUQDFew+wgExR7b8
07znc6bv6tomjfyDGVUEjlQuYYxLqD2ugntNxB/Y1pw=
`protect END_PROTECTED
