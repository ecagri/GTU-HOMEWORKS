`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WyfSFfPKlfigrTk08d+xVSrsLdeIFLWUPCYzPyam4SmxMyWyZgvPdCl5+2lxbDOZ
9SvFFggerjyAlHpQh5tUJ3YsJkmKJ2/RoP4Wm4+U+4QdJ5LDEUYgxqzcerERuQeq
vUKBEHvWShPIEd6xDhtoT/bK1WxjwotuSL1163e01MLZNj4qKRoKJuSIbCWrzB4v
vtp6bkPZw4QizVTF6MGBP6x+dgv9QMLWDnixGWVNvwnX+k+2/8v5gqtlzmIe0I7i
5zXpngdrSIM9rC1nu2pbdpf2Lr7hMEYU9bQvYfL/6y6ew/Y+EEGe2M6T1tcihhfQ
JSFl31qH5xVJyahNb4ClRGpAtfjxcOtZRVJGPrIjnEciMCw5SD4+owxCNXdc36re
lgXX8tUTIsz7wWEskmgzUKLeFlfcpNj+HAO4bbri60qK0Tkz1vBKW/qhUNwltBBw
TuSC72sG7Ibp2KYWteq2s6rHYbW4saukpkxxlfa1euBM3ZsGOxYSVZ7ITTiaco9C
WlwryS15t4sRtwKNwd1+eiZvgWvr1IIuB36cAGFaphkIZd4si5gDkr/q15wuP1kp
lMYkw9rNbI2ZqlfugLjkEI4DbUGkhWoAIurDJN1juiqZC88w6fLu0Daa1C0JcTlP
Xd5At5IkjDx1CuwTJsrb8bXZAcPYNf+3uU3W9VnXEKvOZLPzRaaKzyp0rYtGylJ3
yyg0HUDDsO4oHL91OMc8ypssqJhqmJTf0mCTxd0O+KaeHvSiA1DuLhboZ/d/qSDN
xOCtiAIxxVNH08BPkKTmBNaBljcoXWgAQjzjk0+PsBBmi0mboGrNZX5afxSQf6XE
obcUzFpw70yV3oT+9jsZ2Q==
`protect END_PROTECTED
