`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q4guWZ9FucUjb5/5dytvStErTaosIq/0gxi84Xjh2IETXOTme+A5PAkKiDbwtke6
KQ55zaNkEv7mBqya3/tzKAOEkD26Seqhxy0u9zicvhEGbp818UYH5iBS4ovIlQ/s
xxoYneYM91E1x0KkDJ0caoI7ktmv7Lv26n2kyw8tX3eqHFtDwtYiWvBhvCKTUXcz
SMRdhGZytoLUmaXo8XpjeqrMip4otICtIIRYws0NyEu6Ck4qeWka34w99ooJ7RM3
4gHo8ILR4Z96i1AplCJUd0WV4ddkILBxga2QwisfJTTaa9B8sppTcAw0l/loZ9um
2V/45QZIvMD36oVIt/vSHdTMs85BNr/ZRsFBnB32L0R3mglCrejc6q/m5CYHuFVv
KSNcBiLjCDg09HQN5Gnr2n+3AG2rYre5IctC3PP0DKYP9I9tuQ9toLDje6wcLhBh
OtulnDH5QjqHmnDpi67QWGqKQfjC8meZxqmuxcl73Asi/8QqHaF4qhuG6cszPeEn
W78i4Oi88lNcW/G26gyiby4Rj9x7vHVVxSAzQfGwe+fwXFvzuCJxPnmRU/8C0bM3
Luwzo23ZGD0jT2kYvWfjTFyXMzuDp6PinYKoPG1D3k+urHKn8aoSYQjCeWYCYwjH
2ECNYFQSyvfj+8q3V37AU1/Vtq19jedXkl+FNDn1wsD8YCX0Uq2C6abnbHe+GkKJ
GyFnNHMOAnRlYX4qF9YnKjXhd+kkn27Lo6GwnZDMRYdDXpXgcszygSzTxp8p4DEQ
Si5+TrYwmA/pK7fmxO28IkdyTyyQY7T2Fbb0o+juvKy23hcIpGb1fc2I8x6WlW3c
1ol4Bd3bVdYOd6aqRJCTfOvzNtJ1D4QP/hVjU+Szgu+1H8dTba7f3HwpqrHHwyDO
1uFh7nOQYdVrqWUp+Hll8Sx0xetgYXVO7P2vcFjAwOKSTKP5FgPXn5tBgc/TfAvu
YSdlDS0VLa4VYW9zYYv0Omm6jmpUUXqSQVdLpMP1wo1sBphwfXHCUlcxe1bASiVL
x2u12f9n/2krKtYuYhUeBDt9rCBlWH4Uxie6kAMTPG2rNVX/zHiVCE85aSqe66IG
/wB5OPTBzwuCYS5vAS1hPYf2ijjJ0auUXrynveE8DTRqAtDqJmNbP0AyaP19Zibw
lYlMM4c+dceNZhzQOGTUMIGDDmUM7J86M0b66WVc4CaMAdK4NS/YVxnfvQ+m/LEj
BwrBON75uoXVmLhfeS0oJ4Xz/0qaoS0iRLjqJF7XNrOc0mTazecfmyOJAmx5Kwk8
ipMjiJ/8rJo2e26huRvWaOH8hP0h1Dse3nUpUp9w5Xg64uYfjbK2adA38ofdsvaO
afSCeVdigJC+yFvU2XL0tJSYbJF2VnGSHvXVL1xyXYApoimyM962UuIgLoi+HLtS
YuEaQz06BsyZLDdgGO8oaCx0B3q4GGanaM+Z8RcnKTDSQHybMF77ImEo0Xatyris
G9j1dPjm8JmPsTjzhOoc4WL6aIk3QhkY21Orvs5pyt65zY9gZ8XFBC8uzMeS8Zfg
uhEcJ2FaZuafbf9OHOAU6wQxtGtoHDsKUi+yLEUiZV7c7CuQW2pxxQtDMvl/au19
j0tg1y1V95Ro+Hd7n2a91WaV6Sbr2+Egb+6mZEVBu6464PDeKz6ughXJVax6yMB2
lY+IVA+KlCHjTOe9FVkC8IFTYfwPG6EOKX2wTmxbDQ5jzJppEekZfwE2tEyXKC2b
Ia7rN27IUyMWtO6Jk9QOT83TEmOG6ZyH4Tbbw3TL6gIZtMa9EZDukGb29n1vliiI
ifjswB62NBYg290qJm/w8a8TZRG+c+TGdG5YzmAMofSGZ6gTocSI/dQGz9WPNVSo
tJJ4qLM4LPTQkyWy7ZA4vesASExJkYbueD0rh8bQvCwpukM2WpZjJxVAzkkxXWLY
22n0C9zQBff670ycZXKXYN/C56YrHubU+eBcbJwxA0XdMlRWwV0Ji8TAQ8PRY3kX
z1f1caO/7WntUSPentZ+m2rVYfYAasirR3LX8dwlhY/1BjR2+FPC0W+5Sgchrmso
vDqLIz38nzQ5b0+2/5/+LCaMfudLo0yxXxmviW1S1Z1Prw/1Uutlly/XXn0tN7rv
5UWVo2AQWWZbFjvXs5oVMcoP4CKU+42tRLjdt5lHh2wZ1xsOg1CuYz77tr/K1l4F
LyayOCtwFVTDdTt4Pi55ACsVrYRTtkFaiB8YDKKaVgu7IMi+k/q9k8W5g0SQSSXM
gbWUf5Y9/mUKrqJF1LiLSB2w7G2EGUwWNQZ+pi/pDrhIY6dLRsw4ThEAqPGNEXo0
swBJL4R6vr/vcf70iAypvB0hi3+bsE8GW/gxFJ/iKLLp4mo6O1KW1VFcjTYN9ZDz
QhJL9X3PKSrMDHtQlWfXTsgzNA1NVVKdLfhsEWQEXux0KeG0BNUlopsSrazIs+6e
FNe9cChhY42vIUVtLI8d7Bg7gbhxOGuKFegXzF7TmMY1ZRwuKc9Xs0kN+2WJII5o
r0nqWYyeNY8pKTo5Cv8q5sQCgMcsBknbGRziiw7DUg2tkLV6nGWjYoPn9HM/QCK5
X81b/Yp3ag9aeWqt7R8SfrDNSSiDXmgw+yOOaanqJt7jxMj4z9EXqnIhKcIloKiI
qTNQzEYoVHkqGYfVlTKRyHPnxWTyIe4qeH+I2bn/facYJU+BOnb6jNUMz/nO3gVS
XrTFg1GsIEELB+q7/xfipLR1nF35Bk9J8c1IRGjhaVK18bWvapeERdhWqqU67Heg
pg/ocWKCfHySoqLjv3jeSGss8l0mjH+KuGBJcfsjF6XjdduUvK2HBVSE6tp7ZyoY
nbqpBBk4mAJhkH/IEevsB+oWbRevUSks6rw40UCk9piWZKzcGyq/dWIhNp+z1m7m
9A1L9KzZR+SavQjVSWrrpsyyahRD2u+RjDECfDXPcDOutzNAIPhkDZbKpzl/s185
OgxgNSTVdrky61ij/hwS0YkIgYki04NUrSmqOiVeqvbSCW4xX628ZxmagJ2l0ZSY
Ph3gaQZS5WyN9cTm0t8sGYiIozQACTgrz5P77MHi9jRgG/sPDUBz8zbvC7rIHhgv
YHwZOGzxq5KDy1tt+coQI3zoDD/PHqkEKdwieOkTR4KDCf5jM/nXO14DBFkTeoGL
Y9feyfq1whQnRjxRiElkMJCgggOVtmQdQ8FEI46mDLKwhY1uBlRyVNXyxzeW6CZ+
/pFx6kWHp16OF/UPNWz5s7MeGZdT0Rs/701+Z75GJJNNXR9P00n+ZkZfn1jqpOxl
5s32tpR4PXauKPWkSypcvyDFnQkoe0Xsll3rWhHz1c/LZ2sWlIns7FVSIRfR1VP5
SDVp8AUducxWB7Sjrr8T3HWmDdcXOsIGiVKR+FOBRvwZTpzKMvQYGJTWixUdpwDA
8/cG6X7WH+SxSCy8wPZqEjWZ/WupGD6VlZDJTHXdC/YL47FT+uiR5kMFqq/DKrGh
aAr6YFpw/Uv0NBhsQ8Hqle7OOvFImbApwv5ZRzyX/3IOauLyfJxWsQEcrCqsSheN
ZQIbQq48z45jrsuh4pUWcKD773hcD7JKosaS/VKArSjPbZxP0wLcZMKauoPUcRMX
U5mcuMDoDr03wdMQHaB0lSIXmxCHbEyI4MVsqQETPI1Y1/jFAljhKCboPyso1wH+
ohmcO6vsW9JeTW4fRyxvckbccF4cScw2apPzrPkoC/QtBJZgpzhemS+ib07o2AtL
8XojV1sSFnStmICnPeM4rdY1kP2G/UX3QS2EWeo7CFuDIDO6FRe1I1eWoN8GRrEN
XzxjWgfpOVl5Mi76A8epIy9pSSkaeA1U3ZEG+2knxJKpHhX3CJ0KUn4stZV7T/Bj
eD6EUc4k1ye4z9fQDYTHDFr1OT+XvNBifbILQBX9DXzz7fm/ar6uCQ40Eo+1+jXz
lIiYjzN3BJf+qJcn+llvlGzhi9+jcvl+vO/XKe5QilBztTIjbslqlKw76LRgIg0k
2cY3xmExnXhEoPZ7HkjkJLcLXxsh0bYjYtej7xHxLHcvk3qYQJQ15tkaC11quuWK
fKm79SNbW6mHiPGZ8/+vn2IkJpBXUvNxdl5cCYCxtPzuFnAiNVpAmd5CH18NYI0b
Om0eZKve+PfVvj17JJfpuW2Xqff96YjJ8AY5Ur9iwLIcqOuHbdeNzJaBCTdm4PEP
tpNkx5hiOkfh5vamibdgCASoYu9H8e8Ybf9I0tCL0vAw6sNHjstvePCJehbSiM8r
JSoeEvzDVhPAxovKRM+8EjwadHp8WSCFN0cVbodvQZ039dys/nx30iCPJmYlWgIT
j1LJzgycq3YzdZkjVTPKvO4cDM4MxylVKwE8aQhsXe7A90BOoGN2hMzPlHTn3nfJ
1+5XyMLdLqSA8u6IoOLKteZffb+SheWEjIImTdrL4rIZUyQHTS2lbGobTZbAWuLr
YmvyLyxzJfbQ7aDjfbEfkxce0uoadsMFHoZgxMbwHwphMhodiykb7/6S71quUyg+
Qz/ZtIC9Eq8jZwFx7g05PvFpykMfXz52khlnrB6mrfyI4riXzvDeWvvtGx9JceGy
Rw9gzm2c0ZwtZO+hzWy2ZZ7WxbiOjABGFok4qRcEg8OuyT0JgcmhGpPRxx1GUPIV
BdDgdvVgTp6SY+kGh39vJ1n3RGY1DztBaRGYsXYFSVF1+qmLof+5IHja8sWgxEBe
ZgksSNexvSBdjiHWLqwWbmBp82NRBN5E9iSb27MLZIxTNW6dRZfSEbdBxaZzaxGL
dP8zl9UJUo6fqasc+sIRHbE6SoYdaoBUevzQFQak9v6T6+B4oReNQ21ETJHOCyzZ
xZH5Pqy5vWlXqwkMc6tE3f1aiwUtYekObSnJU2iiFGzgrlq6D5hYLkezQd3s2Akk
zOOStLjhEXsB1I32cVL7Ja5XBKjWjRZ6BVoGH4PNvnvu1bkwzhsRWPm0yPQDIKNK
24PEqmk3ZtLpzK2R9DzD+PyphjnhZM0Kxj8s6bPLJm8InYfaKZQTDTGaK86hId4U
5uu6ia3zHzrkTbxD0jnDqgBYgaDJ8v8sAAnnyjXuYtJNEDlaoObBE0kKqaNSr0yl
H99xXHatPp8o08xQqdWMk1NxJ/SGPaFjfCxN9ruUXQJYQmUWtNtQ8sc0LEsosrpG
KHmZXbGHU3NsNekK2J9vmUvAtTitJAwdIqaSbxBxZF9fiVtxQnlvkyqFVcxi4NL4
bNe/pecNmBM/CSsYqnr2F4vrGl3s4liT0W1iA0cpiUm8IRU2LJlXK2w9d0rDFKNU
2CykFsvcYSKE6AR0C/HZdVpWQClO4b1RTK/jdWYnkwh7EWpJzPxyebuiw4gqVs7F
STSGzGZ45gj62YspbJIMtTddzkiWpyj15mr4+bYOnebOvWWqy8eQ5qo5Gg7+EaMp
qAZqMdDetZCWrzeLqD8KLMmmeWW39n6GjgMa78/OqJGzY/yVJqszlAr2fOzzlCWL
ySh9R+3eBl0UfjrGLpHcvu52Yzk0DHVit4QWHYGDtWkm58QTVWAM7Vl33bwPDOkV
tRtDXtx/5WxjqDHCmQjRgKF73cruabaoNZC9LMG8QrfPHnLVkc3mYMLB2KygWUl3
BW0EM+AQIluB4vck1S9udmSgRXjHrhiqsNTSzJcKtWJUhgv0jZHWA+W1fLvIepPZ
1lippWsBgJLfVY3vfnZUKS18epb3fnA33sipNIaYy5MgcIdDRiyGcRLy3SzA3d4Q
OsnASj1DrMQhlYgeblI9VPxbDjfsamnh2hf1d/7zM6QYaOfuv1YRW3USszuNammb
kxsA2c7N4tQO/gE0Jj72GgVL2iTQeg4o0+LavzClBr0SsG5r1hHVKFROqTbGvxTv
wIH+52ypZcNHBR3eMezC3n2NvP/lWMml7TuS6K5jblKf/HJ6kbV8GtHYibZHBBeu
uLsQxgnbH41VToyYc2qAi35KOE2/HuTaDZ0bga/cWT+CY6uIKVUXgV4b0ZNHscWt
/dmVglFI0o5wcANkj+KgbLHcBX6V+E81JhGXY6CB50CKSuMkCBgZaHo3haL6UFj0
XqVFnc7am0q9RMl4QRqY8j1oq6Jt7bQHf3J3cxEdMm828UCjkKc9KHzl5HQyNZ48
Sr6CS9YofnWB4sh6+8Y+p0iIBiZLNuQxGUp8UOXpu2qBpmjX9+9KsnnaUaq9buzg
9+T/EXyTXW3wgnWbJgDGVjvUQt8fg6+gxjonNKixz62O6Mn9y+2GICJeIwNNuuBa
7eN29wvI5fIBbEM5cofhIz5Jq0k7o8bYeYmhW5t/wucHHgsUkmnKJyVcIHt/L5EK
rmpvoSq3nhhNP2D+AvhS5TPSA3kWF+eA6718onPGwJPVCQc4h/9/l7sNzNHizMWI
WzjXo7EmjBDmeemNf4ymNA5tX5yKr1s2nZATcld/7q+6MCTtuORKBhOKgo5WxlH8
EBYBPF7v0WYtX3Kdwul4YV/9f467M6eVDWE4Mqh3q5edYXkIWhYLXrkWSXQDRtiV
Tps3DvZz4k5nX71nM04tl0bNN7QW520UKcfd4OQR6T0OvdbMN4rVi408gvyt5MzI
ZEHEGk4nA6QpCI5X3I4wVH8Rjdgw2aMKRLnuV7tREcwYjIwQ0WHzN4rRrwS2U3yn
KT+O3FIs4cvbimaQduzp5PgdDFjxCC78eDAQZ28P98cTycX8VSHHvISv1YK3qSx2
uccfcSLLgFwAyXsk4vMMmv/D/ZYzfZQt1acJNW3oj2+VB0XumrvhUhTfxNm8QW3k
QQvzz/VvrS8GUT9xEI7ivitJipHHP9fdNMT/SwfsIvZUCfEFFQbziuFz+DHUBMl5
KgarU4lUzzKMbD6hY3NN4z0//sjJCfnjBKtnFJEpTo61xLKwxH/Osb5z4QUTR82F
2vSKcWuHCfbImOIL6DNBHz0wxQSSS7KcD36/tLgqn9dMYc0Tn4h5cHFV7YcmF9kw
OyUn70pxeb9SalJP8VqwsPATqq1SaS8gR8nzY/e7Itanyayoh0nEhEUn/O8jLd1+
gd0nHXHHj4CY6bipWggawcgis7hTiSnD0w73VQCXlo1W8aOcBp9gr6LM9H6g1+qx
wFpztxjgSAOCaBvQ4FD+JrhgTeTTJ6PGl8WwYI/o3a7C+bF5zAXWvVOw7IDiaSs5
IIjMEdjLayBRcDEz+Ro/rdxwe+uH/DmXa2BxdDAWJpU14+fRnZu3jrsQvgsW6ygI
e2yXBW8ULDVm84VSXJeBDhGd1PD3YxjbpucQJE8DNnKjMHoX69T+rpFvKR80KsYX
PZ0J7ZgyXsog57Dmxp8jDLnCdvJlik1LmUcaZJYfniPuxVpNaZrusz0s5pmgrQO+
QugOaaZOpPKb8sYvwOkgS8pIR9JsjDSdU7QD5LLK4lTzuVqjzcXPMIJL26kkUrBL
SINwqSwfdOduFdIyhxXgaOAQAGTcG5OmvUy4dax7sVauKwYirt7U49OKxZHCdfbM
txlzSKRgc83QqAKfwqwHKoTIuJvBtBcnAqBw/oX3pRIS86XADXb3/bqT2Zk6OH7Q
wFuUpkxtWj5al1euuU8AjGh4fiZEIRbCqP7TYU7L1vAIG7QNcJwmm7CxC4c/lf3K
Xu+yOT67V2OY9aU26P/J8lSnJM/Q+0phcAx1U8HASPu3mqLblzD14XU9YeVCGcqW
M5e+y1/U7FKvAwa2LOFkFS2ZpQwKufRK2YJeZXPa2HqxQIExCAPKpjar/OoWssUQ
BZg36NPf7vvjmm7tV0AE4FIcCfXvTUBIwR2J64gLupthoKUZ9Tw8919C57k8KyuX
Emv/8axf9nD42ghSsTtBc8Gcv/zis3L036gqHWKLaND6z3nVNU9XWS4gHFBV36dv
bagTGIB8SBh8tmgpKnB6eV2OJ8pxHa5ELbld4HjUyM2JaAr94Rn+pHUiV942lcsu
bfM3dP8O5hl8FHUJj79Mf5c8aWhKF7HfUhGOTbAOPBwRREwy4IHHT5H93qmefxpt
4xmYBNsDWuy0OWl+dnBnV+FJfHnz5VUTZX/Q2AYtyCgr27V2PZ4dnQc2RB9Mw+jE
WiwW45cOwCENOVHL5B6Nn2PsHuBARVe2hh2Pu1YwYXW083ox7sZbPKlQUI+NEOQB
IZhfygrLYJY9gW25pkPXcSz5Q1S1XWCPwSDJEp5v8er/1Th6uL/ijKh+j/hWsUcN
7c7aiyLtyRiFUfNp+lpNz7DUlSVUlNdA+6w9Njm7hDAThSLx2scc7259cKzgdOjn
sqhaaQi/tL76Jo0USapgyWa4VnUMN1v/Gf7nstoERrkg9YPpNoUukGQIvKPlgDaw
Y7Q4JIOr81TgEG/9z2E3rPwD+zHbvUdBupZsoxGQUU7QP+3domB0fyBtFtMV7uJY
cy+/lc3wxw3I/dqRRPKdTcd2ZjsgwFNHwzlveeITl2w3KeThbXzYEtbZg+/JtAFS
XQ3nM2qLnXuOl6SLf9qWe8N0iZStqPlI5GymKFaP8vrsezwpvxPRFzKYLapiZyj1
ELY1oeDom7wmC5Ru5aK5S08DaAejLl/NFk+YnmwqPjehfAWd7Uo0ZBcxnGYHrWG/
BjPyOQNEDf4mAQMl1J/1OXjM4EQ8rbP658ivq2XtgXmw0brOxfCi3FTLpDKcfQ0E
ur6A3ZLd3ytq8iwAuE2f1It2IvpKskriofuxXMSwpnSJj3bdLb26wcgc2lmRfFQi
xvq2LZmBfznNMobldiEuMTEjuNWcvjS4KMFHGfItr9k4XNzlWQO+l4VnWXSmB6bh
uKbadj9Emr4tUkuFb6s9wzbdv78tblfv585bhMUzsOoEUeIflVz5qUnnBL9QdKf0
S7BXqH8BkupzXC+XclIoH3PxUXziXG9zO0JHubPFna08qP41fAfcE/wJm7WgdLDK
3QGS+p27i+XXF+gXXT6ADZuBnKVythQKHBr6ggrIVBnhDf1DP/qL3sVuBjAvm7HX
1iPXK+l17t7Ef1RsuWkm3gA3r2I/qeCp9/+PcGryBV6Q6rdWeGv+Qes/nGftF7w1
xHrb2ycoH6TnUzJdbxj0U2JAwnJ3WX6bV8uUv2jyKphfMKV65Az7/r+Av+nQGuYs
l+nd90/EiNPYtDWG3DxDeaBT9pBLsq6X9n21mP3BJrzg3MFSuFyVdUBzD8wIstdD
sVGc1+yz4YJP7QNd4dclP18vpIFvSF6DM1K8AFL15bB35uAiQiaPGs0Q3uoZLoWE
56JPGiNQEKbCM3394kLugY+A15H9AIxsOVILkxMaIlBHNZHgPBH/pZxPWNdPnTni
8KEVU8WRlF1x75812F2ZJ8C3Ff7wJfY7pIv2KVwgHxp/61E1TVEUbZkDCHYYenb2
a3UdG7yllwj2t7y3qvswVzopBAHQGOWIyqAQZDiIwOp3MQCmxdcbmSeyWxrxNHtn
4FX4E/y08XpmB0CvbhSQbkoGK6wC93+bMl3/Ybkf5F1UNPruxhq2yE7EXMjLVJhY
F5tplfwYa7aNHxQV9TBmyY0dpmYyXLtRvm7lgpNpMsNytUzzwCzQM7eVOAMODShb
+shw/k90sSUh+VYsjTZYmskJ/rwC3kEDVaTajd2o0qz1bI6EueG6u6sLtG5ew2FQ
fHlj8Mq96XUz8UZPNSV2d1uDZ1rxnSvkExi++miBBox0uRw3ulCt/j/RJ8XuKlCt
5/7Cz0X4poBx1moE5hTKOi7TQxtSNCw5skzqNBQS5cv6Uo9XIHJeZuLq6Kwe8EhR
Keunh7HAyVCTuRcNreQ+ZeOlnSiX4GbxRoNHY59LO+TIe028fumLQ6az00jzU9n/
sldg5dfc4nJPzHiKK7eLu36HoNkE1z2q2mQ5lyih7AXctszlVd2t1YypBGj++SlE
u05AQsHMji7gq4vu5rEy/G/ivfDAW4GDIfmWmX5T6ib4pCSxvxxjzNm7tqYNzaLw
+2Y5NC99kp+qdslUZiE4CDwbb4PledtJuzV0//DzQpbPSlnSduf1L/4qoAUTAVoE
L1Jz4b9RlrqKwtq7PtOxCFI09CgNqG6JrJuLJNfqm7f6KlctY6sOqcQsLbr9LZlE
thJ4M7+az+M2UPFRRngSlJRkGVmTI0quVzBbi9CN9vwqTrL/r+TxHMOe7BjqGdAN
T7nJ3Xrlg4OLdYLJbw8xN0cuSd0+DXlz/naGDZQWQMOUTHGuQS5uCuyOJVWAx1FO
Su/biQTFrOrqpi9QASYTuZtg2yfyPP52jJKV5MTD1PGSV22TjV9yEG1tZ5XII03U
UjkZkOOZoR8L/I3nsVwFZvVA0r8V+g2EYyxJniXtodJSP5L4CtnQlppgU3BX2b2V
xKAYqMd9SMRdkA3lcNMrmCICtE/AAuN7zXSjC8NxViGLdZqPeCCHR5samydwN7Y6
Ap+pRFkIG7dspwbZjItdKyNyv+4LPokX9jLtAHt2GNJDm5fKeDvTrElmyFh1/ofn
WKrJMwwIjH/RL/L6phAU4yRYqTPbu8vpHTAj2ek9csxN0RDbLjMyMf+wU6h1pXws
D1mpdJCbYT4MZvUPYq7t/DBCBsMh9Jq07gj+YPQ3FlmM93GpFruggw7PxUtMO5GQ
RhK30FXnV66men0dKxqxliFUJhFnMloRvLEEvyPyu/0r/JRhvYatgJjX7g9rDAHZ
KMmV33frJB0vGzZn0rorlCkGb/+9a1QYyZrq2SKp1FexDYn+EnnGv1ee5IZXpdhX
XiOQ+zymgJedZnv4uYEh1WJnPjYRx/vPtCvVcyHMXpP7QYV3sblub/MKecGaeltK
xfsFNSpJzLMffnCTonU3Poy5OXy4a7iFt1QS/+xdGAIUxEv1j1Yqe0vBVmhaA4kq
mDfw4Ei0UYayHitPz6IimhlmyrOUQcYV5rJJneSz6Oa+7qHKFQSISoPYXK/QoQ4e
Yv+jprJP6y1W7hhysPwwK4HqK7jUFOdOEYffyFEZlUv3NtVEnDDFqD76j7ERqlML
tpxkMVC08jwkSTrRnZDZhSDNy+tekwG3lpe+lSikjpykLnYsA7Od/lYy/85nBIpE
Mf0dlwv/FWiit5LkdFNN6NkZwjjeSgItPGITl4DfbVKsHYiF8nP7AAhtJfETvZy9
Ho1q3pEfbdAYvGUafRVs5iXmDdJ3FpKnvtkwlctPugJrkeUPmDn+dvFQcnFXubrg
pQEu6iV7DIooskFQ+pvkNtucXJpIG+9ojloxhwj3U3c56Gq3lRx7ysikBrJdX8kn
zG/TBAOsEa3SStC8Tcmqy4y/WekcD1ifQQixzs1IJxpr42ksS5nJGa12WWHBCy9N
07Espmn/vR7EwsoActdYmB+Sw4Np+86cz4G+LC6wYkVUouRRnR66vxLRRQGFWeda
UIrGxlrCw7pEosK4O4OJesXHmh1fvFqwNAhNDoroEBrmx5J48HoH00DL/jSS43XG
OqQ/mY58MAhqpk5yQIXD5+wRpkMkrArgp1xk5xT2/Km01wi+ww0hW0n7+YiH/cIt
UR+WgMcWMe/1q5/LmjzF8U2r0VdRyq9hv0nc0rX953TDR8Od5rsse1zkaJ40FxCl
U4F4WyuuHug3WMveJs7+CeHrEAsB1f1Zj9UnbYyXxc1+bdxcdd7XHGX5ckAA+GAo
wq8StqJhTqGnrklg0CqFbbfg2FViUMlM6ORCV54HZfCQ5W/GcjOaRhSNanBSB9E+
79NScnX3Dnxwg+RLI4CyQg/m/Ro9mCPVJjoNmBnZV+FLvRpFZjTa3dAqnDf8+k9g
hAPqCi6YHr3y1Fv6hQmj6yRMhQQLeK7DUAiWXMsmTLjOh1skK9aG9JHK6EHFqKgV
GXio6fPtdKzCOxB78JAd86+211y2buOeOtCLiC1rAATLFtiN/JgCP/BfKi4SsHGV
ZcOCV8iVA3Rg9tow6z6BnFgYblyWSBzJjI+aed39Y6eQcK76jAQ6gfhjRQOXfpIK
kpxeF+W2WkjLLsqiHiUsKwuC72tMUmtv09x++6H04OanJYn/5dGGdOFlGIdDxeDi
+q6d/g9+XaNtQbq/0kXJWm+DQwFxe26i0O/ZUy95gNRBHBQPAjf7ZyfC0Gjr3ceP
LeWcsRcDBVp8zRoYo/bu/WJJZaEFXh2VG1A90bxj/y3uQvuXaZiM2Go7fQhQyNWp
tGzP/E9+yDzAPXjzIm/5C2J/fIVZ+r41jCcbEUJWpe1FsIhU1FPlxajnoa8b/8d4
JCw4ad9dXcZzle0HaTe5hzKjMtDRMMwkBy2lAp5k9PR1b4ZBAP8OoIEdtOAxViVh
QoJ1/05NVmnFkj7xzxwwEya14Wds+o/TZjQXPZfhETijvQtDQGoNXS3pOr/hej1c
0PHwnJgsjILbgFj3BEvLDKrwaf4MHLDUxbHS+iYyjlnzi9d65sYY32saYA3soIe7
FawrbVf7OTqOStWHRS11IkM4ruXrVrK2YHDfM39MvR0ibAwadN0crtp3Lr2nimcy
o2wzwOmAOAAdbZjcz9M+gWEWaSnlo1FsV0F7II0LYydCeu6SbFuSLDn0Ti9eBSr9
EFKMWZFkB0CY3yQscKFUrWo+8bSjZoJtpxvLQHZufZPKvZ1iyJUHNdavrPTljYwT
tTFPkfPocnsi9av8wKkQ1bF5PvNiykM6dQFZn6Y7RcMPFMJb+q4CXBJ1SgUDEZWm
vDv1mArFo822vOW8kPtNLxSTSytObWCGqz4HgXSDs/a9JpcpdoYGOmjUj8pjfY7a
8ZWwUKtHSHIBivwybDwnEPXBlNeOEWJq7SuYRAe8s2ZrFD5VIVNK33v723JR3aKb
oYBWJOKxTRur1f8BTL3J9JkLjik/XkRcPz2uNj+4BALnZSicshBknKuDJvEGLSvD
A7TjinhlStqJEPpWRfT4KLIy82ShbW891u4acKZmVssNL+wyDvM9JFXf6cc334r5
8s/74TYZfQHK/56rf846qH/0Oac/2y+9meee2V1ZYqmUi+93Abg6oYBaN3YsYG/6
/n292ZMhrfEUgrZhfPOglxqe0B6QDmRDa3orN+PiYrRFJ39EKjvQv+AC98ApZxbv
F6tRFBfM27SDq3Qa1BFeafA/7E3QvdGYzCF68m/9QgI47/AS5+14xisP62BewL5d
89SrbKgsXLinJCkD5mmhKF/qjl10UxylM7k0aWuK62dOCTpKZ1fYqG5uIZIjsskA
3KrVU5qE6z1/cD0NdWGsg19yBpfObo3rfazDDZqZqdUHIfkus2AftK1bITXitkbQ
7yzGQvpnu7JLd1Jfb285/rDTsoFyhZ/aKpHknMcNXMfPZauTmp5Vf02wJ6upuxs3
X1FUWr6BRHl3Lt3LoDS4E4xWmk7FP0O1de17mi80dBnXqZtuJQD+5A9qIVXSOLyV
d0cOChnjVf2TBCpK3tNpM9nukpWTFsU3DmCH3SorY+AgU4KPtO3sGP+57Qiw7XiB
6NLGibecmGyZX7ki4XymABdi1xydG1w/lKVElQxwLUqSSDAFt0ZmWkLmtcUhatXJ
wU90O7/SrdSmCKrnvjOqmQcO5jkJ2N8whIId5u5XCaWeiZWg7iNSkELTWhMHlqzn
u1Lwf4WoYI264dJlA9FFq1922+vbinfLx4QM4h5W1/fDDS5g6i6z79lZNE3Ag/UE
JIrmhcuxFP8qqkG5sY63fCSjfQYogEUfAAnKPpav98+WbcyRTzx1ThIUhZEbROoV
ACmpb4/DIivlWLkD5xIJNdwwtS+j5wXGf/cdELcRkHKI+FUql3jSF+UMpmJJKYAW
/Sv+hNXwHp4TBC0F99Ivuvk6E3kSJlROM99RYk1qD+oqJIl880XB+Z5mlAKEb0o2
TrrpiTUqMaFbqRqVWATuVoDnW0o0+Wtn2oXoJ5hfEgE2OdKOx61PIAAx9koIhaO0
UQ+Tp0dh0iMCbQSLQJQAA+myPwmDPiWIGY/ft4IfSQFAd5F/nTjr0OJg0w8CEEJI
kDZnfHT4G40jQy882FHhTwfeJ6Z4R9F0S2SMDhKwCXd+u2HKYHcVP1J8fA4DR0hn
vYh4uMdFkXTYoyFmpfxByoTbOW2rw65XGwXHVbYBreA25Wc2tHx0L7nZbS/S2Lms
J5Ic40/fJfJTyeBvvnFPIQAv0/3s/lAOQ4Qxr0x9ZIJyGIXf2HFOrqpVGEUQoE0A
VmeQOTvYOk9qEdDLCrCzmVb2E/K9PrMeicHT+pVx3/9RWENlmm+EsNUkwIt0RzLG
yz/M3fYCK4W4icqWN5kN2IGwkvOPtEnHfTlrRnujMCR7SzmgJ9/KHhCwyQQqLjW2
MMQSL24swgvRkoRHNI/jhCmzo2EaiMEZl1viAQZ1IZA9rzEMPt5YOrZs4euu4BkD
Z4Bg1N1y+C7hnDquNpdumnv9YEzzz8b6zQ0Ulv+Gj3gYDVwj8IPdjGai8y15m/fd
8Qde+lASYGk7ph17rxwbha+IcnwQ/Ngb30mauKjVu5Gx2Ujk7VQa70hgt+Z8hsju
z4DnqXIxgQvgPZXOrB1x3RlyujFGNpEVAKqsPx8MgUvtk1Nlk4ttoFFQB19XRfh/
ooC8ooRPwqJzR5CsJDUhHf41av6jLf09eizsxm7YGeXW/FXJ7PZXOf6DOYIjdYiG
qGioJ43CfatlLKY2xwUt8mGws7PhlhvZKvBwcuxpMw/hSgrQT+zgtPXOKjc4dCK5
N2wEomZZ+7neU2kSH9Vq+2xb+vHJqD+DhqHMGZ4mcUqF2nd96LSB68oXYmIjHMx2
/m/mvHzltP5FxuLEjF6fypVI7GC0bBVbQA/154/XMospVWPU9ElBsg115aMQQ7uI
RaTFnZQv8bZLswZFvFP0wshTzlMSSiX+/kMML7UEE3sVxXRB+mA6k0YRbGpFiJ4V
NiMajoap+6JeqNQqXMTJMsv7HoCVGzCGcDW9T49ys/rrQ72O7qkL0xfx0gVeIZU0
FdM5atouOT0nVQUoY+MxzdDT+VSJSQY5E6TNCo+NJELa8pMyfkXBpxHvluSOuLeb
3bUBwpUQJxZSjdcSUdEArxHKn/2v/m5WSxBokgr9AVytGY2r95IaE7K0TSW8fH5S
g1lhKX+Ay4G2ynew6XXdj0NYYox1uOzQ6zTlSUHuzVXfGOuOacd2tvin0/eTBa9D
`protect END_PROTECTED
