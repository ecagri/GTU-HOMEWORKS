`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jRy8n4UML3mTlQt1m5Yz7EoMZyB8qKYNGCHWMmR7yhbQINVV+6rVaioWC2wJSIit
ZJ3QLgfd5LfWxRR7K58hdYJu9rbq0H7kYHYuRE1ukfpVaHCicbIoItreEr8knPKX
BEbbo6x50n/ASTHASZmiB35xl6rBHmI4gtd+myDTdwt6HY/rT4isyg+3kfl5ZEcd
jki1inV5uGEvbb4hOCkdQ+5FeFFFYvo0FyNmIwbDxusceZVoooEU/Gc2Ff0OGvD2
KD9kFGiam1yq0PjQwwDx9BCyB8KKgHgc6vCBOmPLH+jRwnMaJGd0yBMdaN+zKYwM
+3vDm2uiSo65eDNO7QLyDEaoRu5Qg4mra01wiTAzaeJCYNi1LJS4dlcTqWxqTnfJ
P7JUC/uj3ai5S+Y3cV301pHVXR3AozgSOUdSCpcbJm22bhOLhbSoRObxtHSNeU+F
HO9znUWyPAEiafW8eaDuh3pL0PQqWubNH48qamUQZBQVuJgS87Nr2Fg4AXzsX/b5
HLR+tQ+wa5ycUuWD1oi+kgE0M9aIxe5Hy/+Cg4ZtsIX+os2qpcmZ8c3ToKLZHsNI
LRqZuSYcsUul9WkDLy0kG65WhmEGEvNnHzIGi8yph3/aQqjbJI9a0Prqiygt8An7
wgM8unefPa/2c/ig2aNHiQTqekfqxQVR2nrgQVzw5KwBQJnAU/tGYgd9MQdawIRp
pFwyVDqvpFdpt/FACZWENT6b9O496kMGp+YSNNS581arushqz4NifIs+rcHEYOxQ
xy8EzjUnh0umx0RjEu2YlMFjD4EzfO5EAx1qaRzsU9pcbFBTjuWp6PrXFdshfJ8u
WtC1My3j7o9kzTRCtTTHp8Hodf4Ju2J8d6bTpW++HWzUZknI1WfR/Mn4InOy/hRL
Ysspul1jOs4YG41jieDmTRUpqbTCbuE66VbMYUC43GGXXWliyEK6+riBuQ33VAey
/oLMddqRso6+JIKq8J0o/OU8z5QyUj8u6UoG5RWGwzTZBCg2ftI01f28ICJQkbSw
x3qIqFahVl0+khK9DCKt2R49e5y/Lfi5rdw0hSogNaVU6tW3cY75pZ2A3cEM5R5W
qeBiAIHotwzsarNPSC7NNTIcyc3LCGqups2n1AZM5cQ=
`protect END_PROTECTED
