`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J7Pp5Jnds0445YEBI+3cc18BZY2b2BjlzwGhKcI8jbh7DTrpmuDS+J6h6hThuKKx
g8iDEcREJwJiPua5TF4/wPffwmSELqWhj2Z3zxDGNNN6K0oHrmVUoDHcJnUmEA4t
6QRGh9yfr0XGuNsV/ojoD0+0WvD4l1ge1Gjx+U2WaDSVyF4ZKtzi7hSihSdn3gug
xvk0f7PuJXO3wo7wuEmtJW7dZY+7L3+SQrMxbpC2zAvYHgnLIwSVTlP/Fr5RBdqn
M1hLDScNrLcA6wwo3Jw10JniEsb/kHuRuZbyvikkRZQxL41H/2NibccOLO/XIVFW
hXXJMPiRHZZ+Oj+t21SsybEbwU6bw1IF0uzryOXL6F3Dkiwdr7pLxIJR2vFUQq8m
p714QhSWB3V3uZa1tsL8vvmKRzm8jYhN4dvwW7s48jqeUdDc3bXkuKVSVl/+/Tga
Gucd/qgnCpw8XvNUcXJhUn9lHLi8adZPuvMwJEILzHwMdwq3LTbzrjevv0yURZj0
KTAdTnwKBIXW9plo5z956+Ni5pY3J/U5/7OJD8MV/jwh+MEY7otTLrrjg/rwRt6H
f4KCFoyMFmL8lYUXJbQWA6Z1Tk67qxLLJkNDEmYyjybsSJVPHXwOeke+Yv8ACRe1
QA9OBdhvEugE9Y1UN6SepKtUVUGU/bd+aM7YGotjmKGL0H5wWZxBNhfw5eWC1onp
jv3aUTF/zz5vW9Hhuc30zPg/UUQaLx0J4Gth5nyIUr916/Uog73CpV46JBygII0u
TTb6adSNBXyOBFwIhoLoUqKtBfwH9ew6GyicvQ63NEagZlmI/APr0dGfG7hbugdh
bQ+4/6G23Y6lbDhtGZpeFqPzSI1oPVgTfK1cX/iG/Qmes97UJU94ARkVT4NEs73j
h/sHzJKSSvvvp8QI1E+kZsMXvYkZ5XVa8Qe+OX9TWQ+Wv4D9aKHalGuJU4EfLg/v
WuB0EPMaAFie4EzzY0H2Dd6YhnHUC3/uv692nEOQoy9uAHy3p/t6vOQE8R19on5d
SOBN9yGfuohtCf7k2P924wVjRkhKjIgXWEzpd+jkPH6jW82lp8TA1AfsYuRz4m+j
XPCJXTbrKTnTEOs//sibyuaTSmHCEQVXfBcNyvoGlvk=
`protect END_PROTECTED
