`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RZT0VCNLNcSQOJb8PYua3ngOMkVnVgaadTtaYlea1PPXD6GZhN4tZkokBNfFX2f6
yAvYRIhk/v8A1p/LLMwKwHgrJPsOK3ndIy+k4mpjPM7MFIBJA5SU3PX2UeQJbtuR
F8kQw4Bqqqegfyig3sUNLe16QtUARIoBj7DN2V0wGdwP031e7mOr11aSrpms8Q6C
W85ntu/iEwtE8G4IeFaG+46jnMw/SX9EG8BPezw71TjxC0vO0oUMXkWR6xI1mtH7
9Q3Gt7ckuFBtM5qo5yWXirjJlFJzuHk01uBnmiqxcuXBLFBLJFSWcil+KNUh5zwN
ubWgUY/44UCg5TikuP1xgsMR3Dua5xwDxsdjGzYGR32lgoGiPOd0DL6rPOVUb3Kx
deByorIJNSxZ64V1UoqSxCf+SeAu1mtvFgPRJ2ypCRtmfDhx+LthHyf+I32U2862
fZYlX9tOISfCL6ju3iAPFqsrA21HPUIYv4qJQ3DfetURRC7s5/wY2iv0hlGXnVvU
CnTcxfXYXpDDBqaUU5cjzcWtosG5PUnPTEQczha/YCAocrElc8evzhUDo6KIPj70
o8XIPzrsGyrhmkPPLGQbEKTDZ+eu7FczjnqogHFN2q6Eoe6nEPnq7XEZYi9tgkKJ
20px+N3CQg60y4SE9WZdk4KYD/eyWfd0QebDGAwz4JvoHXw0KdsxQuDvmteCM8bl
ozSSetZ3KcNVtq3gxEqN6CUqnrVHz6/FrifTm+doAP9y8l33H2HHcMU6S54iKnzz
+mqIIvVBEMMg6LnxyWQrXSd4pEbjsH2x+0oBY66r+WLuo0RcIiSEnn5WGDzGzL3q
UajgUk3NADH73kn/V60qCkCnUhrO8Qifx1CGYZjRUSN2JwMslIdndxZ0NP24bH5z
4rDjGpXENNda/MnEFwxE13iarX9JaY6Bjuf7+d9chvfyxVkBk0Ie5cGs1nd9wLmh
J6H5dFp5W5tgSgU/TmkUJruwweV7SkWFy+Xp7yx32Vka1cw0XrHr6rE2zpe2GgLg
dxzox2KylNTVyYs1ydXHz/nwRk8II5Lk40EsLjWrT9KIENlLSZt8sX9L7zTrWV+D
NrADyjmhb+0sinPqzaRm9jS67RzWo0V/GwUefWJ1nPTY3hlwinh+3Ith2nTySmrQ
DX6aGHLV3unOyrbUNBvl7jpq/JatQMYYZTL2gJMVym1hXLMrxTrgDWYlqHrP8P2l
X7vhH5E3Fwj2segxuJ0W/lOmh8klFC83KowqloBhcvSOw+lRoHGCcCgjuU1W1umd
J26oBDz7+LmGa8strPopvNHf1NSY7wG5iNWxHxBbxoJ5Lw59Pk5kd7hisLzGz93I
FxvZAhOtXvUN6/U6pfz7Fkny/5Cga5mouNMYYU82t24ofVTP0gkIAlEfVJl96arr
KCM3jBkT0jJJPwXQIPLUKJbCVz9rECHrpMYpYCc1FcA4UIImkq6+6tDTZNgbWuKx
20nvJORarjU88gpLMFMZPWtiEnJUY+nd+78l0ApGdmZKIeskGLNd4x2AHwuO0clw
409hWV3R3E94nA8QUOyv8Xdif70dz+i/VMYP7ZEdGvS2fk0FTMBKn8EZhtMAYFvv
WkjFHq3dVJpu44uNhVQzcOVk3yBh25cH82xRlBuN3ByYIrk3ff8HGZVHgnS1UQKg
0cqlHoBP2D8491gKfnbZ4oG2T9r+oa26AhoLrSpXqUYpg6W9AfslohbpDL1lir6a
CySpXnioDXzuqyQaNrdEBRsFs4xRZJcXPrA9MalrdMqjeXX2J/gJ6/in4p2PO01v
L8aAnZp7bv0G6u6vGrgEUMazZYOj+ja9Yb1kKHswiwQhzFQ9GqONZXRhzh/rMd/p
qiLDCQXKM+WusoaEqjArtQ==
`protect END_PROTECTED
