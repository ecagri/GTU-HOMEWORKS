`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lVL1uv9piuCZBD5KS16qL7TDObdPChvhduFJr2m6CX3wh97UwSY7mCHaxmc6urK9
RJ/XgAGPLOH65Q0rnGsruAZfdNsaBV8Ip0aqIj/IBrnxAtHxQgqK6FxyaMXh/JNk
Nsdhkg31hDyW72akuHQf39lYCKzOQaYs/IENGLKKWVPwIfs0n2FbMlnmUKfXvHFe
jE2hICqRxvEqnb391NKUiwyVIDXD79TYZCUNO5SGmBtVJzH4Dg9QRa3/fnDpcxKT
HU9ZWcIq3rwaOg4aqwGLeR4F0O1fD3rcJSJTPJTZCa/xARCyirmEai8smnGFkcC5
Jubq8orc0rHlcvXthTXPzPsWc5LwGPsUcaQI4D6BE4vGIWm1xx7x3B7t27BJhkZB
hwPwVIQppg469LwtVCtMPpsNJ3eMZrQcu6o+7jd1jicRuwCtRx9Zi2w2PQ2P+SUW
1iHvw1lXrJND4OutBnRafAjSBj1HRVUNmWzp0UlyBmOcv1scWjl+IuJan5sbdhnK
jRsrtI9eflmM3rStwW5RtrCKgJUQydjoBSYscI98zzTxtQF+L6FVap2c3Vv7Tm/i
7egf6vKQcAaEuZsDsdlW5lHj7DdamJMXl1YUrVLZXJ7kr93Oxzl/BZYMak8u2y5N
XdWqHOxOwDMsLRgVV95ebaT7dKPXWnqm7LrEHPDF3KzH09u+XVLd7KqkBy4ANlQt
Qce7OV8gwrU39IlOeDXhq1JKw4zU2xj00RuYrCDXNER+6At0uNMYdu6YE4TWAF8K
trUcHLyoaPPNz2Ntn9p5CvEO1MbIAyG3ubC6SlP87R2PRUHuA22vFvqCn1CSUKR1
pEPLQUQOlXmJqISdUa9TPhntKoA0qZh+YjvMxckIxH6K8DwTQSu33NRaXDHoVrBM
uP137F6jVfBk7LWujLyJ2GXYBzBodjP/M3vjrGHz+K/4NiMhiAisRK/JZqIP48yz
juEE6fYRrOQuk47Ui1d8udMlRSbzPYC9TdPSy7ALLHbhVENejuwBLHD3ubGp04Hr
OH0PuUhqdVdHC1QGtAt0VQ+ehD0pmWWPWt2ckQb4VOF8A1aeQKrtD0QVnsG9VPHg
0GTSqIEFNAX+ma7nIV9tBY/ZvpNLvFHodmIqps96YOsH7JsFUUYcu/KC5JgiYhe0
Q11Cjs7WdQfSZza0fFVwbLRnrb4MbxemXtpMWV58Q5HoLnKwDJgmRPgMelmAXwie
CsHle4FHHp8NIZx4G4HGuATBl6+kR0FgCCzJcfCspo9tpdQXBB5M4d7MRbHgZBKV
LoUs2lVmL5NoXRJHCOXRPc6DRmIskMw43cT8EvbVPLusgtHpmFq1lr/hjvakSzFJ
J8v70ZjfAwTHxpFVYOSKJHjTblv6NdNWpWFgXTzNwAMwV1tadGWrD3BakJXfzojE
CvSL+TPCj2N9/fT/TdKSbKHPjmHyJ+yCkDhpv1IHKYb6GTdnvUc5AgRzw+TuW5zS
yHlXYFr2S+0mHad8j6kW8tyQyEFrnnpYdZJdJ9CxK7+RYeWwSVjMi7umgAqtFxlE
LeQ1MPo2HWb/vZdrxmI3CS7NHjcZO99IlrgfCprLXQ/xn+3To7Y15fWv9ModFwL4
0+s+MAsTFe6jR7JsBErWXRwxPcbR9S22GbsnE06GAxMwE9MO+1UGZvMdYMU6Kzqv
3h/Xz7WED6UlXqaFW9q0hrQhtPjWBnjVTAwNOOFPHccLA0GzJSnAIZPSVG3l6HHs
M7Tuk8I2vxw4e/jvH7l455yt20/GuNuwCfT2AQrkrku0EwjdFcTY7y2UPj5abJUn
9rI6EIW47QxZErm3W1//xrkVKZYatgeFi9YK+Rf5eIjEoQLpi2fdSSeKiFmIPZ+M
wLsMwjt3WrUu4YgIK7CRYTadkz+6ntkx462wO0fFFeNCOcZ3vCTx6vyn/Xo0Atm7
Kh6yrnWR0NLu/bZQtI3SfwD5u31ewnsLD9KDpP/3lWKrIO0Z790hJz4wwxdyp4qg
xzgtcuB/7FS4EUgH27TbkBlryJnG6vue6LEexHMUnvBJZII0UN4G20qSo+CRKdph
smQOfvb0R1YGvYpeQSFISTZXE+Fw6PNIV1LuEcjUX+i31LCjuiHC3/K4btRh0dob
Wu4SdlAcPYVc+M2hFE4g39Tteu/eXTmaM1BQ2PDu07/xuzlSbCL2Z0ku/1bT5ImU
OpfvHezpE2lPNPMBW+EamlY7N07uZuYKAnxFjF/KR9pj4F5DcMpOM2Ez6yVII3Mo
mzNNw78Lf2uAVRCdtbDP+HVWW9mX/Tnl+Oe1rDa/8lwPk9XJk0hb270yIyrysNGa
XgAW5TPcTuBZipi/BTWubbymj4vWYU898bjVHGz/ltwHfwH6EvxhHsBO4FaFtykV
MmcKw9JfINjL3dS9fMBtftkipppslPcGkOCV+eNpwZREZa7yR/nZqZautLUcKhy5
R3rAJoEd1DwgtQu+8a70b9niI4spOFeIT8drDuMy6/XVUCKivUNhzfSvQKYGgZ3p
htJovJnSj5IoLB1W8+At0oPIajIXAdxnZcg5EKDeyKI82BAscIiGi9Hz4kTiz/br
b/Vw2bsqOOK/SFRI1j+addaLWzXlS2BEaKPCx8f7R4mF46m671ZwzVw+tEUr2rCu
wYIaH7lJjpxTg/g7SbNHrlYQV3rHJeUr90mejUSXnI7P0uedDLJaCT298Y0KkWsM
MgQEfTVREXK05Jg0owhsmTHKitzkb9VQ0o1z+Iqw2q/8kk9BM1+BViViVMFUIzfw
EDd+AqxXxMyhpOHugOntoj7zu6qtVekVcvgroR/EJ1WOoceTmI5o+nXXtEZuvFFB
4JiBenGGI23BOo2eRpKJ18CdHqb9E/mQ8KQTdFPjDhskVg9YndlBJpVUKCEF6KIO
trIBaWx+K5GHSt5E/8kE5g==
`protect END_PROTECTED
