`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8y6JuizGKtTa01CTYxNt1YDug/IQDcc2JygacBa2LOF5i7DiVDZ779Nqd1HOwG6J
qt9NsgSiUwEpAKzgjNHINldUceStOvGI84ei4teQeK/FNUNuW5yNE1HuA0wQIila
hcbbQb7J6HiXUAOorbij3cJdrxB3BMYgkrGN+WR/RRxOIx9PHDjALmFWjD1jm3rj
aUxo9aNeHHyZ64NBLmC/8oJLlp0qfvIxJmIv3sIEg1rhftwiRI9ZUmBkyzJX6THD
TIKWSPQxCBdXc95GS6hrt90srLHGXTa8nD2d7+77l4RHG+1yVszG3D0L0hLiOLek
yvi2x9Y+pmYZ7wY+P3aVv5rj639Zikppu2wIyzShtVM3aXH51noV6yFau985fHKF
DlHv5a/bR7SBQvzxT7LJEh1vc+MmIPXs28HMUKemfhYVM/Mar/JDqHvwm1qHEvjL
2JFEUidAto5h7yCnddj+EtXb2eB84QYMcyV18tX1EO64stjx7/Chp4oM2Nze3IUB
/VnMvgNIl8i48CMkhcBfrKwuh5TCjxam7D/pH56a85w=
`protect END_PROTECTED
