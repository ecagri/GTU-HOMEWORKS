`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
USmIf+MtTPGAR3g23L5gjinmrGdCHLB9dGNztlLmiEQaQN+I5qDuF0DggXwZurRT
zJmTxFT3LTqyXuDl3EaPhUoNKi/FV0S82oVfiTaU7GD0GIZmrxUaPOty1GZu0eFE
M4+X8jIu/MIfd3VhMqNDG0gwoHceTYvt03AZivh2ogrWVD0YxAmO/49kOwjykF+P
elrUZnlhy5alWrJcD4eVV6RUOleAo1rAqh/Y+4XtLEaCxwmVoq8anaM9q1PH3jRU
NmW22Pn/7qGkb43Ku0cc+iznHMqVK4USBQAU5xa/cAqQ+SO3PoXfQ0CaqkZZZnhz
wxfwEn45ea71JCrzZos35qubF66yYI2zi3N0vKhIJdIXytk2lq1kkVy1kJ3PlI8d
2E3nkgmwzTVTnvw6RGiNBguDezqLmrg1UHolifoivGLrWM9LAVlnRDDf7nPPUMbC
WUxN7RXS4gFQmbucdI/SQG3WhU7v56WmjqIaB8Zc8TuhI/xzRDOSt/c4Zyi33bu/
cipJL0rEzUXGxiKySIncRjQd7MGb2HPJ7bWMTogZQ0zT0kSitdk6GmWFlargRZnP
vy6yz0BFTP2/dyWQm0OlworOT1FHYzzuai+qEDARxzco8q9KlHqbIXYXa4d9uKU1
OsLpUeBqTw8DDv8/jeQNHjSVSArpeaB70iLKu+o+9k1bl8ikosnDwwXjMv+z0+It
2wJhJ+05msICvqUMmBZGJwFRNXXEn8He92wZ6NXVIfQ6f7xN7Yh2SnNn9N5imgH0
rALtXze/xcO4zhc3Lj0w9wXCuoJ/RPE87E8IHbNGnL9GsmckD6P+PVD19AfIGWyS
aBfQDSbhv0/d7XIunhd83+OrIDJUvi1EW4DWk5/PChOKrUuEj/AmmjWptalZmkbG
7M7DvMazEySeNEHLhw0ZRZD0wL9Sc1G9yR1Cv3W9fi0zX92w0XLKFTgZj42wkv0B
VNvjxws/qCnC+4t6gdv6lc+NDQctZdCa6UvOH21y8gXlD0H7tLQcNpa70rZt4X/E
htHuA0Ka0iMXSOH/FcODuofXhNSzuuwHCCBLkNXr9zWoEJZ6RaAzPQBdWgk/Vrhn
wSZZvo2Fb7ZUZfSuRM6ELPioj5bOZjwOmD4AyW2988m/Mh0y5vLRgAD6eiBNKn5d
A65VgEadXPiJ3oo+Tp+w7MY+NkGnPTCXQa9cxFt8lHaY2hZ+jl92qwIn1T7ZBcm/
bdRc8l31fdmywVN3Bu5dcfWduCILn1jDlcgy7NBGcaiWsIyTJH7nTTDJxke3XW1S
c9jx6Td8oHMDMbwidAfAaWusAJq8DzloBDYecZNPQkQ9FwonSdgUmR63tzgBxICO
dNuMTmSa0Tv9Q5T/v9XY3VkMiR7+Qb2Ojr7snKa9Dl5WciVa2pCSfsAtJb1lP1ff
HL2qfQCnh8oVOlQ7a6AfSC1lLxhs6ea3IKnMbub2fCFMur7yxF/zAMjpjWr1jC+j
RuAoREvnRBBXnoxAoAggFE4Tm31Rdx83T8su6ezs4Q5mR1Vn1gKOAAQUV0CD6YpR
YTzF0QOJJ1AwmDDY/5TE8eM6wlTB9/J3G3S0+vkXsr7E365ZWm1TB3RM4M0eJO2V
PzDp7Vu/Y5IAAPfremBovrBt6czhXnd6Vs8L3SAhsWZATjgmYPNO4gv/ovY8IviX
MhouVTi8rslBVuElgLViCCbMVG52Ahnbl2vElK3Dbtq89Hj0hHZVbNg4hhdAdy+W
U+VQz+ENc0IisM6AwDtHNjMSjzB896qpqeBRyNudmSQMABnePopYOmQryd5trSIo
ZzZ9UsP0mN+ulVLnt1Cnu415PGs9ghpZj0RBLIz+OCZXWbALEG9aLXmQpc/hVseD
HE01W6iqK+P+k60iPjE32Am2O6Fzqtww4vm7BP3YkSevDuTEyAhIW3WJD457OjlB
fTvW00ixbVaGz4V5bLObgc6SCX/b7gBmM0iCwq30eXejCZMDOgEKPmzaw00toh3p
jTeIfY5gscNM+06YU+b7EsqQVaigDcNps3frBcigIVWYxrSXUVL/k9R01jz0Cydq
fffZXU/eYfXGm/Jopa5fJc4zN+JXmdUUkU3n08EJENNpfm8SqJAQ5UFe5S+2+/9j
+5zl4NK8rR2X2vr5QCMAqxKNPg9QrI25R5+liqv+r58qSgFeoGgBI2B+SCGOVd8h
sRuDulKZC0Vn6nSOu2AnOb4VCeZW9uVS1dTNiFj57zmeRGBHnmCW3BqsnIRAom6v
Cx/v9WAeRUEn+bugc0P4z2fPhIzeURV/h+x+OxHpZy3RG7nw6QGyGE9xrt9waP1G
S2ZFprXqhwY9GFj5i46uvbnFNJQiN4ueUSNLv97u1VB7YXsHEz/G1RbcSXN6Uyl7
Y0yQSSBbiq1ZaL486BhfcEFwdjXQ4F0C4gKDXomekpb4mEtqyGX0BIAfCfDkuO8z
tUDOtIcr4yLjBtMWA/I9FCvxzpBTlAAEhAJ30K2E8JY6T6VidxbSkTAWG8wHQHcl
go7OcdHYf6dH/9h5DbzzgE7sG4ALATsxae4b39mZzbV5IB+HDwW4IqLDLmGGAAzL
hrVvGN8AVh1qgEDcvVCCXKUc02maOTyw4ofzJc7LJA8pZbl//zdWBtZiGwj7+2vO
oxWfK3cqc4hrUG2XTx10XuAOvdeiqNIrI8RXotv67NjhQ0G9+oSKhhEoEid0UZ57
8lyrUe5ungRofa2itfo7E1Z3YiXtJRZA700DeonX64YJa2nQBkG4awEawwtX6ptV
gDM3/Scz8jQgJdQJcKEwcVwYacwTw5bYPzlhJTyyksYFGoys9OR7ZBXhQxviBBtj
dje1l6Yu7ppmZkl94eM7uXdorGwezXxw2uWe1NXppoIKTvj0IuWaYN28ry0P1IYe
Oi2k0g91agFn6vELKOKEcfa59oM2QRllig6yIHzXb0XaEdmypwXPUSpfTK3oHYOU
c82XahZw3GUxygzUy02WTeXFvp97YO6n//dKkBtZZQMbJR1OuVuUkZ8p+UOFvF1z
0/UWxQ8hGca9F298oQoTT0QrhmafwqYl8ze0mfV7QUfq2KQdAar5vJZ3rhoU+a4L
yZzbBBjwmY1Miaq4qHMHP1C0BIeveRU3aVXKBTj6ppXwmMPYumIzziKbzulAmxd7
butAUcWOd7dCKdwmmOf+sfGKN2prEvI0k4Rg1m6QglKJqC/ft8tPl7uC84O903Fu
tl/Ns5LN63aqso2yk15jvrrrZA+ZZkrlOXKb0POShnOeesvWta3iU8JZJEezbv58
rWs2hW4pV9dY6mCk/mvsPAWCbj/P4gORg4G2YqNSkBLTdIzsQepQIidKyhgvmORB
CrZk6DvzIk0vEcj9bSiB4/X0zuzld+OAzbnoW/GJZLPGSnszmMQ2Typ7gQ6lImuF
YAr8wJE8XRVHPxbtpwGVaaKqa0PnVMJ1HVOiBhsjPSw4KabjZ2C1vmC64jIKPeVB
TBiIpWGG/J0xntBsgFDWagYTlp7g2i2Jq1CRl/u63fM5ybnlIxNWEIg2snAhl+q9
G0UWD2g/gFagpK3RMl+vm1u8ZXmAeL9j9sgWYhiHTkHmf1nTdEA003vi3GcbmuWT
QFD7KLtH5xk+i44Dzo5+I7Hvzli/78blpWndrLhyFwk1kt3OS1PY1HPcFmbEL/oQ
ZlYRH6M9pduv5EV5vZjvhRFAt5OOAweogpeq4dYJ5wkcaRQpYv379q+d1SgeL2J/
57ApE3o552OhMt/PVQbDXJqX72IWHXlmSuczPSrCuBSStWzbYJZVspUN4NiTTfZ4
M9SGRIv/vr+ggyYMV7lTmci9L5uE9ZZBkC2l+d5BOAArYIP4DKqRmp10RN8TGSTK
6I3Oxv8SI+8SY+0VaBUGlgbLYnMucqVJ5wIULzGo9rfqxRk0DckNL7V7dG1Nopqs
4OOGMEoIKoUDbWKnMJMtfjkm5nXRFoe8daz03O6+NB0IHoHrJtv+NH/j6sOvc/4T
ii2sWFOVjp425WThF/2D3V2mNMMAcsI49gcHhj2tHHg+AD10i36eeebcDGvrA26R
MH1HY43q75qeXDEisV5DMjScAW74SATriCgid0S45xf18KWGRxb7Gmo+UusxoRib
pxkakC4WFOrTOGxiosGDrjsm6KN6B4Vw4LPCYGhS5m5pFELLYTDC+gUgg1T4H8Aa
XCpXwy+0IF8aXWJ+0lvNNWO8uxWbtLfBS0Jb+EXJF2/sXwUO0EM9CpHrFVv3ILXl
g1Ow6I/QRJvMHXQ5YRCd5q4sO79hZ2u/raaJkwBbFyKypc0NGM+WArHvymYz+S/2
Ld4vTJVt3wNVtgBhzX2bIrLAK/giZN8vrpai+HQiWO1Q1NR8JRLbkF3takZHuPZm
Ep7aHARllhgJcfErlI12mFTrsRJbmFQAo+xeiV80hK9Kqt2+hc09LsYcxp+bWgeZ
CmBTFsuksoj0joCM+1rl7aRiDERpewNsROJrkN9HCVDbsvtCiG+K6GNiNi66mzWb
enEmiY0/fQnJ3h/XSjTVnTasyiI0s6K+Il/2h0fECMv7PjAqSvZu8uSPtkecqX/k
QJNE5OsmzU9QiE8wjZ3MY3FYpPmgA3GXe7jqc5vGs0JZiwWWsXWt9hsgCJNF+IEu
8RU7yuSTCabh9lrK/u3g+69vbvu0pJCGDwNDFp1UagzZACpDr7wAVK60oW4CEU+t
gHTtMuF1isZamrLPEF8cb0g5RquVozXek/sfwaLk7qt7snE6UfT8BIwmQNsuZIOB
6wZD87g2FyzSTzHT7ok8QeD6mUUyvwkGorbctziDlUDKxvKoR31UJdZ3Ehf3is4L
07bKkDVs9j9y456YlE73A3dUl8QKECfEaJ03a5FbRWiiTiIOLeP9eihnb4aY4NdT
ruZzQsJm//3+ggXfjya4WN3CatiXf4Gupao3ybbgM6kgex5JD0Emrm+uerHp0nAS
4kr4v7joEaK/ZnmyU2fj+6EJ2VFwWi4vWcijXQKxW2OrAakXbxtXKsrARug9B1XA
Oq/iXTKDrLpfxD2QJ7C/famiNBmgMVTMTCF8ZJC5JFyQQztbO9EKqTDbcUaLkj3b
02qGNN499sqbNwwjIA9PkIE5JxjfUEWC6oG7jB75Z1/IKdOR6+6JFHkbI2b0Dqk+
qELASbxqgSD9wieEiZEc70SSc46+6I4PKQuhVXAdzOpC7kiBUOeKd6NRiVuyamAw
k2bK2YbdHz64D2E9OXuALkVS9duaGoJncWO0mPl9ubJMfAa5320sfAUcB8r9ROqA
05SeYvvNR1oGDGftpY4QYXq/gWeYfXUAU6BEjQboejJ7Adi9ts/6R3/8p5gpTSZ6
cqm8hGB4ElL7X5wasycHkz4nH53TO6JrOS7f93PfFDf+fmHCd+NVIAbpv29AcdRn
cyMoO30BX2n6hAzEeoHKBFJByPqKZRw5Z01+zKHbpjIr6UCCpuYrbSxG75zoZbLe
RfD2/iPoWpZOMFNuGDPIgZB5a45cQONo0XywAED0WPYdxLwZx0a0Q7m0x2T9/6gc
trz2LbkeEc5HuSnb56VKjfKebzpwTe07v5Av44ky2KZW37nJIRqpVQqrgjWhN8Dq
Cky7GnP21I+dov503u+QHz27gWJGMXksEkli7fdsB0EBAVSHADd7JGrkUeRrrdM+
MFv0YbQ7LZZcnSvpV5ADGIkGzIow+RBt95pQcgLDhK3szqZ935PLuaUAY1kE+LcB
BRFX4vTaToafD5jQP614gLc0zgUihkk+YhPezLm0VW8AUXYz3hdgdqlzH1Oib2eG
+ziGi4TMVUMhrzq2HXBMHvS9uQl4KLboOTci+ezJlqEiEXIvmsxPhaHRtlIQ6GaX
9MQAUZlRGfxl817DluLF06i6G8Md1C1FdWtgGD1a0o//0eXDp785QVP8k8L+Ar6v
fxCCIBKisUKg+WlEar68ct2Kvz8CjLS5dl3WdJZxeN6u4OodGMsdfQNeTDIuEak0
KvTBa5FfRlrPWRNl0IlZPNMKJ8Z0m/WAGsrz3G0P++e6KeohT3hHuEK1GJFizO7N
I9ZlZJa1Fhq4xau8Gq3KeZdv0LXo8foYjzy0qKsaL8aOJYAWjlDJpfNnKPKyuluC
Y+6iEbedaNk2NFE53qQwNqBf8hsQSAPwGgiO7A1tENMrhUALs7WwyAH0Eci5k6uZ
Tn1GdYMT2AtPGyhpU7eRApJPutmH7fvsavDmiEK3DkecvepskSJplUUn7OCaQZI2
LKUAS+18Le46wgDaPZmo4X2fkDEGW+3zpc6k0su6sfWyGoTvZXNGkpj8sVBoMOUR
19eMnpuNArIgvPrCoWogKMmKntqAriiszuxPqtlFGC8wMQvejVRQ+iB7u2xrrpHm
GJSf338lMu/1rbvw8enZIwXorTPyftOpD9TSUHsDyKrjICFDTSMaXtLxC5h9wa0N
0/4ceSchtyLetj9aS1ZX8wmIadBYZvxq+Y6pUo32it9U2dQc84rbfbfLhBNldm8T
6ZRHN/XnITx9rOKvgxNSvVqWKKGly5YnM+M7R7PiVBzRO6Qf67JM6HDI1APX1imn
/u0sev+G5Cka4OgELML8+wmI2V5kzVh2+twZPHUzdHD4Z+Fe4j48mYk/37uTLodK
KGGsMpzuMqUFa6zErD3sbtM9ODGraHa+S6/T4+Y+tWiy04B7u0AQaCggteix7dGz
NTj+rKL1Kt4HpPIRo7QojG/UAwnLsj/s1rvRuRg6CRb94+Wt6uIA3XLESgwSjZG8
+FzyPLbLp5tJkM/Sh0hDvzaUuEfRozmdPiodfjc4uobL0TLaqe1I30QmayLpY08A
1gq1pIeRgOFnP5X0JPOHP9QJkuYKWtoYu8C6AkujsKPtfNXFNWuYtewqNUAAsFEk
NOUwYDvht1AXnbjYAhwqMjLKkaksqhvGQ3z6QRZOqOQASnWRe0WEYdHoU57aZPd3
Y1ogyRxFL+KfmDKwyyB46e/QZfggKSKJUFZVDcsJKO9p71m5TB+m7SCqjJ+YrPyH
UE+PvfRiPXLeOYWfwB9LCvsX9jYtL0BHb1vHPOpQ8Z0NvMeBbAJrlvNlew4fvbLo
GEr1uaJElmpovoRkIjM6CB3f4oxE4LVxvyYfwL/pdBRXJK63DoJ0WFSL4tTw70iT
e8XaFgRk+XhwKAZloH2Ml0zwXK46h1sEsQ/7stmVTYQiFJNMnMJ5EMDryDUjvHrP
LOjODscxT/TTqJmO9RZ4TEiOPb/WeOr06ZhfbgHMYK8dlbnuxH2/BXizJwEyLfQe
/JRIvWR8OXFwFVyctxakNVHmPFRvN3tiJ38H5EWV4AfRoUXh0ZgYEfaI47DLAyx6
QJoTKA4VP5kS1PpYA7QzImm/z2W6XN94KieExD1JpMTfe8wUPcdDImJWwoU+XSSa
AMssObkHrY0rQnbWKxQRoPO3Z4Cmf1bgRwEMdOR7xZqibxnatBwcw924oCN2nJEV
q/dovEhaX9jGyTNCExZyQ44YqdvLmzML1Qm60BOqkWuhhfQhqzDtwEAqfldYP2B6
+416A7AIBAKqjGvNbAzFG5EIJB6yhuGXcun1HRH7TA8RyvaamTmW5CrrBBgaO9n1
cCK2AFt6cu2pISsC5Wjp65ia2fpoq8s5JVNQGjG2Dq7nx17KTbCAXqwhH5Ifjqqy
xluLLlWDbl5066976uhCiDsX2DDtchfJfjgVDRK0vEDSeyk0QlJNhZWuLAZoASNF
d1CJzbyczIfkFYplWyalhX1+myjeBw9NpbBtDMbsWwlZEG4/Ggzz2sCaEwlZfAsI
NzCjdUrQleg1oZ7T69rvnYqzZ97XPMXgCQcIfsY3aRCdIOTYy/zudFW7+MrcAA6H
j5ED82cOBB7D/thWarqAumPmbgBMS+Oi2b/H2ydMY75J35L1ILgd3v7h/mhtzh1H
vSDFZ5QQyi8T3m0O06ub9PAc2/Yi0rWolQDZduToMV2Jp/3wVSJDsUct8E2S6G8g
NliWBD8DVgfsqKBp8e7mBKysInoIqeaUiWPZhH+q81npAgkNTlRb1UagDV5eQ6Mc
fatGqDD9N9cSC6sq7S0+8MnRGjLVQ3j13e4q2p+o11kTuiAKxBwOvAWFvlj+9aqM
ymampb4E+HwoWuNL9ADVz1ZRrk4OL6WA8aVj+e4qMRQ3gNrZpgN8NPqlW6t8CHM4
t4us94se7I/iguvEwL/1YugI7tUrH3j4hZXl+SGM5Az095rFg3WA5494hHF7hxyh
kd8skoKUwjS6neGXdfcsAlJQiA8MK7fVzBOwF4ZwK+3I4Js6eHJthWLrBcTIED0x
Vtfl9WVtJPMynSF5XcceUg+hGvz3cZGg8CnXy7INEgiRLGl2+/m03rgwzQlpqk3+
NxMUW66apKmdWkhnNRwmf+5m8Kjvob9aGYOjSWrGiPfaOrSMxAGmkBUFy2SubtSw
9SxhzHHwb3wYJk6pYhEv/F2BR1wxYpm1AjpC+wecdgVBd/3SYrm/ii6mI2rEhbBM
l0jWOJRSlcMcHjkFBTjHQFv+SqtDU933xfCtxJPaPYthJuNSt/OHD39NCR8+GKC3
T6IDDxFEVjq55WAjDTITI+mjVb2R8qbLG87BtaGMndKDJVncsFDffypL6PJyJFA8
4DS0BbRL5AdPiq9PZ9JIOZX9xUx1E/BRFEISGPt1l+uMHLZ7DgEbNvIGwgZrJ0Ci
oIXNcRZdpOeidIuKrU6/rSVa5KjFM6GsBeCumbqEGy2BFXHTUMDDnQoRhCSs0EkH
I+QGQ2YOMVNyu7uNm/+BHEgYv8WjvebDHZVscJ/1pPt8wmvPSkauoAoWWWkht6ab
sPbUE2JRXuXEsqV9wnL/SbeVLCy92WAlfE1e7XuhzAYl/aFgmiQZa5DBHAQJTQI6
H56XKL+A00pOFB4r2hTwS0fTcRDahKvAlJKNC+Dqa6lwJyqyFFwHaI6i3yp5CdZM
WrsazKsexUJyl2mUOMbs/XBtvyZUHD7goTGrAd+6zpiYWLzs24BBluAeiLNOk8cq
n9u6A1S/5vieqChy7p5CQlu1fOYz3Yl/yu+56wLRlqfq2AVIHQjN8nNjXaSQBlY3
25hiRlDC0Ngyw2Sag9GnDevzBvDU7+jSdqj4qMHVuGjzskFzD1UECYZnqsL+BGuE
+z2mbB+Fkw80qvLrSARVCeZ9JUxj6iNsjmI2ykFc6Gdjxy8kmtq1zEw6Y7a85l1I
iX7Olt0luJvBpIXbehLAdaoV6ZCkz5nKKHGp1/+Q40PFeZ+VFHubdwEiJX5Brdzl
8G2c2gnlPOjV6A95JGur88+n5XQJZGhsPakhNY2dfmB+H6lEmqW9u/y5hrutIq55
Klq3nRHJNC/fLGxQtf2VNRS+/R2C7WdDC9lg/fP6nMQ/BZ6+FnRdOY75OY3FzA3F
Xj61f8V6ipwi/k0dPpr44ojLhtAaBZdFCH0VYR7JQWBJ9d4kfsaEvD9KyqZY59WN
kPlSjeweVwzmrygaZhvrhDufiRPF76d18bIeqiYm8i8hU9NWlbPMLhArrF2Lf+zO
vxV5RGARs8dKGB+Hz5YHl5ioKOwwAMjFtGBjszSa8406oUG7tv7+opEfcmmBIciY
fQ3jSO67+o7ISdQRTo0trspjnZ0OZ9P0PYwIbFkqEFImXxqZfm11jw+RBqCLPh2l
kEOE4mH4GZgaMz5IBmU2Ewg3TMIA46byuBCy6l/VzqQz1wQjL+8+Hvezo4HcGWXx
RWBEHP9/ROZP9EMGijPCXa/N+RB8YtSyeI873x7YqDPlgiojweqMWNq5/vlPi5hg
kdKTJjML8HK2zg9wvFaiQnZb3+8gMwHUmre5Rqedzxqb5633rAgWVIk4YSTP8jiQ
52TNaFBHy+wKM2xLr6M3ptKvtCuFZBuHGtfwYBArmWb6FJjEU2ECCICmBmPVoNjF
OFgzmyfvrU6HiXjlEF6ctjI+ajj/K3C5qpsUzNSxWUMo+m+AKloTg/q/Eijd8H0w
QodofSFgjTOddJbVCASdnV/bCOfCqJg2eNrr+zuRXGoCJRBE+drUDV6RI7AABTeW
8vtNgqZ/P8Uz3kltA1qLCMBW7PPPpotQaE8jMIjrSU7zG+KRRbv3id6niD1mq8Ze
MDvmhQ2F9U68uHwHcXAX3W3rtYkyNpHZvD7ven7GYmj4QXPxOr/DTkjueafQuJgH
tBDCmyP92DCnwRmsFuiS64m5TXWGyn9LQzhq4pwBs93xllNqYYlWjlytpr+VswqU
0v7cPWrbS1f1NAUXxDxLNiQYXJwcTjA5fy4HGTnQwJttyqbiqCPKFuZkEx7PcXE+
jhesmPEhX1XO4Q26i1ibfDKucx9BA9FXKnZii7KIhzCopg7JWXpl/YPOZpGMeQCz
hYznOzwCpdBRyHRu/+qaEyXyVzNKno9oOupsq5z6KR9yuMdYi8ppI9jD+neK+zfD
3cVggpMBTVp9ntkOFcT+wkJAZ5TH2cpzeF/BWcGFxSsdvakrU7jlHVHRNlUpyyBy
NBOLilU+dftHu7HWhtu8nCNhhOAC0yZ8Cc3QIbIKsDSm5X62XQAaExhHap1IMAyb
72TcAzfNnWDuBnvHrQs7o6jpgF8zz4D/3isFx2EvGgw77Ddwzm12BgzNDfTSHpgC
2jZEXZvFult7k20Rw/VmV9SyanJRqxJloesqIeVz5nEvUv53nCSJHfn60NxD/uS6
JwM8zQXWSPjOZzJKmOKl4UkF789UNwnaT/sF0ubUtNnIwNAYla2cgVpG+Oe7bCa/
VfpKmxWmBbX7nYydqyzHogueuztGQylz2H/Dnpulo+3zsnZB1/qV6XqYaElV6uUp
oN1hitKgmjwU8doaYnfgVDbP78+B9rJda7++q8UvJM8dZds83XHSnINhg4JIntfp
03qPjSO7FLdwKc6YAfuTALDmzGtP2G3WMa+TKVTe934WFWYi33t3c+0q4pFiA51J
W7cXNqF0jzLjf+CmX1u/ums5M9WvA1ZkhUONXaOJX+Z/UNpUxzmPx/MmzhI6izgE
goGz85gWdigJkBzZkNY6N004L0phRdc4ftkkJXyJFfvSPaJRxCAPE63PJ17Kg+WA
ozOZeUHYwkl+vqHhfUu6eh8Nsj/LHFUjaoCQ4CN4n5owLQ9tom6EZv+fDhft0KSq
u7RxSei/+AzBuH/e0s2qaiJoKe5UOaP0O29LF2xi3chwcjpFprY4oE8qjbGGjbyT
YsOpIgGbL3EQ1ovfnvGjF8w1yFu/UVfmfd2bKCiqTgkSaREY6K6dz26Z3RBuQmfF
a6N3Z7NcGq+0m3BHGsTrAJZeoxaZBoLBoA3+sxrMn3Gjc63CtcA4KOHL21FUt5jO
+DIcweo9PRUNSzOjdBK19K8pM1Wy8l3xh9BCxPfGzmFkUOyFrMAefQgVfLQHZJX5
s2XKx2mUw8EYidE7cW5/zIHMAneMcWs7yaV9tGQ8cabhxuEpcCAwaxKw6KOKsdAJ
sFqOeHBP4o2e0M+nZ4I/Xnl5HWfYvANjdRI6jtRZwvJQ3CvuCr/6Hh9O8wvnqIm8
MYgIsYFIuoJ9txDgcsiixcJOXM9giSapyzXIRKkS6RRWF/NJ0umUFwGQBNeP6qDo
a/dlJR7LJTKcZaDvRZBpYRa/1zWLFeSNCuBnPvAaQ1YgB1S61zAUB5VGwxzkBFRh
5bTAdNWkf33Dejk3FQEZOGEzctkwIO85DA8yEPfbv9Quy/hBWuYST1C/dbNOack0
59tINSgGVjVkIz6va0OPwm4JLUlePG8O91H254+HaeJOEITYzGpSd8TQZ7H2U73A
8IdIHT8mUlPNcrkMNTqIz9a4KH+D9fvbY1eE3PMs9xP8NeBjj4zqLf7CukynmOVY
VnHx+njMr8VWLtNeBbwrx5OeguBF+5lqHp+FbNPrePmEkhRYhO7PfE3If7A+PKlc
+1Ei1WG7fUtiuW2mA2uWWRFhotZOYnKBKCJ9FtHrTwLaOHFhIywyj9OUNhGtVf6D
DxVmrBpZ9aQkvwOpoiLgzhhYOGTg02MjadfN6M2nilyVQ51UrrOPJhSlmgGArjPL
YPS6ddnAjSY/07hjKXgw/OwFjfkzybFRkjy31b0ffk+LOjioJSDdYG+eiY4ASgpV
l3tqajikHseQgxYVjYneplXASWLypvbb3Q18+gSzXkJDLxRbSm1/tb9JTbhiP4W5
JegsE9O/zqYOBjpyTxnZesuQqkI9aYILFpkFrOD2NF9qjSBLIqy+k4GrUfqrMsce
Umg27cITWUGh92M3hx6oN9HmPaHYNTfXBzPrTNNWmGtni+Vv0R+qB2BWtCbBNZuL
AGEft0ii7zs+CuQdKgRpEFa6xSAUBLBSf4GHOXS39ecZuJWXAskdJv3JNTZGMRxt
dgnYfVpnbhqbZm79bxP6oA+s/ky/XvrJGeEHhuvjlTcJGI8o9K2np6fI+R4IZ3+E
hL2yrLg0SN7y8wGBGXmtBaXxFqFocW+gQxMn97qFLiEen0uZCzNQP0lN7S7SLsA7
PQk9jWA7DEEGQD5Ur1euvCquSoClEckU4SiF5OWGqdCH1X7XRmzOljuz75I8qz8C
GKa1kQL08DaaPGN8hslklHOML09jz7/Bi27XIvjKSiPMaE3YfR9OFygUpvkW8S4l
zIUdXf+mA58QQ15g5ifHJqnYYi1SK4ZAE75yJLJVSDFsiTrABQWVKNQrRFdbcyfG
fR1fmpgvDWxznulk0b+rVvz3wyvh8znlarPlJI9/sVjchbIl0soTuYTm9vY3DaPN
Mdf7S82jd8QUfc9noQ4hNTDGCnCB/2Bp5IfyXVDpIhlgm3sbkPKi5vJ5bKW4f45v
auevjTrGmkwlNIivz6RRQL2H+W97CrH4z7998C7R3aidkmK5yYxJuHeJO4KSuKdg
cvTev2H5RKA3fJMqbBXvg6MVXEe2Zhyx0UA6e5qfXMgYUqjcDjfNV1ifsDtrgJPe
6amENLDh4NQZkHk3VFRyJbtiPF9G86b7LizrYxccVR0OAwwbHHX7OCW181ANWOMJ
b5hywhPbP/S4CLLtKXfdUuM9MuCoLbXpOqwr2qe2aq2tjsLKhlpxYWP5fIcJCP0j
klLWQLgC6UgePSlVdo5V8sotQDvGYFzqQAnrFydWvDxL99kJzSjzosYF/0BUrxjf
78mElfeoA4kencsT2XenmXGgPP1H59JxhzwLMWlug8SDRBj/MOF1TO6GD5TYdf8+
0qLgbXkhg5YD6Ef+OMylY3aDtPm7VzIcSnlNn1EqaS9BmqrbbQpDnM7oOx9PWPb1
0UoutZZPGA0+QhsliKzWk4sToCfikgmRxx5H+JzALECLtgo0s5m9sZFxK/Ta4FZq
VIPAyR8m59s/peRNNTUQaFbuv1k/PiwPEJWwxIz/C9Rn1AbBFeYe5MDZN3MvWoo9
2TS7NJwQrtz3iZExJXAWTLWLMGpvGQNRlezIFHsuYZn8zWQtqdPeF2UdmK0aoCGa
RhU5OHFVUpS2KZeD49ubIXfpIC6GMeu0tkCS9yQAJyqZBJ9BmZdrOQvBn6S1bKN4
kQFx8ge9Q/doVmxhrIyUl6KbxGIgZ/gFZ+sTniBVDQU8m4RAaZrFuqU6P865cYZp
rZDLfjV2SuWkH37st9GFmB8HG/+ZTqIG9Ov6tSl/Dz2N9UVYayat2A8lRck7RjDG
XA44efJpdNPx4ErPXMXscPBuZkTh4qvpdStyjCrp+YYlULKmPppJQm0gfoCUm0CW
1VpJ3oUN498wBgMb5xvwPD9YISP/oDUi6YM5wgOb/KTvuaSCOJueUiEsI3QQ7dmL
ePjZKyeSi+XFdLMhtMistPhYATqFk4XGPCM2tfZTwXil96RrYC/BEh67CN0yRDBf
OBJrx1Wd+NSW7oIH8lc8lEr4G8keQaq/7LnTzmsOPaulIlpHs2/SypYaQmdBKsFb
ggyRCHCVd+R8V7lWGUjJduXEWLGvQQD3csbGSM1t1XWcbIB643csKy+HuASo9/F4
llJ5hwyQ017tLApIs+tZ+mKhVcb2uTrNy9UICWw0x6meA8CVcaj7Ax6tIklmaBjh
7bl6d38/S0faxp5cQLOLtlBLQ49KZCCYhjxNxY0LwQrdufZJgh9tkjgaxM5pKuQb
1S59r/WWVF2iRlNANqbpznilOwsvxe/HHA1EdC0jz//tGImjERKUHAKVtI+SvmQQ
oqtDDoEBK7eMnHxLt7R5HYIRHJpSqXOyBxbx/5AIVGdqypetvjAif/o9n1v8+HkI
B/g48N7QPKMut3/0/FHsKxpD070MhOFJ8kUGJEzOnFft/Nwva630vTZIjTRpNbeL
bUyLHs+WBLzRdmBkxUfyCke0rMNYuGR9DqV97DibIE5QukXcCzXu6uxVAL4Vzmu3
5nWNInmvi5d9KKcjyD1x23UmYbM989+H2nqG9yxqlpgDwrc19Zv603SjB8xoQ/78
5dbUVdL4X8FLfaUwUIP5vVvqRjyZ77v/0O78QlmFcI11rLaG6zRhY5kgDSxItLEa
zGckW43gYK66qofIDoYFlqOdEnmvsEGJWkuLlh5fcvRZ6PZhIIu9qEVwPRNai703
4oJpeYoT4+oYU+90Ji/gjMtesI9fCfw/Ga4wbxO+712mt4E2XxZ7JcWDvCpAU7lV
hanKKSZU+61ltukcA7l7G+Dntrc8TBtm4loliAxJ9RCKVwf2VjTrSzfDOTDW3EeI
TE4NozbyV2xlAkl8IBhvimVO+yGjZTiMC1S+urtklyGUB7qMaJH1YI38vr9TXHn/
83F4/nqDEMFWHKfa0bPEpqTVfMV28tt2tDE8c0iNNMI4EDvBKB6dGsqvb/FQwRjr
+5qcPmPQPTMWzoMcIGqsIWmiRt7hZpiHION7+HfjdIuu9PVVUbhMsxgt8Eff+7je
Fil5K65Xi0qIzIvmZSJ73cdKc/llnl+Se3x68FjCDgK+GKOrNzSjrgAhEq7j6Anc
86nObnfX/P9sl/+QX0VcwXFM9mkoxeTmvnYYucddr1ECfIFExhLOgYfs4jggxlOW
iu9wmYPshLfA8By4/GtVheP3iG1Z+ED/8S7RdZHY75GDbHM1HwswwEUjh3qHpINi
kgGz+CWxQOnrFEu+dNY6gZCu3kkmHHLzIUUBPa4nem8agrLxkz2WmQFaCQO89aX5
rMS/h4GodMiCXB2NHpsZl7sab/myxbJfPI2VqgEvCfCAwX1wTIIe3qGUiOtVJOh8
oeHacavgFN2NmRu1sgzoqwB/qd9lCX6yuqRxeFwko4ZRMSeMW+EJTTGHbw3RjBFU
0pl85YX2YOQtASErWhgAV8S4os+wkI8pIgTlJYRaNBZVENXzKfiD0bhfj1EBjvy0
XNtJE1ybHi1yxTBPxyKfg/W5YiGDzE5TmdVN1oLxDKP5eyfZsolOIRsgGb5n9O3S
ymH4+TbgZnQVTLotxcUMAhL9m7ZEgkE/Vfv+JpYMC04zBx29a8g+OGCtTVhjJMVB
C/WlOlrL7bUEV6PwCNaJp9mJhJ2LtWYYIxLMfcNDZtCECyawpwgXXnLdCGbb4V2H
W3IY5pczcn6tjdmgf2bFJOEIvN55P70NaznVr8bgpIBI33svJCa39MopmJ6nhrLQ
X2wFbUtmbQWxyD2AoOhzKHcL306863Mbz93V4LXVYwgZKI+KeRtFz+PicLml0ATI
FUTKRhOwh/zmspZMGwZexFADd8ZIQ56K1pvHa2YQMl2aqWVDG+W4GHU8Ws2dziTy
ri5nTlWZr8/nn/Ql66mzqg0GbnnmqJopkgquY+nm042NX9/BC8H3hczwMOGy355S
onJ3N3h+eQoZIvz9Z+IF/MLR/dYPnxAFZfnQ4d5I+qpfmNo7ybLgq3G508xR0tFk
+tb/WLFxCQiHnMqusK4yKm38q/EMRAN48OUadliwMmtFtT79QtYeB4vG1QTiHUtr
Plk74XfIO4Q2RT5DjWaf/3UX7eIWCA8dS9mYkr12bW+U5leaGsVnvTYO6jXKP8EV
i6GO+RpQCCjEVPPISqiiqsoBgxLQcXOfDIQzcevw9vwSsLlmB99+pajHn3E8hP5S
uk+KdDGVYlUEZEMj0R8gTAMt1wpicuZoEQTbmt27ceL+8izLUxFtjNGXVtw7Vr7F
PkzEqBKz8y++jbGFMt3tEXUP22016elbROGrWe7L9p75pbvHvrj6v37H3mn20p2d
nZ3MTJFxE+kbsOnN2WGUXDUtzWi2RmYvjfpshXDcXLPFb+DZYLkdu6SWJ+vq7B/B
5lOGkp+GVp9ELvyEtGWlMh5PaD20eaV/mmRxcD4DV/z0SUav7nHw6PT9TZ78Uml4
dh/0579HZpCZvLPbWc3o7FaW1t/Uih/9EozwoffoFBqdv4ipIZlLQMSDT9vcWy3G
urzqFea5FCSTpJjsmKzQU//dTEagk+yUeG5zNrKJY/0hTbrgMeUku2TKCJETzMxm
/JTsB2gocs7Xq2qO0ul0TGrydNnPR3BzHDVM1pj1MnRV3LL1DJiLeixHa8JGlBK3
PXIPGOj8MpJnVfXkG7UO99nyy/Xqwo8JFjVhzp9h+S5WUVMapMb0sgBOznmGLVQD
fFEKOkddve1AWrmGC4B69cJ2cdO5QMZKiTvNMTS77/hlmb7Inj9OGDCjtbGglsiB
jssCtwdR2dR1UDKuTiCkI0Yf0+UOya6jl4wE0FArYBv+XBmqQkeqeXhUPQVLVQJG
Te0k4xbT7MBO3UvsykfeWLgzRJ1gt/Tc4+3wCuhUPbwy5OZcAsSadvQXWph32puj
nuxU1pEsfjCOZkkTKBgM/UjMIXHrULyeznzKuRXM/5YT7rJRH9R8zC6u6eA57r+p
sErOLUnt8HshTD9i1VsiK33BNnmzZCVNvbrtTZIef8gkaQsrq7RBrNbvDlssmpEM
c93e3MeaBYnnxexlRl0bVbi6O2Ol9elz1vuBK144KvRonb63WPy53pps7dlpAA+H
t024vYJAez0tcdcxeInYfm7iFPHY/tEzMY+aJMyJghrK7CVrcuwhbEj6WdQHME7J
jMOKy7/JSfr91996ijYBkJrwVITQOfFsaGKf4BcLe1r+zYpBpozahhRTHHX86ZeB
KO4zLFbyHakHTl4j5Q+IyYMhyUa1opRmkFglBbgfcVA/798/OBVu36sK5HgMM3JQ
bKAHo7V9oNCJgsG992Jh/mNgdGnYflvpgwgFtmOOSYgMHwGj3VQGocriLA2F8WqG
mGjOT8SJtf3miNaAkAh7ISPa9WnwN7XDQY5Fu2w/LbUSj66P+DAYCr8yBdMolQNp
NDnKOR/Gib4I5o88nThDui84z0Ur14hxF7BhZVC7OnDnQqOQ4BOvbYf04bBCUSj7
FQNswofo5DHpGWLB0Jed/ymRiW6QRl3sG+C/Up07OXUTtXhuAyeZvZAdq/GB7slj
StZ6PA/IHrJ9oZxQeZ6kCSnmb9ScfirXoI00SsNhJ8xA1J/YemQIpi4MBiwSYqIa
W6ziJcUbOXXVjOYP9zopnGfBFha4H0t/lUIpanjKkXXhEhefL7ygAYu9a0ZRz0qV
YBr1q2o7TDLazNy405U0gMQBR5BHQZsGLOa7MOIFher89OL+ljJk+2EhLogj0NsZ
u5B0koQw5b9srlDPZLS0b1p/ESiU2afQaEvrR5TKuxDUL1qU0p/snzD62wldLaQi
Wqhdw0VTznyb/DlHWX+TIFugi92+jEROF5vQYXJ1vHNjDG+r3VQ2R2o+djeT2SmV
flo955UX0T6CHxU7FRaH6i3pdk7qQuhUOLptnEbkVcxAnhII2/pDnmXePlFWgfhK
qHtLcPNMe+ih/u6bVF5t/h/btEKATWzlnWqhqRQc9RApJ2wZ06fMWosQpDoteb6S
EH3uv6Lms2uru5eyT8LwygVOm99CA0AKkN4ARHz3NI+Qagta8KogH+CksDzamlT5
SYqBUC45judxfBN1ImZrCh3vF+BGQ04iuHNeOGKH/COLJDEntFlmSdvA6xDZh/wF
yprn0R9gU/08J1FY4JSClRh7FlCFw7sYr6zpWQsFB7Cxtpx4zgb1aNW59MpHIATv
6lfF1z82lV8vOjjBKSPcD7tFlAN4ulscp12SbThTHN2yCO/68Tf1axDR3j3ngV6w
u+w//vjzE1tOTWWbepYBzH4QQrAScqfk55H3tffMDmAidcBmfoyRGjiQPGUKgXhG
lNuMvaIh9bBkqKuy1GhSYpikuk0la4CKiNVaBIote4QdRkqprSTiRcRXH/aWstpa
rrrxERus7CXcFrTq4Is8wpfaFNv9YIRoypBMcIA34jRj4Bd6HUoCOLdIQ6CcPoYI
v6P58q9Lfi2ql4FnxBy6u90B4SGe5SiuSnT5k3qw81DAenuESjSvFy6EbKnx8LSL
O+DTxUb8z1x5ZmcP4qXPxCkt0u2Opy4urU5+goBhkMaxBP9dxQJbGyCc3Jk+xOeW
3jqXHavWaieP38TyURYe3MdzgqWbeugIsNB8aDtafgn7YAzOGty76YxdhD4AUAm9
5u7+RyQNse6QsRjY0UP5h+lkQnMU6rx1IN4heU7Bv077/+uSZnZYntNHpekdTUes
4cKospSuiHjFvpPv/7lR3DrIbd342yPdapW+PnhgZwTJ4TcMjpuvqkpmPRBKkBXk
BNSrPLU5L132ekHEtog93/DgvtWLONMjEiOw8HVQHbHvkY8EDSVQ/7nWxu0GmJhZ
8SZCjR5vtHBk50xyf9mD21/reVxhrbOkCQ4V5V2uT2Z5+CxEl5gKblV5sEIJIv8S
enmDALk9eQnlz5i8jdT2hvGDs0bgkT9LmQuFqb2wcVySoO9FWloQVtdT5GNTWjVH
2k9ZCCPLZiR0h6LjQ/Vk2EYa/MTHst5VQRiuFsqbrRJeFsWnSuZWc2AKQl+qTEK5
k07T9nMlSGQ8O0MLD5dmBrjwiBV260Riob1vOmUSl8yLOUwF/VHpRMGxaqbOH6Bl
eO1qILlrD/cEsaFP9adm77NctTENWj920TywVwO57260GFJlybGM5vkAzXnuxkMM
O9+539ik7HDX3ypC8ZM3A2whQcsXNRV8GoVhV/vsyQGZ5UjGIL4Ns1hws+Iuevy6
0DCvRnOFcbuccl4JiJVoOSrtNMiLrpqH56aCf3pXv7nlFN5w9Sa2u9idmb3WBrIB
dUjvPpH7XJ3Z1N4V1zUt07twmm5BI8AF17UVI8h9dpqw2uuqB/6JM5ejplWa2X5P
K1rsk82nvB0PD8EFr6346WnhcBDVufObpO30JhvsUjr+Ls7Fuoo/dlmZkMC/AnZQ
qAABF3JasR+Sb1Xc5l48vrK5jNzKtXQu5wg/5UtZxOGXiVLwcf3vRuZx6XzEMFcA
AFtqaiKU/0B378SVuw7HR40NDxvFAcIGSJaHGk/vOaSXkqlJNkpI5rWPnU+fUi/C
24p9DZSjsz6+d5HwoBS7pvf7NT6W8G3t4Bcya8SVrPsiNonpwOX7EQP3iAsixRK4
q8Y0ssBrebpEVU6sLwz4IA6nUDtebTgzT0RQu3MfGGXSbjy0GL4WK1SCQIQZnxGA
qVvxNC8mCmWJdHDtsAZXMnuJkMEdctgWNSA4Li9sUMqapgLoKjaxMpGU01eMEAyu
d3DKTfRKs4+1RfJg2gsOyiGaDuWSqB9hZdCdqmnGOt55qRh9GQDPYjwHa9G555YH
AIzV3J7YbmKxw7DTtz5ui/zkHn8eRLXRtWTGGwIIqGpACXpgyBpOrM7u0OTICwqF
RryqGT8if+dbH7r5jLEFtL20vxcP8MfP9F2XBjgBbuConBWK+/SVHk0ebFLtIf0j
MIHPw/I7HEx55GOsUwqygkkUPQ0tiZqmwJSlLUcrlraxhOyjGtblXOj+GqcSkXiJ
Kz8uPhuo9fft3Fb6NxxcWs+zTRIxgXr4PiF5KI2amkFO1JnTSZxTGP8TIpQL/5sd
SDaEmbDKQdg1AYJgjx4+wPY0wCiyd4G2xOMn4zsjZwG3xBOexWmiC53Tyy3k0hVG
u0VpjMNkcTIWdfxoTcNWK2pHZ119F+EiC+HE+v1niVEhSH4A2Xn1RX8gt020Hg/6
PNCucz0ehvXslAy3yQSR4KWHqC9hIAW8ESS6wwtogxzhNRLFUHSxIFV2A1YvRcU6
WrQjdoKDDR3SrGfGo90ImRgY+CCVPn++39777JIcfwK3qUtWGqR0IHass6eb3Sb4
PwvmdMEyEu49dgMkjHAExE8sHKs0LRVHploMf7q879IsxBLtNiyBr7A65chYpvzO
4QEd1R0nIBX6lGCLqOynNdJOK24CxSTfRIp8H54Ln/63F/ZjqCee/Qu2Ugk+x+/A
s0j2nEgW/7enavT2aKavmw+yKfTNltbXENbOzF24hTQavwEfsohJUa2qh9rllSnd
6RJ2KCM6INgE6hy7BlvFh5N3BKCfDEfb/qqAah+FhFhtlh1DkkR9Wb7ojM979vmv
UClr2mQQDmrM6b/Uu1H+Bryi6/qsMHJJt959lR+tsGM0FJwBEQFvt9jbmlyEcJad
beR3XoV5jyttzakpx5lP9/4ch7ohhKBn1Kf5QuvO+rxyCBroAzw6UHRLms2TgMbh
LZQqH3C8t42pC8T1OZyD8xls87vouxeXTTYA1+yBp+FtwE3YzgNNLo9r6IfTwhRU
FzTxsVEGyd7WBUi1aHZmCr4bn5dodmkeqFnEDwOs84927o68kaMcVZvd4xN6re9C
pv4avN7sguod8qe29ZuEQtCI9aHqm2sJJ16nW121Cn4MIOSWG/UQV2Cf/OtWkTL0
bV59LexxjfcswugS5B6Ub9dNeyoS+SWrCqfiCsPTyxoprMSI4jX1m58sd42P5WAX
HseY+oVQ4Fbi0f6DMSenjd3RgVQYCKyaO4I0ecJ2mYC5bZEEGWMgtBPsGslOLDGj
PrEeWWNL552LNOFO9kNu8Il9sxmaTwuQucVRN4CFCLBdtSyPptou12Y0cHl2epr2
/2rtvF80jdn1p9NAzWRbWjG8+GHcn4Qpw+URXxGZl/E1WR29taUaAabkmIiEus0z
NQLBdW0vf/0jzHwCkuiSvhuzwIgDLM80SxJkY5V4Hz1toV5RTB7dybaje2w4N8uH
4JmlYEut93c957tbHq8b4KwZaLkgU8wpPMXpTCesyf8ySwqqcw8cZ7gBaH+ws5L4
oWkNKAfHC+ODCofCgss0yWBH+pbMzFASSKZhnjtHkN1OD4+P3Hc1PumQjgwOZ5w4
jnLXBcS7hPUzyezhIjg6EhV4e3EmoLsrowsL7mMVIosCIyyzTMEmvENpq86MfDP9
0lV1eyoAcnXltrujk0xNtO5fMhQFFNLicGlmWRx5IkQ5ZYIT7kSXrLZcMy4a1xwJ
dtHuF7z1MLT9Kot/v/BWbSURzb90GyHGYeKayLPMETPj39cs7Rfel+I6E5L0oj4R
qvzsYYwfMv5dNCRC0rwjFmE79j8yTeztWoYdPKIGRIzbm2CuMzWNb7/GQ5pLLkGl
XfzCNdj6GNtnd8KbqKzrmWVSKKb/i/eBI9luhOKkwmrdKushWxqwtxNg04pMzumR
+RM0GnyIqAHf/PhQkkGrzo09sHuGOeFFI3gMFPDH/NxDqiswKyvYaEyW8uoXc3vs
ANdn5+Tprn2N6PjFkuQXG36MB/7SjBtNg9q2Per/VxwUjLuh1ZDugYCTFG0XjlPm
iFgR5yjQYEHRQHFjOQ7EK70WnTHw/a5oX1qBy/I//eNYuv50QWhq1oxYgJ1lP+so
MnMUyT95vPYgNC4gukYToU8fo1dxyHgbLAJj/BnO74RVn0psA5ueVAHMg3t3/Yrt
ChQoIxF+cD6lGOUSBkXiLgVLjPG/1J0Tz9WqIa9ygl7hOE8iZ3iZfmDvohNTP+Nf
jysl5NsGMCWoTmY8BtyfUG4U7Re5Lr2sVevHDzBKZsAio7fXqpY1QjN4o+wUdx2x
ZdyHEF6FGWBtX6WM6tABnm2v04WHEDPRjuBTgINVijRvLZsK7sa8jF3YOBUN1yrE
hVDYWqsOhxn/T0RExMlm/QUqTvcON/yL4iSiWrGDdQFtKmjzuZ83Iq/AoICGUTiJ
Gb6CNlNeeI+fke59Dc9imW21ENEl3nzTpKBMWBoqPKZyMR/4EGL6vLnjliWROvfB
cDZI1C2qwKXgC5C8PA/RZ7y6ecVykXFBttYoUUh7PUn4i4PT9WvikOFQxdCpbc7H
EPFy+GED5bRhPIcDfXmQ7OjSySEcPKa8uRauarnu/xQPVBKKSp64ZfKCHwfv7SUG
Whqm9g8NINaNt6a00uNoxPDxN05JXqeqaJbxV+AbKoe+nLcB/A/mHLJOfFGqNm8o
m4Tds+Un81CJIZh+PI6Qd8AZfW6WadFYI5beA42z9oZMnGp/BmjOSesAhfCPjL+W
9nw9Gu1NTufYtFRZN267VpZ+VsSlut8wpLEa6uAB5SdRFNUBUswd0URR35mhDxVw
V963EFSHj3CHfTxgl7Mnmw==
`protect END_PROTECTED
