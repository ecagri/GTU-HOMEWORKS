`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hsk//pmNecpGyzr0+P2/dVCgf+JD3v1gIVRyk75UYYJ1R+9+pTBFoDlm+1cz9vrn
jZC64dmmpah8Vcdo09nT+zMaPSICT/W+0ewrsYVal9Na7rqxX87uuTT/dNrYHDj3
lFPglXbk8zSPCdPWYneRGmx2+2fstuhf/kQXLRfL7NOV1/swQ7AMv3NVvfAMmgec
xskH4oYfTR88w3wpyx0+pdVHy+QUcLUprqR7lGNWhQMT7R13TJKMCrKB7piQVofo
AFZdCp82mmFzeE6bvy38b/aJWY+pqweSGEZHGIvHKss/nAODujf2z9RCRt7zJbsU
LDXRdOv9mjYwPrx24REBgHoNJNGqOc81VCWQOdarU3uWZxxAW47GRTx1K+JkaQY5
gXpl3rnJ/FHAn336WsRg4gt6Fj5OxTwxvtdhm0I9giO05cqJJbgsud8CSyvkSka+
E8D4y40XXe8rHcRVGMzegoidpSCYnuD2RwSD/jhmptheTFzi+GFvxL8V0bfwAUHC
2Af813zUwv6T4GHA9mZp38RzYG0bYHwsyp89Gt2Q5QXcv3aKycll4/eRIIKarAB2
V5w8FEupwRSTOfOTxUAd/9kByoEtpCeZ9vNUDhuZz3sfDOGT9JLO8ssTTKVmV55P
23iGR/dJeRLBhfozfM+Hz/u4dDwDGdpN1VeK7W7i0qiA2BLyj9wvB8PgciCnYVYN
7byXx1M+eRb5b6+kwjY7BdtQA7uNXo75eVt4PyxBnpmevgD1OzomsTp3Z7MANQjS
4NMwm5eK4f0L7J/UjjYMqCWDyIJsssOrgup4sIbFeq587Bxmb6gFsQcm98eSqr+L
AAdIxWJ6dqR5zUiJUgqWtoMPLgVwSCwuU+P/d+lleK65C31IeoLmU9qImQPQYM25
isq9UTPih1TheDWieyPSdD3MAy8u199FixmiL5YAh/YtpA0NnAhB5x+1VPzbkYIa
RzgVICzkAsgCd/5AfIHyaRZ1ihNnJGYJweHK+YpUyjBX+hq8+yRotjAZpByAKEaQ
pFL5m2Fi8AQqlOSGRcmKDET3+OpP5Vb6etaVpy6I4Enjs3J3oeM/geLAXB9dJ/th
zCP84eamd6dBvilfR+rZEAUImK1xlQX96YCQV8meO01PvZ/0J+hdwnnJEHK+Uscu
Xg6MWfUoZXy508aSIiZ2nHZDbFY508sZR18eXc4i5vgKuGLolybFnqaUiYghEsG5
agTP9nqoEInyR4q3COpUsMuXrboSZsfsnZ4JTIMrNhXBb1P0ttp2JVqkgxtFDm8Y
H/TFgiM20hugJiyxmfB31ilzYhwvDFO7ccWa89ehGM4/hA4e1WLfF2bTq80Pj/MD
9ORd0RejXCJnaFCnahWsXOcOr5O7f0OUH2XYlmlALhEtf8dYqAa+c6yqFoariNE9
zSPmCQvG1I29X15pKZrT5vLRnLdhpvRfxgrHsruSx14nrC+vyTe24Fv06pZNFbiS
ZbVVt05YTvOnS11IxpB80SnF8kL79aUBUyoof1PtQ1U0cf9YCtgsCBGnSyCQ/S/3
8F0vEWb+uulQ0igxPIcoPg3UR4uhtdVthsfpBcyNuEYw98fgRorJRYYe/WJlq/s8
1PGFzFWct4Va8kxyMf4YqP3UH0BQsOdy3jkl4nW+CXH6p+LCHQi0pW/pWvH2Q0EV
E+Gxv3XmEEvWRwdV3n65EGrpNM+gUaRFpPbpJeK/EvSDhptqiFh5C10T4Ve2a0a3
sFgUI/iKcSS2o/9ZM7akuyw/M28Vg1sH+IZAq71yQosYiTvvZjK9fpfcR2QE7AW6
eTOOFH7FooQ4WXog1fECE7V37vECMqQa7UMX3Z+6VSvcrMyGWIWAyyIu8cabOeGF
+MrQ6xf113ZCSuUk+4Pl64wgHHn1zue/huKEWR99JKRS+6PD/N42qHwveo5dCE2r
Zib1lGE0WTeghL3RFhe+Wo02o9K2AKCemMeucFPkyR4TdbbJncY/tESednnveNBy
5K+pkHV6KsZMVk4PMg68oiWgTRG6+UnyWL1KmMqHot/j6m9Zg4/NgGncf1m5+26+
NVKfcqIPzQTHGigT07cz9kaK9FA2+z+9LQczPlhGgXZv3xOmb+YJv34yHkpDpzBL
twShzkwpEHVrzm0NpAdnEqg2lqy1aYu/6kgjy3uL7pWjMUJBNH5yCdDxk693MM1y
Jdv437EJ7wjXgU/yRsAOdM+k/R/SIG1iZ1oHMyvzJfdf56I4doDwJ4+9v02DoPv2
pvT0xQo2r/+XGE+/Ftts9AyB91IRJn57oC388h194wBCkdxstiefMLm3Qv4LS8HT
33gidmNV2lDrWGjIVZkKttvE+gU9zIli9oNqS+UJmsASrXWbJzzEuiRacgV21BNr
kW7hJfo+zwddBc7Iu6zdw+H8ZSigkr+/mEx8aifLcMmrkWkVqhFUDGVwXp1QRIZw
ItgAbbtf3Vjj4Ykyr6uj8xVUi+88LrNFGnnCiDMwfKuGohfO0SZeDmgpeTCg4QTD
YWuwNsJz00MZgAZg9ivam4ACS06JTajmKkYvLfV4x4cKupj+5elGxhcLfytlSOQM
PNCgxOYjnCr6h/YysO5fF3H9hpUvoVDVK1M+ZXNMhvomjw/nYHU4VSi/QePDXYDb
RAubZt/KKRavVJqcKks4XWA7Lc53O2l0kNcABPaOQqJOsHS1A4SoHzkVYRCFlWcK
ZeCDyVHRiuTatWU/JooQsIwgg/SvhIOwUv1eJdyiFgG6vn61XhgPew1qnK7WZ+44
080CCts2XD4oBLvDAkdvVUtCTLx7T6dtJCNljbj8UUQTrLRQAMGPpuHA75iAks0p
TsfLIvD79saW/IyTG/RxyETiDgAxwd1FUHuzPyUobt4H1agbtuJL0m+mnp/EbTM+
6xXAzZKevoBROL45dKWG/yIXKAr8EiavsNoJHVrP2m9HnwgrdOhjcrVv/uxIp88+
y54YNrLb8cHNYsowgkHMbFV7cU+4yXM6PuxG+wQeAI8Wms7Yb4qn8lZOriKJASpK
+Y6s6iZov5jcKvKckNqPqbd13m4IC1ILH8eRDNJpF3jOcsWvCD0/EO8hK+o9dH3m
FCzA9BXLLh4Ka0ScDoDrM/HlZjwwx6yoPCHcN8oG8hwBsoYGVwmoH7ADQULc5zb/
79rmx5HmWOleGdJmFzTfN6N9W8h5Pk2ntxkHsLPqyPzcPENodefEz0O8IvGT9gO+
qIboSjqJzB78vJoJ67FeM6uDu8ciE9yollaPq+mnS9y3rc5Vw1k8YBKnLKJAj4xe
8VK9/Na82REFyIDt6nS4pwh5WhisVnXWtlROGPzqc0uXyVc/lBXdGLGVhGsVv4FD
a+IuIMIasmnGbWdb5MMuEgywO6/VYeYhxK9cgBYpDtqso5GlTqx6prdPgea85BNn
0fqcudU123t6TURgQI36SW5VSfIO/BaWN86/Cb0wqOzlA75ocy25iiNEZkgZhWSq
m06of3ko+4UB8CYwtFhjtHB863WMdb2JyCIZNnRc34wKu0Wc+FK9+t5kDAiEvG/z
4Q9JDAmTPMgdb/KvJDNH4zlHw5KIg2WNCg+SSo7z8PqN5yh+D4zKlCA9ZBoIx2dW
giiClPwUAR4EzZI+viJeCPWBGEqnTcpEwt0odrLtihbRZannBtpEYoAmqybTIiSr
yDR+x8VW8CUfqZ1NRjZe37FwuCKkzHsHfQJg6RiyB1rvc5kNJRY/EmASOthNU3Ud
Hvtmmh3ENhFdPBQtJevjfUwA8+KHPJef7Wl8Lv7mGm/Q+bTPdJDobuJLs0btzhf/
auFDe7WdRhHR+frVOvtswiCkSYo2d0LLGEWmeaUddqyeplSQNtmhl8RLwRFQqt9V
JXZXlZ9npF8BjVG5ULtH/DqtRA9dyuqp2ivC7cCPLz/VEDZIn/AA1+tly769mFhd
Vhu7To4A/5WTLaCgar2xyrVNG+4NXzRB3U2GgNzQkSpGmvJaaYpTKjS3yNfLxIoA
KW7XL//bjlPyVZnTFjneoB6C9rEmJdK5VWjYBxnsDBY45lLd4wToOV59ZodM7NJ5
VB7F1VmAMjGMXgi/gBwncZcQsAU+qE7thiAjk5WPeFY7yvj5g4Q5muohhYoxhPBt
iO51qFmv+d86YtTkOs1IbF75HkyM3dJvtr81cDUgGKcR2zTT8UCA82jicePSWbM/
YR1ETAvhE7lQm7oPWELRI5+y5IAl9vfr0vFtDlAD26DkYV5DXjnWtutjZmxpJNe6
8pqj0XTa/kwHCG/MvIWixnhQ0UwggYOLMTF3F9iZh8Mxawc61eXPVVA7tHnh9r8Q
NBEdUT9O3XaYlsL8Wupyk58osB40tSAyMLt5zzzLxvjjvFBSOLjSzYbUimAzg4cE
2XmhmmSAtb/Bz3/Vi+zXrEO9NXp/b+AfwpMIAIDqdVxYXst3KybBmoUAes04aI6e
YFW0aqCjS/PEZ90FELqE8qxNJqtDTjt8R7+ZnWZbAqih7/FVEgDBRSBdVOa60vGN
5CGBElU6IKRXxEra4Vo3zJ+RJONOe9rMXWGiCz2dvpcR8uUDobtS6cNm0DPGl/U1
vlbT67UcMUMAzW+HMyrdpYHvQgg19nJ+mStkyZUlEyXljI5DGRNcnAQ5h56aFnoi
3QE3UpNhC84/X5k6v8/FEz9eSCDPlSNTUskoiMEcLp4IwnMd1zQelX2J/ml6c6iD
IB1QBEJS803r5gAm5daq2QIqa6AH787Yfmok8ILmFbehosW8y6BQuwpA4Xu1ZOEZ
w/COBES2uADySjlo9LXSrs6ZMXr7R1Z8fWJ3gv9d5PZSFspd1N2avObtWzFvAdv4
Mb9mDnnjKYVTzTzu+Vl0aANYhfFYpS+YO4llJk0RV3NZJRuXyv3iylQcUiVA5vNf
3EdqKryVKJ8ZVzkhLkb+S+KU1UVcKrAgJdbtH2Ych3Tybxd8yV1M97EcUrXSYsLI
ad790SISdKIlRrODxaMOMY1Mtipz35oBylqrwPkHhSGKSKTO9aWZ1powTxdDVLtJ
sRMDrTyzpzzbbnMBtxt9uc9AExHwWbEOk9zzuRefNv1tqomNtPkl2cJ4CnmTXQSv
6d61yqvBYNUUV/OoDli9ZNjgNudYS9NuVRpz1+GW3aUKdfesLI+DEzMd8gy5ZI5r
B2skbLfAyEO7GX1TnJA7CXc6nVVxFoTI8aeQCxA/+aJuo7KUhoHfSgw4JWphaRUP
h6itgd2HvgjwtlESYaXKT338ZvevNgksEZ0PfU51fLGUFcqLGM+l9w9OzAzzOokE
+h4eycUzbZpRtcpLzBzMU5apZvtL/MJyMMDkwgKMmskIJRsZ2kepaSrF8Bn2tE9b
eMbbpdMWdHMl4IZDl0GbVqDbKXl5K3Gu9aJ1L4WivkoZevoGSkjWgBNFYcNFcBxk
N4s8QU9ywzcOGOY5CfZJ5y0tq75okdlH1XpvFyk+IGRVWPVFh3JZ0MAs7QmqDYYO
iEX3uFJEL9YGJw1lpb5f5cNmRPlRISkDeJqMwc73qr4dI8rtysFsQ+eSpd9mRGd0
KCnEd3n6GySkW4U9ABYMBV8Y1zGi2GEPA8h65J/uPtc=
`protect END_PROTECTED
