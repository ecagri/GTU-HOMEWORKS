`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9lzDjO4T0hyWrmB6qzkvuUWBdZhYu6UO7bIu9Rbhr9nwTkyibh0aTYsFvoxcmAoC
mdYUkjTK9a6Vn9G6aeTy8hgAwe+Wm6ZqS6Ox3+0AxcuN0lxYqx2IvzQkRhHhb1+I
+GKSryJBwTxmN/YH0Q6oujvWgeTod35LZxZPLNrp9rDkzaYKHcjR78+6tSxgv+Wl
1Xuxdoew087BADM8p369Ivv6g+Y3rxoZiyLGtGl7SxLQZtTZfxY2InY2DF6JRT2F
xUPHw1L83gguC1V818+6W8IMymBAHbllLs+H2rfuuKo3J4Jz2XidMKVi1j7JLHow
yizH1C1zZmw+mvSRBAcMRb0FJKT3cWMNMzMU8n0aauWdpbY8VFJGbdpjsZglxwZs
w+VMpIbPX47lTihjTb7dhEgg4WLmsREh4LTIoyHg/6AY9XW11nMaPdVNNYHnkH7G
Ohdlv68wCG1gz9uN4nu8iG4pG03MFgMIyiVj/IbybTxcRscd1bQdmv530YRtDDMJ
ZejgxC5Z7Mn99yz/NY+PiNhduSwrsPjNQG5w7jYofmziRxMWQWHCTmn6v8X5YsbS
V1VFUIXhviMoTHIf9QXpYHxyMmHg+kWyTRqZjZYxzIZAuBDN1gTnl916phQj1R5c
G5+iGzVNL6At/9rtkYPEiAdfQaVnw1q8kchTNX6yNxNly7j2ZuTNKxU2qjGHMM2g
rNB91+od5YJN0LsyQUSpZNasXosjlSm12f44X5sojcXkdoqNUnnYsOS99VZPqq0B
8C/Rsg2A+yGCDR/gcc9vJC091wLyRQYz5V8jZ9eFMqemfFpx1D0Le5adBGXHarFH
6lUt4KWI6mQzPGYF4chnyoJkR7gEM60ePenRr0r50lcm3tHO8rRobLaTIOq4G6m1
eRXmcCJ8Ng+7ypvBCluhTPAtM6nZGuFnqaVS65jv0VL7M507glOD4uY0x43ar2eU
QRwyTCB+NAgJ52+nSYhWXlCheL0T/QSS6d6VVYwM/0AKYWPfeFPEuMEpRQWiRSuE
TYHxRBlo2eihiaZ000mOBJU6iAZsui6fhnqZvVMBvA5baClhu7VxtT81zNvhdLWH
X5rPpdp/o6C214R8ARmbddPF6AcAqXSHxu9G/ts7bF1qkwK7jtCOaE1YCHma/TA2
7p/iBvhFqoHJ4AFSeTL3+MEDhQC5uUkxt050wltBDwzN/ptcO4MklD/AHQoqXj9S
bOOVcxT9obLzetaCH15/PuNPwquJ/rd7B07aqYxTVjg1sIdhsrhoU8cbZ7Us55Ho
BKocBhURw3dLAICbmxNnR5lbByoKqtzxRy2QijCPCAPxkk42tn1q81onlv1IYP+Y
3DVmvfTMw93ipwlfUtVTttdXYKcfU0yl3ZgreSkEbY/MeNcFLR5dyoUYzi+9zuOd
LTRMA3cVe2R+KqmOOZ6jJBfPUxBS0YovJmJN9p+6he0tpVzTlv8rn/++rwZJWJeA
u7Bwg3y0I3jloljSwp8vlgm/jhCHPD5PJs8obBEUKGjjrm2WfCguYeoyz+VdOaHs
pgAQxI0eEtj7Ro0DreBvh+cxh9U4YdgewQ7r3BRF40QdA6FlD5WIUEw1X3hWn1la
XglDTzPF7KSOqiYhN/DNw64ohbpO1J6jvf2Iv6sK4nTFnPhsTcPE3Q1EkGBVWfEx
Dp/jzZoO4X6xsIiAB0wjUvehv9Mm45NxxVPXX/1Cf8fXOay4LYf6Din/UfUg7OrC
GvOewUv/iOAmyTTxVdlP31MhDFPnsCOnmGqgQbWM54P/H4O63jx+dXNCHA+fKsp6
zHztzHLGgYtLB+O/GaoIkg0gSOjH7Ly69OlrDT3QwhdnL/Xd08BOaBthuIUgEbVN
Twuq5IhnNuw+myBHwB8e7BAtyJQCbelMbb87y8EJZbm+1EezrU959xmiJOQjzIUV
wn45dgJSf9mK8L3hv3emHRbZPwY7jIkdfW+SC7+HRxQE0YlWzRSjVL/eaaxHn0sq
V00vgpvNa0rkIPy/KHz2eIH6BnoWLkqiRqy1Neuyv07YeqYTNZlne6u398OC+oij
v7VTo3/oPuJfTzitoSYkqyImkcf0gBc7RmPYvqD2EhZlT4lkOC5T/3p7o5Q85DOv
lBPynWMiWjT4Fl7fBKijn39LbGZ4Op/fRRPFv8njr3+gqp14+iAEbOxAAkl/DJAp
/WM5MFUydO5J53qI+BhqpHhvnPbuJzE4MVE/Z0BKhcal6RF80YBSnsHCqMomz+DW
JzeK33RgyTYWpiAGmPS8P/S678Nkn/79rfCUqcJgKWCb0/LzI0V18E5rSMBf359a
V7cv5fE3ozCPbXt1bdqid7Cv20y+0FjMPIzQOI4z+cnqxa7+D6CmA+59bBS6JeDD
hK3jZ6Hp8DO9XTLhxKP7ztZVu7arnwofYiI7pkDUICKUv8+MmIKHhi3e2pB0dRBi
5zgi8qXu5WgpmSzgjSyiNK1gPOG5YE8UX1dSScYs1ZyP7UIeIv+SHbfHDMhkRxbn
LMT3yo+QHGWET2uilDCAS/WoFBd+tZQLvljwSEhWj0g=
`protect END_PROTECTED
