`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fTShXKJv9pWWK70F6ZSnCtSRU9Hi0lVon4lF0Z3rH1+4sUSgvTUk1A2utnVIGLXO
Sd8RRPGFRaONrngnIN+snQR75OEquBgxqeoE3qZM1T+Ao478iQ0JQtdWr7c6dtyq
DEEzyEaaUpbXnLeWZDxnSRyFqjVeW3kWce5vUqUnpcQVyvhs/a0IosN5bLraoEsq
MB1CK5csETQc88RpMXxMNpkyiS3Rb4w2pWaO4NrO/gHQhaYJ8P6h0mJpg6ai8Q7e
5IB97QtZKAB5tuq7eNkDZVbP6clQbFl3xGDDI1Ccj+Pmq8m6ZqwehvyXxCVZgp/d
XPdCgN4WFBRKF3UJrquBNx7hpLKSFRD6ra7xmGviydG2jSwDOnayFSj49Y5Rvb9N
4XhzswZYbk7gkIGmcP8/8qaeF/3hdalN7ASwSoUEOKoLkNqFiGvTCzyh/1XLli4F
a8EW8P7t7zvH2M6F647oymt6zhVWv4fDgJjjeLkLkZoC59kRd/ubfZuDrjtyHMvm
FInBdi/rrdT0tnxkxT7fFhB9USXXPsj5mlaoLBPxCiyf+rmJI0Q2x0OCsL0vMK0A
1IbgGbwK3nHkFHD0r4SDWpuH7/Cb8Hlq0xFDijrmy+e4CtJ5lotHMsvK/GvUzQRP
su/Nge/JNFT2c7S+Z3O7XNlpIfhwoKrYc4dp19sredGcu1qSuASp/nY27NE/mlQb
oiJlLDpv4QBHL67WH2+i/WCIdaKlYydXaCQ5X/hdVrwKK2pVfTAcDgKVBAVZ3XgG
ac3hF21YFu4ZexAvHiqn2u8nXKj8kfI4WOt4qPP52Xx8b0Ar2HIPA6JuqFh+g1Df
P8SgBqQVzH7BPnxATMCP1KIShdgS9cajm9pZy9YMjTa1Im+1u37a6iZm29uJK4Xd
yYIdDlI9kEX0HtzYI9ktVb9OufFs75jUWnn/wZ686j8+G+wu7YbQi2b9RZm5FuY3
iJ3NyATlXltLfIQS/ADOJbTQJTvTdaHU0gyJB2k1BMc=
`protect END_PROTECTED
