`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pica147UxMbg5eDAI83iwtr+PpNyVOih4knQGU835pTn4PNJX5n/J0xRjk2v9g1x
V7VL/zmHhWlBabU5BLILKC9e/j4lyU+q42aMUMTor9HC/RybEaR6ZHqAmDk4RxdG
IQV8q59FVsfJJ7L0U6x+BcjP2Mgursx/9XzEbQnQszVqm+7FKcvIXfLk02U2w+I5
Lv5UGeyKL5tmsjwW/q4/iVhhe99IVsNAi5SE0SwFAuwlAxD2FFLRhRzA+g/PA+hn
TiAJN/X05MqNujWtNh9G1lLhV1rd/Op8SbvTYmzNqDRM/dh/zI+0mGP75AC1R8C0
vp/Uf0K4WzLyyzACES07e+q8VsUlsiELv99XGFFg0r0hgljyBYt8oSyZB7zbJWww
jyRNrzg0M516tK0NhHRypoFXOlDiC9EWocpj/VgGU7h/UfESEEIi8NSN+X+LqiOg
RMmvwyIYQKGKjBRSykm4QJIJCMPjvsoMyGaSQpQ5eUBmA9F7VLuwH8vWxjaD8rNN
Phy0BPRJzMo/5F0Cj6TZOsAQ+OBCV+AhnM8ICUC0FZcPsH1WxrnqGRZUiv1VnKmC
lxeJNEm4GU1tcoHbpDIq09GaLsvRme3bbu0Hs8NiO6O//AphJoyXktqvg/S4ENA8
NZtyohNOBaLNsJgB+3Pq+uhUlfo1H4rXB6e0fha7GEjwXbhp7YZzYmncbVx+iULs
TMgH0GkZaBVT+clY5M7fZMXNbCog68ZzLBdPXiHQiwm0GM83LwP4zFVlq0iFDZCU
Rwq6FkcBS6DoekwwntUedO3YGsxe1fTXUQV3j03aeUk8+pvh9QbC69lJAZ5mxV7R
1Mvjqa1ZLFJJWswAYEICJCkQs8LX4/SrnHMpnuEc8gswpXIpyxSHXpSHnXPXxJcv
XJkKt+Uwd9inQa4jGhzQFIatcXS88vVNJ5KihU9LIIgolxBQFQ+zRYkbck8Qm6S2
AELz3uNf0neb+AEhgMj9/VC9S3Wmlx2vU0NOuPoJ1yOyEehUM/nWk7D5vqKrEzXJ
M7OpYcZf1L+X49ukhYIWIQ5Kbd2QpT3GUxUibkZkrxPZKfCJISUmuxAotUgkP4u3
9GmyE8gGuTXQWnHnQAncWPMAyHySW9WrlQ+4aAzwpQFAQQ2Z5+m3YpKM2VcHtgRw
X2+JWVatzmlJe0MdWvx0pxZUb6RVQr9pLMsu5/5r9fbxmwdFk1cllEhd/8zfF8ux
Q1qa2N+K/fnT1Hy5fV1FasdUGSUVcXCoMT/+Cv2iCnSHjYARYy7tOV0rB7sw1xP4
kwQNt3cq7Cq0ZafhYgSS+H9Fpruuq+KViq9eChMIzSCnlzAE7Tin92V6xZrYQn+m
SMkUhwR7D58TH8JvlAaKk7QVZZAZJyveqnUbwkxvUwHYs29lEoA0QEdzlW8C6Nm5
566TltI+zr2i2O7gWwAIWLQFmzEytZPk3NfaCJRX21FwJhQcu/hm/R9bFPSjpsny
0AhRoVOAh2DOGcLAHp1G2uoMNaCQTWB9on6K2EDYxURgsufZthcAguJyxiX0ca90
YtQMt/57bQeyteAnpDFsEVGLqtk9WT0jC7ALegzjZnm0yoqJr93QURXLMglGcNSZ
kb17PeTjMSMcs38UhaHqM5Iz4YbAQWDD/ziMwDzOvl34jB5hYdM15ZE3foJdRJaN
RybzvA/2z4rT/z4ndvZxZp4AarpPHZgotbG74IVmi3Ntw8vESoQGiwiXfiMFpIzz
iSZnoqDvsm13yQxOLRuTdfsnYv/TCz6YIuGgrGIlcR3S0E5fE4TfYGVyALSb6rTH
X8E4Dh+e23JSmudkYWghGgo2P7QU7EA4/duHq3kkx3zQK3+89Jxpnblf6RRagPhL
2AwSSPFDfAFdXOXaJiWyaIhKcR/YD7cqy2UQZJuWvWspC2aj9FVWKOVQDOwKUhGC
VlrFEdMTafmj1qd36neviW8wIDSDHC9m+QzlVecKi5FnvaA9A4SWj+zT5m1Shz0A
lrK/ZhPdTVBRIISPj9UTaBfUgCTRhhLw6ELNXhMmPVtiFUtBIkKMvPV31TRK0MJg
iQUqNl3CZtalFNfjlIqYUsofoHxdL27FF/0JNazIjAFUJZbcMR8K1cCStsdSuHBK
m94yvjvS2M2AQcbR8NHTDMATPybfZ1JxBrKQptuGiHRLrvKUZMZe1KVm+gmuONc9
Y3Qegppl4YXl/LTS4P40sQV2vl+izD+BeIQW+4rZTesY9SWGGlM16EOswYTGAaS6
niEuQBTjI+QJrNreanoTCBRzjzC2QxJqEs2CxyGsyNFYTqdLBhxkkBPgHpY9z3Qg
YXhRn4xhfXeAjG2cTVhWcW6jqhn6uUYfaOVAvxkYUMd1u9pPyB+stTo+WClfeRZJ
zhNlaDVLinZs+Gz8XZqTDMfiBlmlcvqs4HjQSdfW7T2Xp7kIHPqBKXrmDWbDLnkA
4mvcHh3y7zDQgrv5k9XKIFpwuS8pFfYtz3ol7X5x3NR99FiOprodvYxk3MEFI+LX
FszHi7LAa/1V9t7E7OZ8/PAWN0KnVmDamishQhtThrpVCYVj3FMFeBIKJLsEEi1K
ZnNRT85i/rgVMee2nPZ2I23eJ+TJrFXQLfg3dCK5AssWBC1W+3dpWeo418ln5iyC
M602tXpfP9Ly/BRp18H6vwnn52j4L3bOaGbQ6JIw2xtOJFP7nGM310c80//t/VYZ
mKbNKHe6sh6KjmcD3xY2SVwiFbh0Wi7+vAJbIrD+2vhs/zX/SwIMWihNh27hxtp2
RBUAlzU/PovqVTHIRosb2knU492L4vO4Nvjr7f2ZK7xlbwMbEv0vDbFiM4bdzit4
4HgR9Hhnm6EIfrXh8acyNDft+CeHo+Eu2IlroyC0LVFr72NJHFSo4bvBIKabH1ZC
IjTZF/NZoQJG3DxFejwzjfF/859+ywo395fsKtle519z/zUYn3oPZviZOEJAJwid
kAK/2K+6xYJZRFDYkZhqHRDBjwWwvEO44INcjuxJJNCYBm16RJimvygz2vvTgqd5
Lau+nxD3v28xNBUTyjuajVanht1VQ29vUR6pCmaG9R+2A1qFXLrIODkzKLArJHl/
olW8wG9AkuM9VFaUrGHlPCwiYH/Pebuu5/8E6f6SXjWRp/m0MjYkqS5Q9eX/QB72
V5QG9nMHDE9HbVLrmofJuYtjojrSV3HXhlrE+orj24v54rz7H8lym5xLCKMLlQ85
TqOnNQZxhV232W0UitpZUtlHNuDr7dwHLyiBGtygKr7XM0N+g5+n4Q+x59ZZShVB
V8oJ1jPdNUEAC8Jg3gO78J6Xd/cwg3KLt5F8AW7BnHRVlZEjvgL6aMO347425Hux
NXEXOSq7G/zJ1WY4rybSgJp0ZxZbjbT9ic2GgCAM+wbqfA8KlJ5Bjlq7K2lWT3Jk
+zwbGDI+lojqG/eo3Db5t7dfXHoq/0xKvrmyHr2Ba66N+G/kC0MUkslaOJI/v2DX
sBhWPvtvwDFTKLs7fozZ+USxqxCe1GWJaBOssQOrO+E6YNeZ4IUvgHJTosTs3AeR
T1mU8ETAXBfiQC2VOtNiRT41UpVizEYf788YkSWpM46nOrn/ANyAnGaKRK9iC4Q2
uqsm8Xc3ODAn4ccUNb1PAQmCwoks0gbIPX1bTCivMetSf3R82lwFAbX5l3qZ8+/m
/irPQ01LfjBvab7yHSOXqZKVsasJfkS5G69f3XAbWQwpIfj3cCa6hs/4EC20mjbT
lVZcTzZOHtWm0hOxdKwu2TEDYEtFwcCOzGvBWgM0JXXlimP+hppWBpFghxfJDfo5
WelWa3h6R1aFEJGJH1dfKNRxtTK5Cp484dQ2YZE71NUzQvh+Gqkepr4qUP8Sne5o
p8ckd8hKc0nefnmwlETA0JleoYiXW1l32nx07cx4gl6TLrwqNVgQUMt0cXTHEpTt
Z1DIVQzKRNKG9jAaLcoZGptHlfBOqD7b06zcCzXgszSFALuZfIP+RB8ntu0u+2/S
oOPaVRZD/f/Nb6nPxvjrsxX+5fIvb2RoxcW+0kcsmnNNSGfKkEPh/WpUooE2MJzI
U06gmL5PTvrCHDfZuZR1rQIFd8KaoxCKl4yi//VF13Vel7PA20V/FBqhfdzVAY+h
QdZ1tlQzKbebZkKFBDE7dafhr/bICY7KRM5jN5Wru3mKtenj4NMoUL6tcxGY66Dz
n+s0zJV+mb4+yOd3tH0GwmT5bMHbbe1TJ5lDkeEhaBEhs6Qm3T7x/aqx9+KJKeK6
KtEpDfY8NVTNbdNy12nZKo8n/fbRejnk+ID1MSh2CGM68kyH+TtCfWvQIdeIrtCn
j5beWOO1uLadMlW4rbF/rdHY1kWST53wng3mjYNY+rIhKW/5Ta0jwqtVHtY4aNHD
zMAPfAWBIjT+tLf87EcF1VZiiAGsE/CjCVd6iX/qkSMx709gEyF1XFZKL508sdZw
bdA99v6cXF6cJ+A0aajWsjAccrFCaAO8zDXgfCpicXNt57IL7yqjgUJ56hSfFO2m
CU0EibwH4hkwDcRI+GvdGEtg+CUSEnwkwm9yTEeNsQ7sT+JulKv2v6sl5FlcoaKC
6dFAnjnE4Jc5LB/E1UtLcUOcVn0vAHPiTGK9TlGrA2OMCW06usr4ooHwiyTD+1zT
P57AmpQC0xjV8uiI+5JSJfXWB+0255KnKEmzc1RBFjb7WUHEHC4iSjde2F3uo1BB
FI3DDZ64052SBCU6ezchXVgeMo/7RG0IAzr+QPTQvG/3JagNMa8Svj/GAu+anMvh
6MwglmrPPJrQcWtgxdtR9hHmAlA9Tjl7Z69w/xR21I9NqdRx5BqV8SL5xZ18zUk4
vfsH0/wxYsM7qAAMEEv0vSFiR+7hQ1m1Av/I3I6w/Ice5QwebYy1ew9hLBgkxmOT
0KIyVJd0apvmWGUeG7ow9rDgG1pMtDKzdC2tgwJQUTOB4v7+UJBBkFD3ShhXYkRq
qr7U4/XqAjDAcCbemBzyljYQPit1OSPcmE0/GYuWNpq7fIlD8IobVqAc0rtYRlUc
DSunVvca0vHwq9zVtgaAI5DHfEe0nyBtBSAQCccJDnsjytR34aj7aGyv1DdSH6iY
12rlfWzqNzqkRIEatJee6lgWlLxovkJy4KrOE4WePxFTezmutBd57jKdrbdTK7Z0
JE8Hkl2muPn2AsBFJ68Y+yDMHMeeP4sErfKQVVg4XNI4COn6baCry4LqpzzIILq6
NBp7YZJHjIWd+KU5TTrDKCljRO4qtpSlTRsUPWCxat0Nh0gWL53IqsK7Qr+CKgIw
JonVIxO17EXg5mz/mIs+eL+q70s90R7pkdIMr2ACQVYeAmWyGoxTDy6tNYKGJUmo
m8XUJ0X8Zv1QyrJPH/R2tSYVCmhtTfRieRbIdzhAXYk8uB6jv2y54Dz5+GXLMiFn
O1vqwEBdpNQnySaEIffArpH2+BR3yd0yWlxnByyl14Vuw50sjo87/xaf3EK1v0Rv
cVT69rZ/+cjFk8oeFwFI9cHsF9LpXUUSu3YB8lx5O2/iy4WjR3qts0Qog0ATrj4E
Xfrz3P/DeV6tzO63EfUe39FBACUVBG8KzI+JfSwTsW3k4k3I/y7nGti1XkF4aC7j
65EzIx1vmKTnbYQDb5G+o5eyCCFXQXS0MxdHyCeSkQa5M0kGfzZAK3OgnIOWPMzf
YrHvrATz46f1f1t9bbAfl6p3IPTNYleRj4nHmwmYpHAKD8HGkExrEcYeBiV3s6IV
ygwHfv6+W54NksSj5XtLUK2MgylKTfB96J5bG3tFbnOH6Wvo+aPDU7/KwiqPGTY+
cgr8rts79e6moFaZ7FfZAXNa96lTf2jQZ7K6uTbKuD1H2GZwDUWQFnhn3tUMJ7J3
oZPN9Equj0ATAkWTjb2mmNNyPUxCTJI03s7i9VxwdVJWyBE/gDPpu726aByr6yCa
oAfksUeBbkc/LEKtA2NdOEaQlc+izWSrj6mX2YJ9HvOhdGW1GOnXNbY36USFsNxD
nCXb1rb9KsuVuR11FBbOD90x9AAHIbCG5toFJJ3kYbHcPKvvYBtUtIVU7c5KkNGa
bFVJOPk2kloWU1VwMQlcEFKmXSD4PP6OIoZeaGmlzPvRpuSPHKqxeHlZSrdeOV13
2Twgc8q4OIeCoBGFqB7yMMFT7e7kvu1TJ27pvV1zzyjoXkCIyPMmwdASfwM5qgJX
6qEJpC9b27r6AsAwYq/7+Eem7leaHSNs/7PgCCpRwMIJ1DyAkdD5vKG01gB76kNB
TDtmKLC4+u8/lw3QJNFSNJMnwxIw0EZ5KHK+7BQVKyjABNdSp2GvHop1vko1aIll
mx0UDskbt5AV6xouAAZBnKdT/HJdRgZfn21SCWkA1BnyN02NvmEzxMD5W9O9JoO/
/6mqsbgZnauP0oXmNcTyoNVZVPwmSYLseBtwT+3JGpFQKOWH7fwvdtd3qCvFWtDN
d40YCWi5BdN0dr0cjsaMVw==
`protect END_PROTECTED
