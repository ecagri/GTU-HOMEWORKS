`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kO5U0e0WTBVxHW2l5G/JvgMqm4AbNVCinKgjyY3OMLlAIwxtQG5gaJWGcSoXbeUO
1n7+YsjMvfHvpefF6uK6KdNQxbxve7UjbElbNVxd5O2yakv64uRyCKmdHfJpJ3HQ
Co904DjaevlfFs9oBnGxdQ57rGNNew5AIVGV00i9SXOUZqyNBOuoFbtPYvL6G8pX
tPZ/b8ND2OXWc1pL8MPQff3HvZfZEBypXak/jsWLJjOLbJBxj7mhE3ggwlef3vKg
hM0LPejUqXqAd9tUHZVjA6xCdetodEzEEYO/MEURIuYyxzhRuME8fUGEUYkCfJkG
FO15EroC273zWjqKKMcXXOw5ewrYSJY1tGQHUYHzRl5LYz1d5F4fuWBUwOMha+ii
u2ZXhgXujAF9HFUKWsPtwD1FwVHSRAm0/+Hg5hxvVQsG/CM2fl66s9sKOIV+CLqN
akmE9cq70Yi6kYnMeUI67/BD+8R7yVhDNdA0aXnNA0kDwsofHvVrvjkiMHoZ1Wcp
MinpJA+8nbULnAsxK/JosbzxWAq30NvOF0IbG3QwLpGs5Yl0+ZmMVwXGzeeonOEW
29kwbjzZqfPivHmOA23VIOsid+lsiySbWeTjXGyQI2SGISbet99YCxU2GXhC/Njb
E9ytSJfHqtElPL3/jS+FhXgcbWpiqRueCmAgkReFtJ1yquMg5yrVobkLpjnEVA7Z
esNFFoHaWDEeefdXizM+NocSpR0lPV4lyP1fBFOz0z2/f+ST0P3Gewjt0Y5LqkIK
dQfWOXJXhkhn55Phx0PdfP/MN2ZmecWeQ/Cv0vBZNbLetm3/8ET1ZBTO3EIErNt0
pDR8FWtUSG1E7WjSX9hKSqQNgAU2xFiWQ4CfRdb0iE6Pv98HHYdGKxBOURCqy4Oi
XXPzmTKBE1yu9JdrXI2cTJweZkBx6J5iqR3uspqadwUv/QS1jD5XmWuyLkDOzJqW
xPYZargcYIV47/SCDCtz/329TC7qsjZ6g6mPnk2GCD14oi1TZiOpMWJWKScKYWuE
rBq0CnxYUft5uHepitWbuIliDyjx0tokYFT5bLgMJmnR2CYyl/GympJYFfc3Mk6q
Fq0VO49IHQy/68NNX4sUbmWZdKw6/Am4ADNYjXiU/QIsxH3E39BGGNDeuQX6feVB
msty2p9LE5pL7WdY+LoKKQ1DRuFiC9tiYl31K1Rtn0Rg0UhIo66XptzvfAdtgo6Q
yPNyxV2pO6cVt9gDxVxpXgHnDAn6F8DvvzreDalCgCkKspH9xvEwVJh3okjmUVaF
XHq5nGwUiIzKdNxb3D5MLPXHWgL/rN8/DNV7n2LgfNDknFUqE0Ejhs9gY1oDiAJq
LnWeZXK8xjbkJ2FIWr6w4LHQpfm5kvORuUqSFC+UYFWmNnGfr6Wh0LHIw2flFziH
DjPcaj97OWp6950OBNwr+nJEo2XnbkK2k7igKLBNYhsbx3IMwqwXQ3SYJFs73Blk
VJOPGNrwOjAtbr7d/upQ7Ykq21CU4QjrQA1CwpBJ9OvTftq163+9DHTGubsCEVya
DsCPdaJLHTvuIX1SJsGdEQ/O3aT1MuGnxqh1hDj+nHjPbLqpAlFeuUDwATp7bdmS
hHSuoIisjs8f/N7iV+JdE2GhIo/SQlkscXvjMGKE77lfV9gveFWG//Q21ByXBZgN
kmCPz9M8VsTk1FT6iXSNIjNB4uPM8o+c1Dpa9kF5QzC+NAWnihXpkqhb2TtFWPTE
fWCbbV7E8BDm6TctyDNW0+P3GZOdvDdMhPHBVO+tgzToh1Xkw6MpyTmwrHAgFc/z
GHi5tGCVJOBSo6vxdeVys53GLnxystjj8c5Int1mkqTXT2JdEx+fElCzJK6B1876
N5EpNeEM3WobMnZanVj51K76wxnUPaCeE9Dv1xsgu456oJnrrfM/ni/5CsPcxPB1
KWYnKCj0pB2zUTtWn6Km2OaexlJgeO1uLXtgXQ3/Fuj8k4hxoiUxLbngP+2Yyyny
VfnA+hJwEyM2U4nA0NSqbIteBN/HEffIODauHK4DLBGeXBOgOGxEhaNWpvR7oc8v
ry9RXy7ZQgrDaxcvqPfserBYC5gFBTuOs6dymWEKhQJNQvRI9zDiZcUky+gtH8wU
lq94oeKItFmM6riML26ujuvIW09BAVXh8yNeGNwe6YFCwTAvZfNyzJT0REiAnSGl
ZMHzkbgRBygckc7ARreiqRBA0PL1FSFWigCq80tLIeNPRLGJmFi07bxPxQaO2p3B
9Q5wUn3bg4rCaGWO6vxo/HegKO6bNcXW4XmYOltNOI/AyCsqrL3B1GaTh9IQJEwH
zzughgi9B6CSOBvqSkXX5401fggoT1tVCuzmbVoE77Ys6SMv02k+CiqC9Glo+6qv
B4lFOSn6yUq+CjbHGZSpwFcRghvcUj+h+lrO6CJ+dc+iyVrQ4SuJnkMNzwC4gKIn
FHSxHUkOFyD3oXcxXAJg3YbGMykYAkLeKeL34VHEgYGgpInpbwGzB5ZScpjqA/MG
lN01GLrLKyy9Ng64kZ1+aGNQAZl6SUncO9iOo3J4wamuZRRH6wREzPsRTPX7qaeW
ESwEECp0WOgXFaMbMKKRAMjXDbiOR64AIBb/RO2EqDfJYgb9zgqikAehX64CwxnN
WwTlaad/k8EIz2dTcqtLR50hQkvazRMGceEgkMRwJSq5CtFL5RY+bxrk5+NunhgH
LBgEcPJ51/X4EbVFCOep9ocKnPX0kdw0Dn9j8E2Bc1nNeK4PoTY/ldOVsJtph48l
JjQMeOa6U2DMvxxptmwfIp6EThO8IEQQuZkIUmPPvsSByFnlz1ZoXKa52vGUVSq9
v1M+s2SyvIl+6aasHns3wLLjEa2ZT/px22s91NJVVCRcBiFvbMtP123YiEVGyt8A
aQvpYLiiIF9g45InvysI1xBsWmP8xabHhZda06ZFUc3LSBP73zO5LPAg76T4sO0i
oqiAW1LPOY1OGCCvn8seh4UgCVn0s+CL1uKezGBBbYpm45TYG4nKAWDn4WQCHVJG
Xz9Wbk3MX8AKFpaQZSsECNC9Ffa+ezISGAPYUFkgunXCBFIozMzT6/4Uh8bwHpCt
Y8mtHwDfpc79aQ1yYZJNx2KR84WVq0bXL4enKKtt+v/OErTsDR9FR42G7S1meAAO
YVjPO+zbFIQ3BMFx7ZnBTedDVR+toiWPYmgDYyhLWjXJYS+2MsRlJQYi0jRumao0
Hzdh4hSZTIEgv6sSnY/JTvCEmyNlgN/zEdP+a2+8lceCW680DfwJtptp5SNziP9b
Eu+gTnSw+IjLjNt4au90ZpdEOUK+v+bcSb88daKesgVz60nWbqx0X5cM2WCJQUto
PKlOE7bJ3T699NyN1O+BVeY7dIDJrrW0ofwn0lGTdMa6keuQ/VppOIqZZcmrnCOP
/EFCiYL2iv1wUd8AgEbxgWI9vIvQbx4VVX+ztMYZEg3q3vH9vZBkJWG236ZLHVEG
ky62O2S/gNBI+3ekbmcHKGKHCumYgXfI8qd+tMQ/ZDE+Fm/sMo3WEzXESmB/M3OV
kWy2ioWdukhfbR59k0qZDfzOlm5LY5QGe1cfazZVxALOXF/6XChzpcgZWZOS91hE
nOUXm+/rAB7arPgEhrE6yRccA+3EEUumuTHHpGVbcQFrRukRewDYgTuWglIkx8Ye
Dl9zdKmycsb5NqlLVp+Jl2+axyGyurHViUcCS8vFeT6ehvsyxaovDpMRWoSXUim0
VPsUz52LoD8g4UvnBzinpx825xNiuL/cNfBOBgt5hlglVDkBeU+uijA9+2t+9ODJ
EuzuhTMCPdz6RSxxhEEAILl57ubobaNOp3AYVwHYGfk/xE87ZxWKHmDtW+Pq9b3y
uCqrYPE6wjAwvMeSIXeRcjid0soZAulsNmfvsb3uk8Mrys46VIM82hbpv+REsZIv
Cgva/DMyqCOr5RHFnN5URFW9yJY/N1j1sGzewClPK2qp8mfvHnJGseIBkkvh1h5P
06AJoblzECRBNtivjUVIrCr/c8KcrxAW57Do89I/4D1nok7zjbhMIrxZKlNlPygJ
igBZDcx8XYtlt+U9C/q5jF5uHrWPFqm8P1ULVgHDG/c3sGfZ71eWanRxYSgCz36I
hhGjWoPiuyg62mv684SM8aWmRwX0AV8RJHZwT/+33vtT8T5pO3COfcaz3nHwF3Gy
pZ+3vXxodoqcIQ3uN8tPEpZo6O3XbiOifLk5VnuVkHmGi1juQjLuItMy39mLHgP0
vNE4wDz+msZ3cdaKe9lUTr7HDTDaWrXLKNSNvIilXPZwxrlxy4kZjbwdl4XLWV7k
5YF9YzeBBcZNl+GSN0ZePrUfCJKQej94uOsBPd55z703kAm/ZSHnY/IQ2rKmKNhH
fSr8dnqaP8Z4MbFv70UqOFpwx0tmotbuX1ui67ZNrw+QjC6bP3rZ8Lcqtt8+WNee
0V+ds8jwERQXQja8tziJ7dGhaGdGtBcPOLAqsQjw6v7eoCXLZktOoK/+HbHbskP0
rEIDdYG5YktTA2/Aw/quQu9Z6K39F6Y81NVHf9ebeqwKYMHj4vn3bB1GrnlNusqQ
OHQz0pK1J+1t2BPj1PKv4te8erg6XvLzGmlp68X14cz+4sO533c2kfOlPmKg97WR
TtPpAGGM6SSdVRq7o/LsqJ1pMSQ6A/xsjBZMIZiNjbvS2W1hUX14oNZCIyO0vTC9
2FNNwsulj9vugZoBGjdik0cqZg7kVYP0ZXYbbBNeyV3V1XhJekGNO5KeiHRn2iwi
OVO8hTRFSSumYehlmP1UfYwX9gMs8w/I5Km6iniGYyGoGVqT6G7fWbv1pTLlPorb
CqIXfwtaskZ8zqDWVFD+CRVjAqiEdCh9sL/EFQPMBsH7OOfZNpPAFXwoWRc7eV7r
RD4a/L0UvUxPP8BNwOkSWbUI3Xv3rQUXgXLwL4QNdV5h5bfr3QuYYUkUpzA5n+Kx
/oa+gyAG1u6lglCC/7Y/hRsZ9q6jMIL6/9yKkT+tplYzpAL6d5pft+2VYlmaLMVR
JUz2NrYRnMVbKF/WNBoTZ4LTK8RsqN4RpD1PvqX9Cpbp06GHd/vwS7QCqngv+7hr
KSDBGNqMs/jUCviji8mef6ehoYiniyBPZEyt1n8JegHy0osGXNn7zRATf7VXuUFe
xrQNO4icAjV/kBbkQ8wNg/Kal5Yo1twWSwAmaMSmwmz/tTFdzYWbwnW85Z6mdJ6h
3X6ejThVg7S/vDOf0MWQn7AZ6F3PVerVGeLU1fx9ahC0o7I/Kdpoutb5Vh9CzaFa
dKUEIqqfzXWV3dfTDyhAkTV6PyC8PcVYYss9dtYvUl3FKReQE4qNY7oqoGWx9lUg
FvBorCMi6C5V2J9LxNQffQtXDIaNwd5iCFj+G1YDaspIiBdr0Z30ATZ/oydvXddf
DIpA9kVDvK5wDtmtSaUSJ3kTNwjQAuBgEHVg+ywY4L2Qgir6p9vKZYLAH874Y+MV
0VFZwoDSr7j3qLWMPmsYbQys4yOoX7NdWRsujqTEQSbct1eeyXsgmPckPOX7LUnK
7ZblfliU5yFX/8hIP9pGnRgLhGyAMSe5uXhBMx6gVN34nAGcsQ5I7hQeTv3IZmM2
ZH/DB61p0HYd1uxgsCkRepfTIeoZwRKPMXHJX0s9G4Tehs1VOxCBFup36NwigtDg
783yDVW+aVFpWaKAIluohQDS6iXcOz4OY+uyHy6UG3MGZCRogAyDni/NWCI/+332
3bKHuqpRE7hKV0nUZKHJ5EuTZuA84PR9rSkyaepkHoecG7IKGHRz/s6vxzHkvkwC
oDIjfMJhzQaIl73fcOT6noabu8kGeYo2IOvQid+aon7ScKvfaD1asFz0O/KYyifj
ei5z9Ql4ufk4g736hulnR2DotESarQ49HwFWB6UACKr36Fw8gQTtEfpN9YwPXoD4
WsFQ+F+iUZOpZCTuSreIwJwGkphmXJD6jbic5QLMXinVgNufrISv6hx1fp/ySIuQ
+YyPmqT6O5Wx1MdKgZRV0hWgjX7gD8S9ODz9Rs+/Zr3MS5402YqvvHldwotD8q7l
u0av3aLO3e+uMpBlANVZfyZyRRmK3yUzYRFLoBmw3yayweXoKX0pt7adW2JlsCbg
DAqzYYsr6P1m4G5lQ0INx5FGS0F9ew572qmi8kSGD+5FX+VcA8xjR5Iirtr6l8mI
s9dkRwe0r6sHEeFa6f5CiMLhYcTR9o0hVtMg2zUYg47rSE1djIv9rT/dRa+4axFz
RfQhxguw+qgEDjHfi9LXNyut2G42o9O0x9U4Cxpf7z0YqHaOmIBoMqj1qiH+cYGR
uhyc6Vkh06aqB8tEKDplC0JOcbZ9CfViEYkvefHQaE6/kHmYKSaql+/ui1MZ5R5K
Xt2XLBKK3xi7pjBnvQHn/zfurW6RUQjwhToS8MpxrlJ1VhUsxcARNeRHsjwdcIhW
JWGfKbG6r0BkTyGNqQPSMJWY72LIpcfvMWc31Jik3VHHXGAMPE3ix1gSRHNuFNiG
5YYDOEkxcDfRrM8+jQRVokBT/Xx4IS0fkPgwFAbc0BjE2K3sow+Jx0Iwc0t9XASV
2clJWzQGtkOpz/FA/dB+jfEX4OX2J8E1gbDJSDcVfszjWp+Wxag1ZE0ZK1NGvYcp
6dWGnOwRPtLtT6jUENmg6V07leXXegZjoJDDzumUuILLPPL7G24aFxCxBUhoJddS
Gt78GQWP4bPbr73Q8+HH7sucbRcNju9+lzrg1dH1sg/3G/wATkk9EzoMtniTEABa
ee9wVaQYSDFFVTyr9BlGj8NwI8b2hfzeUmzy4dBa/320amTeBkY7nG/AJ7uPOLHo
c3EXhSAuG6y4TqIwRzm8FamW7+Zg/4IJ95wcaz1TvBkjd/n+Jjp0tpwDNAdwzEJD
WefmSyx2O/HFSI01gstZAo3w+bHQpaDLM+NRPUi3VEKyIVmbrQKMFTSSwGcY1kv3
+IWQEGkp28joRFM6Cs80MTfX3ElSq3e06/vKstpcO0OsegsAJd4maTxSrMRd020r
9GwEMm8Axndw3/M+9+ryTFCerykiABVcyA3x8Wh4v/E8EWOGMKKi2J0qBkOV0Wl2
8W5g11k3TZBLUgSIX2sW/47l5N+F7kwlKurNw7mbL9hfh7irSRcUnJ2/hL3YGKpF
YpUGIKeH0fezTFok8tKuGn83dRtNRvYxVRklQZ9AMqsIJrPnpKDvpYPRF2ZDsb/b
SXpo1hKFGdnBajeREjSbwJ1WgMMfcwGYsSFu/XROmqixYHzuF9YyLvvQlQqDjnrV
v9nOtBaVBpuXb9gb88vhz9/S4dxHHGN1BWiOxeww31t108qfdxTyX+zr7fUQJy2u
o6up/l+Hfo8KMWCMdDXPJIIbW5cMFGnQ1dK/wegRi91JWVEI221uOrg3hhJiH0K4
ocnrvrekNln0IRJc/c5G+wmpOi65ZZahg+CWHZfKaSo/8xEGmtg7WU1H2YXT1iCL
0G8t4AQtzW3wbg827xUrQMlJo8lKyrinVt5D0CjXZ6GPFKw1eNIW+yhCn9PaVeGP
RUxgsai+u5bfDWLOfV5bAJIeFn2toyoug0kcHmSQyWS/ADu0q+UeGXbkhkfWHVcI
e9WnuLDPEEiXTb53mRbhwq/fx5Ximnp3zc3NaTARQlxYvxU2vYnDOvaQ3NDbxFkp
A/IzaO5s9H14LN5Ag+IuMYkDFFLDgLlvGBIOTFroMA0uFdZdhD5AQBF8aoTB9zDB
w6lYBCGoa7RipSAmx8BbT7tGZ5yUFq65IXxfepx90Es0FR4qy9WZBtPBJRtEvjiM
VWvDQhg2oxZVCIM9lotomolRdELcnwHrJQtWH2buztm+dChVtb6Gmf2Jb5jQa/Yq
AhAh/5MGQXvmpuLSLnj78/dvM2hX3qVkP6S36DDaj/I9YskwpEj3RuEr4dJwyOzO
f4sjx7aOWWxpGZoEn4kZqXNYq3ivf/vgy+bzuQ4Fuz+RvdakrIoE1HefHf58YmMu
znX/U2ZdLM00L5fGmczPirXplt+azWLA0ugTCROHMHvdzKoHdjEqKToi/XzWw4z3
XlQW0O+dlmHja2kFtj/z3gPEIp5mDZFgPbwqCZ81qJatNQfE3shcfijme0fNpQ7y
ON1+7JQgrLMZU40ss+GZYQFurvaDShTrXGtdvsSnp2ryq58Lp7jOKnAjWufkdEA9
HX5JoLVzOTUO6YSmw7FmtLq39g4Z1rpoR4smtI62mIIiNVhCJAGhLhRLAsLY+bPM
s9SIFppdKAT/TyujBjpyZUWuVJjDj+Dlr6J+ML1jbYu9kq81e/E+oqd1JbWcOhHq
8QRVghMtphCwZh9gRZINrrIoSkGFm4bZFUyvMyECOUCJ8K7FgQpp6sDU2zmFyaB1
2XFw70/7MALkLEJygLJEoCC8f/jzgUfakRz0MNRyZxP0jHooTEQve06R26yEatco
8MLfL3XQLgKVFYUQ9wb3wMPIO02kiSf/Kusb057PmuEBTcyvPYxZm7J2zUxf2Ndj
N4o51aLLvYOcBBR1FUdj12PqY6UG9f5LqPI5JyQVLMZJinl111z/akBiTWfye80h
D0HXwFyoghHCU01VtKH1Wbh0dXzgM1196jvqS9eTZBILgTJafrhb6asPbRvSd/79
dFQJbA8Gh8b0YfpROtS3Sg==
`protect END_PROTECTED
