`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PGTq5Z5DruvO51AEx5r10L/G6rQkRiuTSOgCjei9N76ueRrPCoHCBiTH8cRs5g6Y
cNcVJIbkDqxyaoTER73msmt2NRbvs/ohXWWl5gZgqR+iYQmcjyROOTytC+5tuJSP
XFBSHMx5ufOb3AK5G1fgg6p7Qrrha7VxBP9Zz4vBzOzNXmg8/Q+cNfnYAw35tj/J
nBdy+pkq0MJ8/4L6G/1zu26tI5IjS+Fg+fDymt8wYUTzMl8YZigUeijk5SUvAaBE
tk68UL88IyQrJcw+/B1wuS1b2dGQU2dx94V4f24HGwHRwoyPCc8/OyyWeUHML3Of
a+Tu6/wXa+GGnWfr36JL/9llPVLTy3xM7O+eyaOtkRWFcb0huwxX224vNHZvSs7Z
vDKDIPJyvcp94Je4vLux8jlNldSjYiFBEwwsuno9SWFV+S5dSq6XWh7ZBDQzIHzO
26UeNJrzLDnZOEl2dHPgH1kzAbtGsUTWkmxl42mtB0hXgmurAsq72smzprn4iVBC
R8klInNg+WihdNSp4IZRMCV17SGAtquKmxv7QOBFUFub3Ze3XqjlIERlW85kKYc/
5CNi+VQYdPhlzUvnAeoBe81HVv4QgxMMNkhQoAnIsoYMy+JURf3mXYjAXG6wIjJg
AZ3DqN8ZvTXSIdKk7JXy6M1kEmDtDBf6msBfmCWOUjrrMmkC1Z3pNFvoPdgxmoJL
W4k+o3ve05WnCNDIwl+g8K73vhod1qhv/ZJcpDrMbGGrDu9KaBShK2BElezR8sMS
3FldA+PMyuFj0qDkn+zDu6sMlLocMCzsv0fYJRxYsUBH9QlujixwL6GZE+lpkq8J
`protect END_PROTECTED
