`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xqRJrJHk9af5clcbTyKg2rFnmwZ/jLPsKrKG93wLqZ+oKw2XwtDFTb0RoAyZh/ya
Ug50Oex2XIFCyD6hckLTbKsJUul0IM4UMOmGK+a7n6vpFMqTbZIaZ0ESvaHNoXhK
bTsfBWw6va3Qa1FNzND5c1PQSlLV/0tZkuPzlolUAHX4v9W+L59Oam0e4pngVRen
rjoKY3GRBmWyo3T5p9fgvRc7XB/VcKaB2OhBjsBATXtlhpZOQJqkWJxg2rCIBr1d
Uj8UluA2jjM1AsFUlNoIkE4VPcWOtjcwWqW1CIFs8u2ZJhUIgvtQViQ4mWMo6/GT
3jdUTE0DBCoc4b3rsafzEQkQuLLiFbnZtqmJrM7lyXQCRfJChYNcrDREPaT0yuRT
G72Gjwfavx3iPwC47hUV3D84F/I3gbVNfccwhT0sRq6GBuHyuD7UwWdsSMEEok+J
fzrhVD8OqN0Ga/mg0YIgJxAivMC3/cSGRVd+pNjGQCBDI77iRJ1kqZ95NhBU5PWl
bOSxIr44OC/RYlwbTJ0cpiHUFgvu5O6ub+I3d6SLtNB2tttz208IZFE8re5BseQm
oYhWvgXfDbmXQCcoAx4k1LP7ADGO2jVObZMDpbAw7oKuyrdatsvHYEuu67M05uuz
wdHOyZ3t11cnrw7hTuGiZBDSnbQGPQdmo11AwtcLhUDoUxsCwejc9AKoy1x46HMP
HuO3hqqoFDObdhjiYCyh3C/anXoRAV6xUUYdeqC1QhwRnT+WEcl2n6qzrMEZkiKs
oYmw43envtoMZOXTnTdvHHPza/f415280EfjgAUl4SOR1EakiiclKF4nM7xOxzhm
hmIzUpSroCccN8J+zO8TZXR0ATO+PmT3j7A3Pl6rAZkCw6vDYQy3cHan847f9THV
`protect END_PROTECTED
