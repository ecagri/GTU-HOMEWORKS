`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xPxdc1OzkZbjzuODCB+BFTlA710CyAUFLs6fvj8esT71/RZiug8BKV4vHeM3A+9X
CpLP4c0IR4oKYkQstCJfWZ6kVMceog0v1gsphJ0aD5ViYgPwjuh3rXK6PRZYApcS
EYWMbdo87F7Ws8IB3jyWVKKVhmlAGuPitDdMNHhfXBKSbyOFL/f7/wwO69O1Xn7B
7ptSl/AaD2EyvTQUwv6RESXRf8XlBerMV8TVVG0De4OWz/o2WTt0nbwAmj2uAidW
hZB0K5MDOU3EVG+cS7KYLsbBsdb6DZwVZdcm1WkjTmOt+tJ+mv40HOfI8Uz5l1oe
s65e0pTw7PUpQ8VtSCjyFjm+tIkd87jALYUSkF0j2Fy+3eqUDVKbyjbDikD3IDY1
gt50n5M8elA6TaL3FNTBpiqcRz3Qjlz4tA3ARdx3/15dK8XXVpA1iwxPPy868Izl
BflhlkHbHegVn9HQVKX1aKEF0BHwbH6N82845M1zIBB6YguaJ94xY/zgHpl9qmCC
557RTooMJaSbnUedqFTOhA==
`protect END_PROTECTED
