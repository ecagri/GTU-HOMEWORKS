`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DtojYxEkX3iUSqov/jNe9UdP11lAbbaLbqYh2pCOQm/drru5dbTUolON+e79y3Z7
0nESuNyaRnQnY4MqHPh4/dpeYDyl3JaPzWHs0PfCxddG2LDqcPUwWkFPHSdrauht
6TOw9cgQldrJkBKBCvqnzlVFz3jcSzyt7S+8mTaBwR96rHfxV2ohzPfgFiWJoyET
X74eZOKROhU5JNlRyIKM8di/6lLMGeT65Nf7FklRhvUHyeoBPobtBbaD/Xf8US40
Y7TIKBqceR0FfB1KfCykVy62zjFzIbYlu9HQ77HJp3/sMTdGoFVXBzOWCtRAzQvm
NAI3uYqE+5YomV362o9GkaNEifMmOdsFpeeXqr9FB9lgxearHeDA4H1AieDNz4pu
cRRpnE5mAiZmDYyatlQa324hjZgiSDthO1MEjtaN2Qp9c649aznEOU0MqWKGM9o9
mpWQLYlMX4gm9PHo4sHooKtI0NKvAo2HGhkIVl8HUMEPXH5cY9yz1CpMMoVd8xzE
2OFANa6e3L3LQ5pHnTh8tFvM5lGJcKOtZhrvayIVoqwcwANGVjRBhKKA4cyoZbXq
XLbcpRDaAvc/IxeeXSSU1uZujzk02QwPGVNVP+iT0kqEBUFMpy0LYJzulK1Z+RZ5
Xs799OVYk8b5TUAEP99mNLklmlxLUL6VLUoRzO5nLVNesTrKzE6Gbdzqgx8sEcBd
90PF40D7WeGbrPEAIRtb7ZU7kjKeGzX0A1AW4H9atB6JaIFixwztt1imvhJRKjgL
whvZNdMoD9PnL0Pfmg7SJbKrJlpyFlDUTpPK4zQv0rNzUTZM3bMcT7oE0XlxjAdU
CIMPlJVkwyriydWBN4PsPjLUuYVLyzhaUrsNWNWXI4HYILNuMs3XK4E1ujDR3Phz
EnC3zGTSQGQNlz+NOHGWwAR3iH6FFDb3k5R4xq9RCxk8BEqGNFxkk86TAaqj2AJ1
GjFFbzXtICwXlCNlQY4Y8p9KSigXMEHcqrzwYTTvv+bFV5i26I3wyEBA0fq5sbhj
cIrnujwCe76tDVrzzU/DmStSzreFRrnO4S6/j7677Mo4+U8EnVW6bPt+FeItQvOG
pRDzaHRX91sBtz7Pdpjk4J1f8aVdAu7oYA8IMLSuke9N7Y4e5Mm8q/zO7ln/J7gP
nO8llZu1mhCFTBnlrkUJn80bpqFfUXAIkgXS5S1fjs1nYI0CmffpNlcKSSYr6cTt
0fEfuzbN2QkSCJkIWN1uGb5ZtrLzcIVFNloE763QDzc2SRy4GPmY9/gGOQGGv4bq
`protect END_PROTECTED
