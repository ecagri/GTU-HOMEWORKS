`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wpE9U8zVeYelWEGLoabQdIJuWENF3huZBmH+JNWg9pTRK6Q/lFliUMa3dAQJljf4
VClk7cxmfCa8RCHnZjHEIEoo+a2dCMBQURDFr+9E5TgheytTBQbBAYJ08CCw9fLL
t41h8zx7dwPh74ej7wvuB0MK2Pp6wyW0MZ5sEy0CAUNfqGE5uNJ6yAPh0tdK0Ed4
i+eOdRyBukJ6KUEf6EX5PZHem4qNLAWiVKggIveubwvLVSUMhICOOPUTjfth8roe
3VDilh02OBt4xbTrCrdbD1HKTWCgb6bMyqtVdJon1pqOJrhkgLz32Y9jc0pQ+dvO
Hq4GM9Mr+qZt/YQ6jr7UiplSIdKEPHNFvxE+qR+wUf3sN8Hg9H0BmrgbWO3ZK8mB
jQdbMv7A8iXCWrkLUOa3G5cJJ/fIGVr5q8IbiVLB8HQV91101aA/nnVIAEgKwqGM
IejHcdcFRYyWa4lloDq7xM95ZC04RT6Q6oJZZYMvtvxLTERtlQ3iQn9nH4m+/FZ2
ZY3PIPYFQyUZ3eSVDGu8c7+0yJPXN6j2w0gc2OotxD1kPY6jWK7bV6b6agHCHY1v
kJIo2e08LFShz+HEFShQAyD6VpYHPD4lWiJO8dodplFpLhyxKv5vHto4D9Jt6bjN
3sZgXenvKC79J8eEt4QimUQUPdr0gPzc57Gkmc7oYQUMeHGYTCVNbBUS1ods6yuU
W6cj9OtaqjUIYH/Ndfxf54HihvzTLj8gKDVcTYgfroUgzrOG5TAVjjJvvruaFfHh
9Ji2iq9Fe4tPSf0iSnpSQCMVl3D8cIxyB/z1xzPRWD7JOofaONmzpLWR/IpU1egH
jy2TOt3qLQRogtLogW0+SeIG/FvZOkkCiRU4U4jV75ZjNBUhE0wXlnO9iKLcn0Gm
PRW793qYmJ0+W93ANkoKmaaRhvyXWLrpht4WLTjKnyOiE2XygOTLRS8qGsFA/m4A
VQ0uoIdUxIssc7RlynSYiccY6Tfd+81lePJzFYOrNpBoUgMx3NR2KfTZwpP0ffgR
u0gK1jX7ouer2fUkIWgoifvgnCYlUxrYwrYY4NGrPxdm7BT0AIWfxEH2iPE7OuMB
yD4RxCBXYZoGuNdmndZVEyo+aq+rv6RNcZRreh2GjIBueUf3xsEG+YrXNgQnJn4t
2Hv9gyy10x7blz4Cfto5bbn1PtMB308Oo77vOVhx+j5Y+xHeUlaG+w9Z/+AuKLhe
dgKUFBZEVTGMVF+ThS6B1K3r0LV7Y+raUC+HtXecLvUhY3WlQ+aukq1EG9aGJg4d
XpvsUj8DCuRUUgEqWHgMojB9BBw0uBqjAxz5iwsHgk9PL9EZvZhAoI7Fa2N8t2ay
BYVaT9hwJvEcGWdM/k/zOJODbMmAP6jC/Kp4roMNZy3TxCMtUEn1ONbo9lCzOANA
ojw+SicSvE3idcZLtQohr2iMU8VqFtDN7XQDhbVWCWeMnCVVsvV7+CF0/WxSnKOh
fN6AUocBCz1nOF7N/tFkk4DIcBYkr99xhWrYZ+07cczfIT/qNaovPnjJyJMQYRcS
nKBcYrW1BDFaim354mRoh1P57GD75sBzhqE2UWEh+WOlgv2p8qlTFzeXggchV10h
fvQgqvjr9iKHO8uddpyThof5KYed9vUog/y1/8L67N5b+zO4HhFfgm/ts0D9CnlF
3uicPbctrMOCbj/gDkghlfbbygpT1XgXyEGjJQTeePnwQG79cJvFLlfinxRzuabn
q95BRHTSPnyvl+N4DswKhSY8kBURiHU0DsEGTH+kD/Z2NNwYkoDlXSQUn6YLTAMM
Z6PONgqU812FaVY1/DCZ2czkrk5ENuzGfxg2ETgjfcalO3yW3SmpwoxUc+dmXU/b
l/t2+YqnUM0PJw8s6eDN86DXdoOURb3N+ymOj+kXMnKhc7kectrdse0TuutHWSLA
qeU85KxHb3uNR1tJ/k7/vQ==
`protect END_PROTECTED
