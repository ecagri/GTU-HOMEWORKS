`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TVmAB0hJAxsj63TlijhwnhBSdE2S0rIHfLaISQwcsxAvDBIlRslESL2obq6BOUrg
tAoDJPawEO07mYJRWZ6Aa4Y+NaKB5cbHzz0BGI046pkr60KeSNxSFD7FFXch/kRG
Cn8B2HTLOa3+5K6QELV/FpSg1p5md3tTJ+yt47EVRyfY/B7xgszEghpuzz8An7rE
/fs3PTTyZQffuXl85+/9VKV4N6eHXYeO6Pgkb1E2othm5lxC9bCRLsDXegNnH9/t
IBZbEPwjbICuc3zI12GaxEsR9Ghb/QI07VSqWVDadv9pHlyoOTmKsDGD2ho9rNa7
7dAVYaPQrNsAiaEkUNtY63n9wJ5W0LI06EEhBKlhZqW3Fue/XA+eTRjo+lTwo9y/
LPLjY558pjwfvmvAdjr03IuHDOnp4PkVyz7W5KUPhRFZZlF/SWi+fMfAj3KBr9n1
DyFlgB+90otQr5+07kmrRlqzkl8qS7lpEtiuYGHK2IpXnVGf3ubazx24TCfOw4qF
oc5GfoCM3ZV+Y7VCyREjGZ1SMW8g7YLotef7aoyNHvwNRJ3X/uUjfORXymeoGkQS
/sllXi8XjOqlO7P4gw9nauLwMdZrUl31EwMfgjXHZlG0Ef9jQHST1tEj2EnEI3bd
hUC196BWWsVyEKzMMAqrg47yU0U/qIW5M3Ia/5KYyCjQ0SqCqXVHfxIxtntyj1EJ
XGNjdfzaw+LoZYE/TWhWMEIIeJ4wC6tsoVxcxzJuWBGiM4IzPeszV2gbG/2yFQR0
aUxEBz1Y0SzGZrdgxrjEj+jn57OJ3gsS4qgOtZ8eznWg2DPHx1lCMqVfklZxYsGr
SNpTOU73Eg96FKBzt3kklJwnXyF9nnYd0kZP7dN0V03oP+PxCw/VKTs2reyTGMVn
PQhOJOWzqcVRMj+8rRl4BNqMCHWrznKKJ+rVMMeWcCG8NeuOE9busZ6qUA9TN8AZ
sirGddwZ7+uQpMAGKG+RRzZ+H70M3+GLMDeGu8LQaaC3sq3zJlYpxeV8tsQa9Uuo
iKa8eP4otwxf7eaj2/rvlw==
`protect END_PROTECTED
