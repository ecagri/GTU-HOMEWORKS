`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KQcFIWn1NWhMWRJM335NZLM58aJ90IOWNjyLHnm4s/k5MCgv9FPtzT3u6PEcq0W/
jY7wbUA1oJwaxBt2mRfmMCEkHJZAMPR4PbkYiKxJl2xZbJopBkbUcuHpPOhDs9Pj
dWb44905J1x254KH6sdLuR6ktuQ6MQhvuL5snhGlELCgd4zOKqMTcK6giztAZeNR
HQkvtXXazGWA6FEb4rmD8qlcQX+rXgnuWLBNaKD0A3ZJ4sSlcX2ZrDnxrtvIiOm4
E3w/39VTDFCTsODDb7nVdKmL3se/g3uM76m+hRkxyoswcexpqeQZZtYeTVK/dwWS
5uJTOf/ZabjLpeONPW/y6MSbJw1gDCtzYNvTf+P8c/R6P/ogYMLOAmHDotOIxc3M
lCK7VqFQyWsvxaeScTkcdfL+LxKouYuYYjr7qLsypeq8VTfGsQ5Z2/TJhQjzVW3n
9rF3lt2qV2XvtUmqKkZCcsesTIK/jJJXXCRfk6+2GWiyEofU/qzcf3vbCUDck1kI
w6vKLaivAPzbEgsE8wO2c9KY2QQeuGFs2CaePJu93gAS/NwpXyeh2EpJlCb/VW9A
k04ByZeTJzn69ry6PTs0gMKtgabx0C/vTkZa5FVtSrIrHFlWGom+4jMQAOPoVOto
JBVeDbT0ZJ6yzFmuhq1wUBneqMTHCbH6b7pTzrnV8WhwcVHVNamN+e94aTpnQiaQ
ROui9ZYBtN9KShOdHds9Tf+zIBIH0s3at3HK9l5J4LhkIO+Q260OOBmw0SEvMW1+
CYF+ceysceRwBG7zw9rmCA==
`protect END_PROTECTED
