`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E7QAAs70EOlJ5ZPQHRPhRyuA4gz+DOBxvfz0OWaRfycaMFP1igOy7eGrS5V+izG3
kZBETRgho1tlaD2Moxe5cXIkiiF/Q4XHVszMnTqkDlMmZEaho9b3tPtW4QYZB28O
SCIHO7UyiT1un966mOz3sy08ZhsONfPXN2Nc83pEGGoZHJ7stTJzg3JDcxRKKFw0
x0NvpybTCRa6pd7oF3QQdSzoDFR0mtQSHukLVIRx7nelFAs9s/FRbCWBN2ERUMWi
zGN70WkKEVoJU9faBt05hTgQVpBGE/l44eBYH6Gdgk0eMcWzRd6C2Kf7LYcPl3Z5
FXSEdT2rCA9ygHrUp+t5+iqMsZzAEXSD88y5xSqhoETQ9vFGcsXmHiy14QmRidTB
2kp1gD5/kqR0wGkpyVkNyfwauB0ofIiLE7HAgWNsM7AQ/tAfor2La6ZM8DZM6GVQ
+pQCOMEae0miqK+pbtsmyNacrF6blDJ3ZZwbXd1CV3GidVFjNRpWDOCnoTf5/4mm
B5uGhLoHEo0ahQKgH7I62srEdZXKGJUCGXXVswmE+vyTsiXVNqyV09/dUingsKs0
F1uNG2qO/alnMpTDbTVKMe3Kn4nV4CWzAlXoMcsM3BI0gSzh9cDTSqejWOXjyUPo
FsYsy5lrkkpnROhwBsaptn8SM9Vqrq7MkmAH+zZ2d8Sj4w1HogAC5IG7XVl1RfPC
Q04S10tmkaxvAxvXiYOME5+J04kpmz8C6Jy0LSLGzKgz6veOl/mumTXDSFMckNG9
RTEsg6/gnDxhve+5VZ6d2GlL2cTFvZuWPxQmuJt6cBtnQAAXbQY1B7tXfcqvEaCZ
ghBOD5wUSjjzoS604p6P2i+lZ6xN1FclsGjovJLHpJVGvUPYkAMA5EcZb651j5ve
xgOmv/0JvunFEynDqJuLTD6LPVPLSNyaFZmK30uGstxpWWLxZJI/PBOJzXZNvYfa
`protect END_PROTECTED
