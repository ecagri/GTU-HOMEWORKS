`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vr2pxmJzw0Y8LyDXVkPVe4dmjdm+gs16Ct0RBlgztXGRDCHuDENS28TC6lFw2Q0c
5gHeajx1YF448pdMKaY+IjrNBP3O8TWx7MyRPzwO5UM5QOPyypqJ4Itwf7UgsWLu
ylAWaTAen7HxZN5P7FFfLON/V64JVdBIIu1VBL0RZArJgyloufdxVGRYdDiY3EdG
U/OchrToOA4bvh6ufoZ//Msng3in1NR7cGFqHpFv2VwngUQ/QL+xNgjVLMa40Krn
oQ7UWALJgz/vme7p90rzOl+ZVe9uXz5FfppnSCURawXiy0E8gWjezA/V7tpH10fq
OF5DvfNTHzvguPtJ6FqQv/7DrzyM0WoarKGcMOAF73ENk71J+s5q5Ct7pCLTMB6G
6A7U/AVyQzWKnSn4F7yjZOt+zFHH2UKtBxbKCCCCHheag6uvR9qhu/+8YiKfikRb
spp81RzLqlQicO2REG1gD5X9L4pIkzDQODzcXJtdHfQE+zhfdwp49pBLY7/W1KnH
5jPRXIELVMyQbv/V0o6gk6qRnJJC6WBbGOKD8MzUIh6PMtDgLXyuq4ysm31Jt+w1
3Z595RJKmqCRhqJe8PWSHGB2dsCRbZAYx+hf6VztuMJQriiRlQTvppOX31IDIS1u
Ark2rZgJyKbSZJHl3q3AxOQdjzaDp+m3SF8Cvv/CcjAPeoSLGheJwJ5QU6M8C/Rp
EPUZJHoAqs4OzncQ/FnUrgo36LG53U0MRQ6Qm+mRihF8fUsZFVZe0SqgjBWqkZFc
qWilSEH82wiSHkG0OZN7uVEvIkHgguURtaRooHfnfrLrw8ahGBtn+0guXVWfJN7H
xrRMYeQCtNuOEFvyBuH5uW2UkmT+XBbW+gTpQBu8HEHIehJKdKSaAzxS3jOQfP9e
fc+pSp+8mne8HF+ff2c4kKFl+Y0Kha1SFb8zOCHZtNs+SGOdZ3MKNLqbWZrQYgCS
nnmhlX8j0gxPLpYHcYgDDXeozBW5C8dMU6/hQPRU+kQFhtwzFJQQTqGBZHq80Jl/
XoXC63Ki9ZJ2rCAzEnbBUIiubjPFi7q2k6h1uCsl+gGtaQD2aEoePJIorgm3uIaU
Dikj7jK+sYgYu74MPHMAFMMqjblUEna+71z1qc58f9edIX+6qx98vIbJZA/8mpFD
PscM+xgMpz08ES+Yzch0otvEL5krnaLDGug9vRWpYMZZ/RelN2iEIXndfK6nwTQV
rngteR0zfDbbjJ9Qk06+qDdAK2oRCzEAskFBEKWDy4QQP/6PKQ6mjuLJedo/Ie88
dLp9F0xsvnPnvI3d0KfSiNzSXgIAhXHsTWB+/ighwgKyqff3etWKWVnxBjDF+qsW
IGsC0tjwSmUwHf9xxubDwwpbz21zNGSs320u58q1Cic6gnmx4RDA1aoWd7MzSwAF
S9KdeUdzJ72naCq7VNyRnTjN6Jy6ZGOC7jCQ5uZFtnhJ8WtPkJRB+I/7EegJlGSS
PgHj9AFMsqDGCOKQDO3tKum5GH6pWR34nZiJBFUCsAvsv1+aJXiBZ1c95sXnXvs2
`protect END_PROTECTED
