`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/vl9e9Tvgl1fD38iO20i8HQJBgp0MDVlRkK7T1muanzMjncYs2RCD+WVhqqLfae/
Q8e7c3ye/ULpWW3kESXy5XJuVGBisGmHRWpP0/fXysk5gmOe7BuD/vPsxkIcULI0
06v7VRzZM9WKWyV6hiDJFE1Zlg6LISgX58xoNa1NpmISTAs+nKamcoAAvymNtZLf
mQNzxMA/WcX0qZZJnNTBo9bEGw4a/3lqc8kNAmTBz0brc67U5dE0n2qsxo2kSSlC
PH5vGwoZtDoVXuh19+1ZS/ZL/xvldi4AKYFEzFELRKFU5R0BeKExgWeIyeKY/Th0
T9wwmfL2ProXLaCmHnptJCKiqYf3alr9vZPMl8nDP6m+I7KxoRcYl74LsQaJCt7I
ycFIyRgUGBTG5gKc4eBPwlQ4ILdVvwocsEwOSlQBuTO8Zgz6pcdKwKs9dcRSV9WG
ATauTRZvay2EKn7nfZM2yIKkZ/lYd/blMqPBYg1SS0U=
`protect END_PROTECTED
