`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UbN29LDpYb1NvqRL+WHxdTv0iDyDBMbebF93WKiI4/DquJNrpLbbX7nor8Vqdq3u
99hV54aI4pf95uC+jI0W7wD2AYlfhjPRbC2GytMtebp/bMa6zL7wAUHJzPNrCxfF
KoNkdn4dBTaZkakXWeefugD30rW0w4+2ZM0GGW2N6ehQIS45Zpp3/Gf7YnSF2A03
Rd5Dc1pRHbhj1kIOHJfIxCmy/ea79El2nWHIhIFSZEHsJK2J0iDhJKU3Mo9q7wi5
8oWZugWYBPexFI0xZtMApBzi1YfLJ1bkfDIBiazXJUG/7pLU6LoCSgkSFV8zM0Fv
/PtXn4tUEr6gs6bFoHfoFt16ir1ONak5neUGu6Y26CRuRWltLocavoEFwinu0hei
3VSbXerXQ5RnU43ZbOLXoeNnHo6Gjz4H3uwdQAE3BE1Xgf74og0nF6VuVvBgNR5H
htYel5UDQNOb70Xl4jI8k6ATjjSDnabRBkxeKguWBYI=
`protect END_PROTECTED
