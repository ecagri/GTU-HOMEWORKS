`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mS7/eI+kN3zh/hWiDczyUH36E5pNceE/NedLFBhOKMfnFOF2ee61shNZ6a4Fria2
NLy7OKTtvUXJrKVRimR83NkG6zAUZOJI5Ootc0NF/y1tOdcx07LyYSo2qDoefcIZ
Uj1NNOnxuUxCU5Gg/m5D3NUyiJaa23eIlGJG5er8kKfo4uu7C41FZyGrY4cCGmjs
t4BmectpshorK5D7ijz4gr5hVWrjcpfDy3D9++wQVEAytDJY3qZnwNBPSE6tKNGx
04/X/jnr4OyatzKCE9H69GxpwbDu72+Rz+IGfbrf9EemhAuXfCYKVtcWkYZEVHbI
0w+Mlv/Ptc1vnV0pgg2+PVsQ4FfcE1OCi4+f0CX0Y/M7QZg52oJFKC+hlSNqtzvX
wi4bdlJwiVpx9De0eiDQ/VNejMU3OopRgEUl6FxMxTw5Jg6/Kwtdel/k+KCDiDmz
zFJO3SGxEQhaSfhWxD5Uh5/RUUM1KgwqHI1vdm4kijHlRppTTOI6yJmrABnTqG3q
IimlXecc4rSIP1ISNMuD7/rdeE6YfzcPY6HXHihNkszblNIf0CaSvKlc7AIvfbxT
AFhqMFHRoYj3fRJN2gqnED3r143oWND4No5I1oqCZ7woOawF5XhzuacJuvgdmyMB
MiYxbck7uGH9YJHCIo3GEAdLGWnb9kWl1JARyyaZ0XuyZH2fEVobJdM9fpT2zlgr
IJUFG4OkvfIhdRy+arn15bWvsML9OFeSZzjwIy7GiNwhMaNyZjk2M7Yv4SdBgjAK
DULBdyrOdXgHtaSufi1S6x8uZ/aSi3W81w2bgPEzemm2ehiKPFAdcxRumAisPJfP
ez+a3NsX2X2MTTkI4pD5TO3kGV6NqBbJvT5SWhg6M9zQm8yYqwbadwfsg2KJCZE3
s8nhLOm3uUvTZSBfD2QOOMsNo47PiMeMGB3W9mCwLxEzXou/iZqMjpPqx7Ap+D0z
9w1c8Lc+X4EsGTUBIJskcQSzr56icC1Ga/ttAGUSS2CsFS0rB0eR++LOBrelMKGH
5gPz+O+NtqNflF3odhDNBaS4tJCCGCNpPmTtwoTSq9sBgmjW8I1jKThA8pHU75fC
IX4i/DYc5yL3rzz++NVJfYygKFeekuroCPYLHPEoZ1cceG3VgD0oeHqnjjIFlYmv
yyecVs+Ap1NeKgAUrdvsEWxeufWlziVdjbRUW+jhRL2e+FXIG4iy19RF0hPQFY7R
ddnlHJP8bLqGNn1jzfPY2tolb9ZZJhxZWRqNWZU0oA0BD48hCuGne5TKZyb3ndfB
dFNYM7yxhlYQ6dUpK6E+1yD+fF0t8OXo6IkzUzk2L2WDMGupuXcYkRp2EeSp3+wA
zPqj20cBQ6tAdilTKbhZaGqMUX5qB4EQVugzevERxl9PmT0qvcdeCwbVCMs0h2YV
68qhxujldZ00mAjUL8PiQn6LfuR1iVYr8Cf0oPc3oLDcybJA/0kZ1c5Q+4/wg4mk
l+qCLLSlP/HTjmJ6oDCAqsb5MbRY+S5kTrp49FRcpmGz37KVeWGWtzZzKmd68KMd
ugC3Rfx7IeJBFH/ASEqp/pXY6gHne5xC5ZV65L8CT+g9TlGnpaAoEGfE/z4mkH/F
RgnjWZd75DrnByn8NTG8H8QEw36wMMA/71jg1fYxFs6+aAI3zgcdpHRM6E81iake
ZSrUEVMpOMb70wM6ij9aEmsxCDycB6ilNkHfxDBFRIKRMNgv/p6DhZuyPzZ2/I41
yPcjVS2kq63apEUsyQqo2ErkIy2zb/CVIS+8dETH9thr/Ph+BRVodWZnj3bP3Iui
/B0KfzCOeYJ6YAnrp2MMLxSk/LSEN+ijJLIao8rdcOkAKuYjMRFDVDapKVXDEMEL
aI7kC2QaVs3MSlWJ/zopgWMBWmg0uyC2N/Tmy7lBH0902FUdBKAMRxeZIHgrseDo
i+Ss80MyFDrjocnNipqy9QAPZRaAPxigB4qgFx8eYGZO2CF1nm2U4cMv6mEbHRgm
sIv86j6+9ZfXrTMdUGsfNwkCs9B4DSTPTaaucMVGylZZBZZBidha26PWMkGo3MgP
ebSe0XeYhXEE5HlJ5fHUJFRwPG3j7BDZhYKK2kEvI/MaBMRAyk1O82Dki4mY1vKg
NQJNqakN0bUUhGrXvlliqPdSHfLrRttiR6JGArO/hWN3AMVPAvbqsZrZMfuGSKzi
l3NJGHLqXKxaIxbB/ItOpyZ733tc7i4CkVGsuvz5nESkbgu3uvSnwYzqSnYAOufS
aeYQuqTbptNpGaUPTbBUlFYjsSdreuDahi7r/8tDAGTHaUETLRGtP9iSkB9hD0sh
zkLm20TApQwtiYi5lrLIH6iHgVN/dT5mr0gCBAe2uLvkYp4lx1cTSCBh2SH5uC0Q
F0z/yp4CdnP+cATfvuwetVzDrIhp7p5eDvMaGsWaKtpyYzJWkhR5uWHru8QZFKTF
dkkp8bqaok0ZK7SiNXUnLxjGmDtc030HClHVynFHeqRVmeGSAalCm8J3Z85BvvIu
JMvF907sEXPKUiGm1Yt+z/a0WD+5nwG8t3y5QxCI70offiwS6qkPwoRJPGbEkBHP
fPMRwpCd4jel4R+s+RvR1+LRDAWivka+50fDjPYoLEiD6DD8ESfi1t6coBV5fZMB
Lti+/nOiUJbU+UkC9XSAWOoIEf8Qbfv+zGQpD1/mrIP1PPDs1/mBmtfHLrVveOPb
7SMSSyY8qb5gJJfoLaTdbBoIErGM+xgxOLq/FGKXxrAtPxHAivx2uMgvB8Z8plSJ
j8ah/y+ws0I4l/X/zoWD8yjS4OkI4lJqn2DUNWWRMVUF9lL5rDvalTTbYIdhMywN
ypaYKb4m2yVIxFpEDBxL//ANgfC/2eZEsMqZW7xSoLqoe0MkAWM+0AAAjYov/J8f
T0s7TF44WfHuZ5tnieSggVf4dHOF3/c6TCaAqfPGN3AlJULnGeZ46wS7/ZBbGw13
GELDFFtzRAfgfTheZ2D0HRf91QqSAemalVaDJ5zqeBV11vbPcJZ3aH7JcZgT+QYD
CrWHQueDxTLhbgBd+P0J/6LFGX/nHIQnPWYWfUfbnqqpmUtnKTbs+Lv4cBcDPX4e
XTaOQ8OSzSWqv28h4vbQdA==
`protect END_PROTECTED
