`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XIyUIG7MsBm9B71hRtuyu12oWA0figp93Hc4iidPtHtJIxsbNkAO98Ei3DGp1L5z
ga3lrsqHRypwEWm9V6Ko8ZujXKoX5YHdJ1bONbbqs7Gr0uhTxwM0w4dt8su0sNC3
mXD3+2H6LOBanCQJmnaWS48oVE1YaMkFu6RD94Q2mKKPHewygs0qjnmNToNbkoE1
VPKh5fLbtMz8hOgHjGvqq7Jhce80c/oxN7kCaOpuiubfyQ393pY/8k5YG+awAQz1
iq1kjru1WU2ZNuh2X0yhG7P48YjbXj7fKw5/1Jc04GEPI0meiSVHF15+jfG8V78f
VL79238ZjDg4GKtKum0tcOOORFKmnJp+rguSYQBwJTdW/AeFZ4Avyt7hrbI6wcD/
119/ASe2tocsL5gL1dbqlII2ijMX8J07uooXN7DqkwoBdRoRjWtTNxsgquLZouOC
S1H2cjPhGFWHlxlSgaxRvCcZ8KMrfrUg3/Mkv+k8KR7MtYGRZydzMN820Tahm4o3
u/z0my3mbGcNXYxK4F6GdtjNXA4y2JyWVGFWLEiDpotzFvoL+giRIzYWbFXoGTCT
a/yaHtkftn9At1c5B8flECc13PcOc93zfTOIHnnZ7Ce78S7fGcI47L5EfL3tNeS+
gQhmPmrIX46XF38ygWgqYFYTBGbRZkH0wt0XWDmEN3DZv/pNJ5/yA5g8uJTqf/nM
3Ttkc5PDExYz6Kp5blA0t94tIp8V3DPlxBSYI49Heq3w7Kg4pqgecS5jJv6UdTBB
eo3rMXfOZJFa6M+tM3m4gjra146oz0YYcc7AWV6rmpnXAg/nYzfoEHxHKsVnMIjh
9h0PC620MTixezLnjxlrZJ3laUqn/smhMfY5JtzplZZ4W6M8aWb81aUVYfeBDzOI
sfyDwfPu7JZv9vR2ilO/lWGnPMuVTxbUKe/d5nHTyyCDGQCsUduYPxmr5O0eiKtm
Qwy0uRiPWOOUw0GhKOAT26Kat1CD7g+Jh3eHXQw1LXT2N79l4+0aXyeckMMtqVDy
dLO3HAeFYEHJguHo/3ywHMD7yzUby9YrQG0K3J73byfIc1YsXJw6qvtPZLp00QMl
R1l1l++dmCLN/NLoj9dc8lNSEe+yYQeKIxxeBcx/dsr0sluS8gJa8PtjVepFByqS
hRy4kJu+jkBQvMLr2CAvj0yF7tHlS1wkb/hoz2AhIz3orC+/uJdtFheQodZUS3z6
R+tR4efLtqTy3UksMi38dHAc92sc8lRXRnXxZkTUp+xha5cT2i0C1j3v5mOFQZZs
C4hu+JDJJ5sq7SVxLVWJkpEuyUpdkS2Kg+td0XlVJPtKwdPSFkEWcXVG+QIC9n2T
lJuJsI23JOx+Mi0xhWH+FwPoFRfZ26QSF5lE1J7g2PT7lnFluk3EfI+lN1N5+NUK
qxycfVTiI50LO6k9QYlMSKbF/ZqQTmRCOqqhlidq0n2OXYcNITom1QxWMe1YPF1c
LDqT2E7y1OTt3qttYHQW318B7v4Gnvtgy1RAjeUKcNPbupOYW4SOgbSCcKWYwRBt
Vge236v/TWveHnqcb3CZ7DzWNaCNj/aJ1cStzHTpKokHBF650Gf96HfrV0GcSqgS
1erj44eLb/hTNZxr0+MG022bburbkUkhGRv132kZ7RFKc36ZnjiKRU/okQjuoR9G
`protect END_PROTECTED
