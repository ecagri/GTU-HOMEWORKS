`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qibOuFn+awwC7jYP6nEeBFglPiD6/VNGM7RvMZT5Ws2SCVr8Q57aRT37yGhcYo2F
2SjKnXMnR4aOtdp4MyO/jmp57Pfuy3KTOly0Zh+74vSnkgHZOwuD1O0JF4rjUuZS
un6aKSNlxmtq0v/hARpFBj03fpPCFRFENjsEi8rvrinjQ5VYgGoC3RCcCk8u7T0I
Nw1rb/edJ4Cbi6qpR7NtsNAoYbok0KKf75YC52FXgllWgFdShSHPFenrgOJh5lMr
wCJVRCODoU+aUzVyKcOi1iGlTzB24Ndct+fyONApjK1+P63WBg/1Nqgy5oKhufaK
42z1kE53hI+58xoZxRRlUYrYbN17NwdKxq7LOYhZ35bbO27iWmnlKtbK2mDz/9lX
0n7O9fH1Mf+l9hPuKDgZrVAlx9vSUrojGXdd5csB503XDymDxWAR3+oKDhXeSjLL
Drdzd6gBTiP/Jt1crOyoCXys5NSnjU9aeK27McIaBosrBVbhM3wEUb8HDCt/P6l/
AHPg3O7iwZELA10/I0rr67T5NeIi7URs+w/zijjviyVXox8Qe8cYF/A9SZbn3bZR
hmaK7c0QtORk5KgRSmE0wFVYqRn7tSPIi9kWYqo87+2Kqbi2+JFP3+7i5L5YPrE+
oKo0XZX6s9mvqAgZ+SdNugamDw0NfXoDJJe+GJzt9cg=
`protect END_PROTECTED
