`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2UyiAeSOqjqmiubX/SKxmn4ewKUJbTRDDH0IwjRPKPIlIJGYLmlEAxQNboGzYnYr
fsAI5jbeh5yNz2MtlxgtyqnD/oIWgubNfNZ2cMz1nf5u8MYD5yd1kdK3VuJ4NMaI
C/bjxdmPtwmpCZk7mcrqrOKTm57RNJ9r79zXAtruHalAVRF5c3mQlpM9D49mjHS6
tuXAv/hyo3wsHb4V6oWXdTBXwD2MHxf5RRsX7me+iEQ1tC/gv0m82tPkzx4cWlph
jWA56KSmC0YdWDsJof4LHVNkSidfPn98ID7Fsi74pJuODfJSQ675kWX6L/WK6Ul9
CrmTE7JAIe3acqkkyj+mjjsWtTcifLqy9limGtkePJebO0tZtdLZH0+dVE/e0zOH
0IZU+urORVWx3B+yHJia/zruFlfz6XLDqZbPWDBy0+iLv6SqNiJeRlYC/s/m78hL
EdiSxmPtNKt5D81tu+y+FLFA1cXM2RSCq8A0KDiPBok9hPD16Mv1RB1DSPg3SHnY
LJK6iNjprstRsDZVgNXNx6/QjIC821YrhuNnNzRnDl69O/aOGq17DLS1Id3ejOrR
7eaC0qYzgMD7LIkBJSwT+AhUCIQYpLLsG1cGZezhQrBFiOT02d8J2s4+lwk5jCLp
Z9h1hsFn116Kj1kQFD3LXY2x4jo4gRnhVBYQqjR8+OnA29hOw6iIsjITnVF1JhWX
tUmK7Zn6dgLnq2n96DFsBQLume7/y9o6u/R7nafGw+q6lal8VR7//eKc622Sl3iV
`protect END_PROTECTED
