`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MW814F9bg4UxCeF9fNIxGZEMBN2WYykpiwV9mV1kLtfcy0IkJ3sz3pUfnl7gK/2t
Ls8j7q6ZyJ7Dm2TVtXsN/B3C2iIqHwv4K5bjSbGlzQqBBn9FPhld9k8u0gmFLraz
OOCUcowzbRmJodjJHc6B6yXMGdT67S8UFKwnv7IUqIj2j7D9Qet6hlrMDwLYF/VN
ategnjYXgvvJ2L1Jzut66QgNfBfhoK6hej3NRMngJ6V6FB68cml3PlAjpJvssaAN
G9kVk/rHfOP2CxoFJEKIRGvSeGSvkSsAXy5/W+HI0CoU/96mMC7uUizFDEPnOx8G
3r+eltYOEwR8+5yGebFQkTIUHhwNHun+FaGNAqiVklet+J2avVppHBVnw4+kVq32
Na6DWqhPzd/MjLQ6Q+K5nspTsDyF51mCDaHXnF72alxqNg8q2bBQXnBUrkID5hyV
LyedJpn2TuykJ8CpXAUzBD6Wok3uC+ClKmBiD5KnVM1RhLaXHgg1gJ0ewKbomUBK
YpYWov+r9Cdsr7EEjkrAcbirT4fHAUd3Pz8A/qbBHUfZ7pKevmOS3uXkGD33LVe4
oH/ihwE0EFatidfn2LwdRL3GnmPHprNg36q9XjN/YnxEjBj9d0Xvmct+sMf0jhw+
hB9CAYCSRfD2WdGJzjOrXcqBKanONszDY6AjSq4G740y6jWU+A5m3i8SKIiddcWq
7SK6YwfBfIPED9sa88bx46W1N7hk2eL7bHoS+fuSJsBVDm2HDc+EXduP8VKwqhEC
TNYVMezqt4XnxC2iqzskixwdCH4Ytbjzy7YBd00AHHcTsYrz20mpGTVgBJ3oPzaS
HAMMjor1hDklQUZ7PFpeabRU5VQuWza1fBQBHrOIs+ZCOkIXXxnX2ZI5YmoeU5b7
FAPC/yF9p3VI8hA4ZaPbBovUUhspchgCioca8f+nZvQRSk0fK2s4Z9XQyhMFVoM4
vwUT6ttvbOrJXRlHCR7/4Rat+NG1VOUbgpaL/H/EIgv5g+kJtS/9Itf9rFiByB1o
UNOmiTHFX6jPVGcJCnNHbnZj/bhvuF4y8jbqhFgQQ3zTY3O0UvEL7//8EdYznXbP
F88YxkuBZJWIlld+NW5pggk2JvU7uNAKfGSF0gfTh0gxpr8xDuZXgzWTWzRibhXd
D9pAR9ZN/YjOmQMwjB3fYhRIEjNTSal1VYVNFOpbSFTh4FUmyAsre/eJvficr/sM
K6v+isCGV2PD/3NcvKvY5HQCkX5B+QMBcN6RVHtRC8fJYv4OoRq9KQnNdse7UHON
0vPjYLF+6KSxMqJKs1hQPlIyoZLc+JPtmW9c4OCv9FRk36i0kkKpMnDRIXZpVVAx
YhTPl6ZP5TojoW4YoqWfYZaDYw19oWA3Kco8G8McfMNoQbEdxiL62qtHkfs+o5qk
JYcvUjb8JWWzMZuXDBkXq6fzBs+cPfhrTgODJbce2z4nw4wMFJ9UQe+jpz7d5BGo
cmcwfg/x9P/vPg9xwjXNfcQqubcbb1g2NB8v+8IVtqJwe9tgxIvxHZEmmTdTmCcw
wpJDazjxN4jmGCZl5SNgTvNmzbQbFJqPRkhI2buN0fozPPjzvciiMw0okmxZpM+4
O89DAA1so4KDvcOmlXKL4WmVogu6Qypg960PtHZq42OJldtVMeC/TbONvRxK8MSj
vZPr68/D6KVL6W7ACH7qE2dOL/Gz/cnZsZmXh3ef1MZLydakWDWn7+9A8lS9jwlr
njECskvNk9R/7XNIQI4Bkm/SmJRt4V6Xz+4PDaLhgWjT4E5gGOAySwBLyjINseDa
gNflbpTu07b3QPJSjgDcafXn2DUqdKHrgk+cIjIxn/rWv/WpKVQnqbtmdYma1X0o
ZS6OLvAcf65U+/PLCVdYlBV3du7VygnVvkIUCzVwr75FFkTHLUG7ld7mQScjQ2CK
WawwUiOlIvFMlibcLjE82l55lGd0n4j1sfQGNQ+nIu5T95T6HYa9HP1gtS0IEcd9
21Q7EfP0gBI45yUv7Lm2CwS59jj6lWREPwv9Yo4q7DcgVMyUbJ8Stz0m1mSyqhqL
v0KvKXpumv0EtGfVjz99Ly1VlrppCZqU2Lk1eqyKxioD2uCkxpkuHmc1NaWWIbsL
EWX1dRRXnkbcZNC6cpahXtYti1E2/GOB4Gkvyj9uDVn3iM5z0dOAbiLuPSt0+3eQ
6huvYKeiog1LgpgDPJDCaDjOuJy0dpzkhqoULGZfLuprbC/ewNu9GOc5r/ue38wM
iyoMLp72EBwteNTNJE4/kEGaJuWgS4w1fPQPesg1cUWdgJs0zvXj1y1aS6TACA7H
C3tVF5oSp/TbzgrjX629+OjbuUUGXnNeRKhnXFv5xZRdmE2HMOYFyUuTPm7MAC9U
GamWKt/vuqfACxiZ8iAQoO2jnDeZpgHVYk3FlD5HlpRj9U3b0+OcNvj/N/hfVjH5
9aWxMHY6Lp7bwr8zpXFOwpZv7zq1bERIMlcszWp9haQNRrCFxStq2k3n3ARbIE9/
iK+q9U3rO44bdzcj+hVAHlepTXst8HcR7OJrjEe77tdTFsVQV22NgZR5rH8ZcBYn
I4VG7iydsP+12HIoXsM9X5FuBUO63XLKMYOiL96fyW6Inq/VsP7UJ2IBN8ubodSw
LFSH1LjlveI46MoarjiILfpAhaxRC2J1YmKe+r0ZFEDBLuD5t1bWQjDUdA2ViZpl
2Hipa91c5+SL7KTCah8eudN2Sz0+UvzI26wldNwhzlYtXJGtLF/7/EWl0w/TozqT
RdtFoR5ZmZQgUHFrOPHaLJ7OyKk5fKHpBDr0h+2X+GPTM9MkbfDtGE079zDT/2SJ
0Yyh1W6+yCWNt5Z1/5Ah5WG1838Nw7c1r24MuU3MzylQd0Zk0PeITsT8f7t5o5kH
DsK9890YlfvbKKooWVmBc7oGYRzr+7Ke4LBiQcVhb66CTn51vtcK7LwRQ1WAG0OP
vXZ2Cy/GbrY+FUmwOQlSM2X6U7s8tWTAi50Z8pwdKKSW2GEqEyuV8zLE3iH393ZZ
Q/lbTlv/WXzQlmP4XqBY6VI/z0Ls6ssp6Gtys5KP2vb6xbuFSBv+5hxp5EBzUmWn
RzgvakdEz+jaFFBNZf/vSA==
`protect END_PROTECTED
