`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fpFTyNOkG7YVZwVAzSu3x2fwGsuFbhiHQn/Lo6AMTsXX9Cpz1w1npN18aKNWBYcv
w+VI3u9Bht6b5gopPtr3gT6T0tsjqV3G05TSLmRGG+uNJUSrIeUaWq9zTci/Drgs
n6RlwXWRa8JGjcyfJnN/Y1SlaaLIzsMsFOH/pmovt0PHaI2kv7d4whV5Rxdyf3Cc
xVoHPkknOzMqRR4DSAYy+hPVENEgchwendGQDsDMzXDUG83X261kPic/ki3lm5KB
cAJbGQ0Nh3BUnkGQeITvlMgM3kDEvz8lTZUyfobjfPrJ6TJKiGodV+iV7rm22VQb
AZhKXMHaWWBn/X1gRnLsvxiUTAjkueI1wBO0bVO8pC8sYC6Lme1pCYSe3yr7PDm3
+63mHnA/k2+su03lQwQz4rT2JqFk9Lv4EhVPrK+R6YtuXJi7buOo83CWWg5zlqDM
MZFPgp/hgTT3WPLrSdfJNX9oLH+4n1k+v1DU1Tx9RmrclV7LpFf/jNZl0b/mlklR
8jngK/Ty8hBG/3FVPmvyBuiTdWMRS890Q5Pi60frgezChUTyAtoa7rq/d7XdiREh
5Q094G5WPVdEKXqrNjA31sB7X9sD4lHpbad8l9/GG8OUPSmXolaZ2kvD5ij3QaAX
gdFZNrbCHs/cEUkaLvnb0uwJNK4RO7dAIXV6jXJnR1GP9WUTkhdh3InIBLQGa4Ho
pToKfh0i+MEoaCitABmM4noXDGUJdxgZ/lHa9Ojx/xF0ySNfIMkQEzO+4SbB2CVk
AdYh3a2xkBbUISeAwYXV3HcR5KGt4y7jlHbejzvQ/RVX/zFPFJAOgqInOJqK/XKB
q/Ky+6FKfjSSr1gGbfgfofFDNqKMJS6n1R1VbDODek5H/rhBgF+bulJ9on27sWoh
vAzfjVyQRLER5D1He3zPtOukzI+8Vy6xYrtXV3WekOqhVyEcpkKV4ZOs5TV57mB9
af5xJ8avnwNmmi6CcFpRoJ7rrAwLNLIBiJsxk0KKtN7iy7tncfrmEOSz7F7WWipR
j5k0uqRJKmEuoVQw+qw3YloEgcaE5Jn+g1blUOWENzb/aCe5/T4SmuHOPU16HQI0
dT9S1QegqgkJ76Hq5dswKMbR0Tv9eNvjwTejZmg06hlwHCUh9oPCl5qgdH9Fwobc
+cBTKgNHJyfRsqpA3eMZUHMAcsFYIFc88u4F7PhpOxRS5SDdxrY6dddvjclqa2Xf
NBkvOsffcujJnSR8TCnP/hDwxIUohismD5grUALbkYS7OqZlzsw1tpXzErIr/yZJ
ytLb5zbHwqQ7CzHSniXEpdTOv/4+pmia0FP+wwCboIw3cdKqm0u/ntGLsvTshsLt
fQkUqkmKK+RPBKqJM2ebBUluC/AxGug+XcvcL8Gyok1OqORPKD0uJUlwTbQxObo6
E8xoKVuCrwrwIPsFMSPahPFuRsKXEmFNZXZgBPTBcOmccoGnXFRGC2j1UZbZ+t2t
a+8/B+IODgGB6Is2PAOZh48fIIBNiwTp1UwcO2+AB0xMk6KSVO7AkJONqGCQLDvh
w5FHg3GWmR2e4GMHsNvQnpNRx3E1EPi5EVRdFRvKFfAc/FctzxbW4qaxIuk4MWAi
GQK/6cvKPUBc2hab744hCFaFul534/tyIPKKBE7z724kkY0ohwv04id9OzF+bBAB
Taqw7qCm+sMsr4Om85UTjR5zKdtslJUHtAatP9WBz0Zy1Otwe6qfAhZRteEepS4G
2gsWs2Dq96S1VXx+sXGzHmxQ1K654VpNxMpYDNPuMbsR/eTY+hmFHBVbIij6nvVp
jD3m2L83ejz8YJMhp1CzdttOTo9s2ycYh7fpQ9nsLxyhhMfYJreH+hsHtDcYf23L
1YQZSSr8w3M9mkidlh6QDxaJp8N8yHERXJQhS6UpexSVJBbfewY0roXMENQXW13r
33SSHZNEZTUh+i/+Y9UzFwiRaMDGwpagYInqy18KJjAm3j6tV8VKwOupVwt5CGoo
dPTzYNUbdJ92S27mzHvlZ7qE5RfNM+PLEXIp6cB/W6DNegS2GqjkMU6K/qzZ9WDG
twPiouvBN/wNAZ7DRcVq/slmTIatgxBQZBBrfY1ZK+4fUS809sTvVs5OqmhPnIIf
5iTDEQ4yGdKcQqM8ojvbeOzPlhdBpi8iiwtjl7Fbv3Np8Xgmdc6rC5JDIpRX1QpO
/oL6hdgojlrGfeoLnIfYZQ9smqk3Z3Hw2ZGCf4ZNhD2yenKGS4Y8PMdsfE3Auww9
cL1FY2oe9s0GLjwzbYv2rrDDMutjJcWVn15zH+q7TfMBuvX39sVRx5M2guPCUelC
bSezChTFi17BQ8kA1yesnEBeBgQG2cyZE+vRcjrWp3uo5Y183zHkl66BLQSsvFKs
fpnE3CQ8UzTuq6yByQW+3KOSokAKPK8c3HFSotUGBS67l2jPTW5cTJey+xyn1dUc
xhAv3NvC+vqBC1HJnPa9E7qrYZsfvsatyuDkISmiRPeFQGRd6ywbq3QsH1LucihR
MJ/nqz9TMbGhxjT5m/ktfwcxjlsJC7didet60dIVZmwqHIwasysI7hqvJ020czdN
e374Qq6pSIarsrT9hDo13FxAdUGdrfg/2tQqHSnsFQTMvVDOxyriliRAY6yzkYAe
kNaykdilXqKZ9/EPdSfqlUBn0dVRrEZ0xkglcl9V8s1IhQUePnEPaYqwRGoG1qER
JxsMOHsb1+XOjchu1vctIyOaHB0BwCjmAwX+blgGLKZVrPS0arKORjojw20KoNMu
VbxiG+S35k7qju+cSclmi5/+UIHqLJFpCjE3hlO1FR1G6nY3HmsNCWyyzXqN/OsW
LCAAi5e7tDYxoWLXzMuxBixD3nsdFLl2fAtZeaXD+xUMw1fYSlVgfSp2w2rFWj5P
6tuOe39OtwLW2oaekBABHFofAp/RY1MbHylKFtpJQjHrT0JTrFijwllmKrr5IQie
mjBb8XoKZDmcTONcx0JCsi2V5bCPEr84+9SClVc/M8oUKm6t3DNBG/KZSvYqPGXh
Wx4cAdAVH5kftPUXU7KeBpO3BLrHsYCPJd/4xyEZe9uTZHSg6RHxPeCYPJEz4gl+
ocDbc+BT+6693Icm+yYb8dtdX5yp96QOCRJvtSVkOovL8XhZGAybV5M86qS7g4p/
jFAUmcDyIf8Zj23BMYl5zrHrgPs9RnIos7qx4PLJmUjR+eYy6c1kRNbaxJPQayqj
4QbsVxkOaKb24R8/3xAxd9s0QEhDp2KMpxCSY0hvE5QMW7oZNCCVuZItOMrZmwYA
uVT3tJ9mBe3xxw6aQM9I8NK5Ampd18vwTf38q5wHBs1E1NkVhpo2tklR+7s9VLA5
xBccKUiWSdxouhYy5Klvbw5CJ/zmT1WgahEPOrfSbvw=
`protect END_PROTECTED
