`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kWgP0Raj9pNFiffuYmSeQ4+V333ShafdEWHdES0YIhfcraT2PAkXWXMudqrfNtNo
MaGdw7NxAUAjPnQcBH3P7TYHbj2cTs1tJD99J8646a3J3dcCdsAe8EBMktM4EnKI
LbyUCNXBR9gEeJ6ZBHgJ2AkWAzAavabXaiRrEDi7tP/cz1jNg26BP9kwpm6uSSye
wuUxiVEO2PQg7mBIoMIJ3EcdOGhV+YWFYc58OJsSUmbRYYyrzE/y9JzneWPyGWgB
rdzOZtVtgsAEk70bLwD2/jkWwNW+AxfqY8Hb8BHyHmqCl0V0BrBoWqEjH0ticMro
f/UOrJn8Q51ncLNlMBdRbYX2VWpIKp4XbwjPAi7E596sjMqg+itPcrbKI+QMKAZw
CmhcmHYgnADD8vYkXJYYVyCjIaRHKB1g0XPY8VI1iYjAuLsoDkr73W+vZVOUY6cz
plk3eLQ9QaMh6o6g3C952mLea3bbS2T5fIaSLjrSfZBf1Xh8k0SWAu2by8Y7UWBd
Qng8cqt76KCbKCyFUBlTzLBAWV1gaAB2CrtV1SAmu1N8c9oS1H8UQb2TP6N1CyTm
5OwMtRd21XodkfXQtJESalAdLUlSgnc+Sgw3EXEY5GIsTVhTk5tSaRJyV1EF4PeA
fq49Cpi4IHQkdIdaUmukhOdMu6NJYBffHxhg6/1MkpwmdWlWCPhGSS/6OQHAgY0N
szGkLkAteuMgfkmF8HdsKJpeLdDHqdv6JcGBKo/LDbHR7dvQkrQUrnw06jF32Y4u
Rr7AKSCctyBJJ1zvZvXLx1HeZb0ZF7TwRtc/nxfoC/MBOEuiPSNFq/tOYjymtaKu
SGr4SSyDCY7YuySleTgQDCmV7dlWCvmqEIuNLQAQ+gTbN3BKpcEZNt7TaUqKaKry
PBFoiEvgnS9U90/CMYt5oW2IHdrYV5AxiJZCKw4D3OHHmabymD3GGLZzGWvAPTyU
e2Eki8tdHq7nnbiJnqM/EEKOnoYOhCLvRkl8svJWv86CiNrdT3aqbD0WCja5E8e5
PK+GR3gb3Pb5Xuk1jGkvx+H3zX9Sv5Jnq8fPa2UvJGYVbpKnEC4DSl57MomI7d4l
7rsX6X6VBR+9WepgLs5k1kF0fbpbGGa+gZcuKPbgfn5PY94DgwmzRfq7jYgMpGlP
UwV3JRHS7HRNx3HNWt8cmclHBL/JtF481ZeOwHKL9FvlwsXLimctcEC0kWr9bjKt
bCleImfm8e23ZAOCEkuAh4Dt/aN7O40TserLUUJVVgUnvAxWmunI6VaCbfhAFM6e
7f1co+aRszQdhBBOaRydxM5CdS/uj6YPRedlUneyBInwhcjosgeAorrTTL+e1pCV
3zVEgbb7IuZ5ez49SndYLLIWwAgoyMXIqP7MXrOBb9++3oEs7az08nrW5iMryDAH
beUMdsd5mvxU0NhbJ46M+YvmZjptC2vJR7KZxNDkTZOJ/KK0uq94t826Qvj8n76q
yTv27kSx8Yni5kndRCQMGswslGybrZm7Ih6r1BDo+BQatw957tOy3M6qAJywcoQg
r4TzmF/Ni5/oGPVHy1nzUHjWGFQ9XOowpOFSNu8V4fHEbGjz9l6PlBoKg/X5GfQW
ipgLFPSRTuDz3q/1gR882NRQ7YXb570Drl62dhm17255imVtqoCtk1sNemy94/d7
WSvwTlLHxkdnLvFTdebmEzCaj/CoOq2xOP5L80AedDn28JaWzPKJXPAkgvdnBRe2
gYxMgyfP3lcZHRdYzCt9zGsEXKDPCD4ngQN8wTcELSZCMVNXqgwic6tLuRVnTM6h
B8jStq5Q0rLk+l8CZTIwdBfh/7+lwTAl5HQJvX0TGg8F29NhWwDu71oXIro8hhVl
DOjreTaII0SzBVTSVXZvD+pyWXjm6pJ68oPyceso4R/U2i/Uu1LLv/qJKsbQq2mg
H4YHxZ4FaHqZX6qnPzDvwy+CfoNSV4wMQS12uJbW8/qqcFc5SyZ8h3vejF+N5YSb
b/2Kce8bLFcECiboamlJtYYPIX3RMkU3YFp6zIlU4Yx0gmFqV3GmvpYY4ef3fdCY
SXojBUqDn+Kyu12AtiMEX+MQw5hjmaM/tuL8nQrPCJjB1AYF95zadALxGx3yycdt
JlXHqwyVQe8nyPn/gkdlmWu0s3MS+C1aJCVD3+OrxadBbax59664sNuVeq6epSZu
9TvAzrz4Kw48cyTLpG9OFfwwCw6KXYc3FRye2PL29O4ITW5FzqCSD11V5AhEANtS
4JgQQvxYWpk/8hMDjcfZ1xpsSShK62y+WCoJApj03lhb0emW+tITofr6NyVG1qc8
e7KvHmnwU/WV5JfPtlQmAhtue3SQEOCMQ7WofxK63xBRNcAvTVZ9VO6WXv4+9Nuf
LGX+ltPOsBi4n0l3Nq/bYNYaHfUUnsUof+4hpT8XiG4pht3RXBt4AkGxni9Mbl0Q
A6DoJP/u6QD9ArZD1JezfkmOqMGgjsqT8YVb1ZSfr6KdDjwcpyy26XDHmHMXU+Mx
YGYRQUdQjEqvVFY1wW1K/7yCgvsXRZazTlgF7HTL98jrT9tcY1fyVrruJLQ+2nWk
XGLUQQXrpn9jU4QJCk4AZqybte2wi1rG+AriA27IjTd76hJdyoOQkh9+zlcpJS3r
GdOAy5DuxI+iJPBbDEepSY1XqW0U6pJpDyp8QF5Q8lfURBpRYt16q034Cz89SWnu
IxrpiT3qi6dEX+65ndFSMJ+PJkdINWevIBlGrhpQ5Hr6Hcr1N6zZKqu6ldklFT4A
YnIuml/gon8VqOzqR69fKTMgpCPkmLRnPEXFqEUI2dEY9BSbd4cNixZxbqaWOxBr
DeQPU1hfBiBB5hJb85vua4aqENnEy0/Go7Hq8aZM3nzkGfXxrqByxGyOB8xYGeI+
RcIrrUn2bQfJO54RACcB9sxz8o1MLDRTpCtEkxyskyTQA2z7P3TRptugPeyfkV0t
BYhB9tiIKugqrXodMy9306rtjrr3Q4UtGzPEDouxW5SEDnTN6PD68vmnb9eQWy/W
+2eo2HevWFiaF3ZBHjO8Dzmj4EsVqYDlp2hDQ//kXtrKxFzhBFdOu9K+XqhcHc6e
RkmqLzgVYHHXSEBsPmcqU74EF03kZ9EVf3DUypMjnKK5ThDkzTkrzAZ05O5hu8Z/
sCnb4tuwllKHHUzpK4ZyHlvK9JawNlwtAjxvpS5DR9tWHQNo5tB00Ai8DSE1PAnK
rW+r78X/JDtr5A6sxM4yMVSAimGyfMI3IoGC7B8g5L/7+Bx39wi5hbdmzkK3DE+Q
kWneTJ9eBhpvzhMU/SGrFk7E76jyDAdCyNeVCJe6oIf0+XvSk+f64ZX0xfKvgA0+
9UbSUOXEkkS3GSgwnCPim/jWH2U4ip1F5td3GzztfJHhAr6mqU/q2SN6RgRPZ9Md
CMO3sfDNEa1Np5zoZ5/7j8py50FPw3uCy0hJUugr3yrQLuH6mQDHc+9tcY6sqAR4
ZjfZk3zwHve0Ub3Ac7egHIriexl+w0qrPnNG/hTXhFvlsbcRqpBuXSABwTxlK6/2
z/vp/kRT+TTFbWioLgaGJD2KruFZD6QIh99gumUHu7WJbCT82HYgxzEV5wgB/k5o
nzs6om5uXGEku/TkLUafy3yRKnJR8bTLlfYAfYqzcFoahYrG+1ibfjksk9oKZYCc
lNBZgAlxwvkz91++pDCsb3+dUeE5PP4DdRGzlTmx3fxwca14La7XCe+wZjvl3xKa
Z+2gBeWu6zKJ623+g/oIEyk7mOZzB2nxuHb0zhBI4NqAk7tY5kacJhXg1ZvNy+1g
hH8EE+1WLWiyPSUozK9J/CgP/xzKkVOoidmcDK0Y4iRVDRzzcXn8JeHYyEQnW1PN
EAplVdIycLwDETxc6apNA+Abd/nIm/a2ttMoofFvDLaQ32QCywER10/Y7b3vrEL4
HTSbs4weI7xLDsyEI4TtqK+s2tTKlOQjdGFKy0EJ2yKRaSZtsP2wWtggvkfiXqZS
V6413EwJSAgcz3kbkPHnVD9GHb6YoiMwnon/yy0EDDuk51cBuGlhGTABcHrvB/gQ
1M02Z4bspkEbizDyzSJgasTHEcsJGVog7P19wUeyfR02UKTTeUUQUxVRn9v7wY2g
M0/Ez1QCyH7iyeEBj56TcHoQW1ZyA1DsD5m3lYMGhWWP4b291XtKj35XC4C9Kqcv
xCd806mgXIAbn7pgL31csgU7ix4T1+qdyqrLEIOK/dxDGcZjcNNCMvUYlKM9mu4A
efz4bA2M7lFRgoWcFPViWAUODbkdMEEnRG/b8dngi5WXoMwfx5hg9olr8lZ4kGe7
fe1ToDQ5LK8YT/pgeGgm3M+QV+udRrZ8nf2UEKTwnovWAnRSnDuwa3DRsV3cMVAF
VTew8zX4HDucajpGzzaHdmVgTFrzwozMNgmICrkNw+zXeJj271hRLPRgr0kVTkQv
wW4fbBvQFWJ7r3jNvD2mRdz9T6fnGRpdpoPi44k8G0mrmE1CHeZcJh45svgAjmBu
hJV3z87ngjPwIgDEZxbQVY92BEwhDA9Ov3udBJZhnsWIQxO3eGk9oatuTN3M0vDP
suZKszkzsoI323AgY92IfcuFqXK+fO8ta4eZ2D27qyhxoJ2LJYvohhCiVW9nxNrN
Hstb7iv4y7heWKzBzjLyxiRmUfWOibnlUYCW0mzz6G+ZIVvIobuzIgUI3CW6M3kB
I2RHgHfOgVxRfMe37CEft7FVxM93QE9BX4foM4/ONGsZIcWZq46qPgAzXqBJZZat
9keP5Mq+zYPVSSIYJ00jVdvx+23KWh8bVoAHTFgZk4Ml135pRv4q1Gy6DBQqnzv5
UNsu3i25vbyZM3KmRfsCqtLs/j6xaxyaIfP+Hkyton8bhg5Wsl8drxJJXZnPt8sB
nHXpe9RvrF9buXSKtjxqZk6uc7zjIuRY1NBvVn8LXuGH7MTBOXjjIk4qEvwR87gy
TYWyOYeg+EBd6fTdydOqZbJwRuzMQIIx2k096nu7ptHfnlc3fS+REPLFz4jeLHTm
O4QunBVQYvvqm/1BTxQyA6VP504zRErLZbr/FGPUuj3aER5ALaWGBNV7NvjPj6no
FsXeYkI1tmWJ3U5XQ1Ed7ODd7mLFC6yHNOX7/BAHyHBnisrV+wUWFTH+l1WkGpRv
aM6uyn5L/CUrXMafkmq+9X2MRc5JViCi81YlVk2hZ9pkrmQ7pN4hXH2YXxAJR100
YKyPLhDrcUdPftR7O1/Opli6hd0TPhqjEdSo0le1K8rrAlLG98V4DHxq2xWDv7/X
brTatUp1IYIAYDhq8+qT4MKbPtkKdLtFHGq389C9mK5Y0py8SPkj8/PyrObsYrE/
ZosWlOCBxbMPICzxpe//gO+S6yRCf63s1JDKNeBGyGbej7rLOJmLZAbVCOMuWPiY
jLSNv13O+I3G9XXrsy0AdD/bxX4d3g6rqQaH5mARrFCcV9AKgG6XOWPEx3QjJ+7I
i49vCYfbLYkeJaeVSTYxV/wlweExYFe1L8tFx0zPasVwjpe2El42RT303IxNNkjn
ABGKE5XDc69YldTUJ8Euq8IJszn7S8wUfutxs9C8sIJUmxpOqQB6IYV7Ci6jBfoT
0mzOJXMHyxoAIPCoF5sJyhrkmz8K5PtrNVHxmdkFTrxUxvAAEpA0hLOwk73uC0+o
5ZJjoBU54j85BqibRxNDM0o2doVd7WoXwosrfmt/6eX/kG617FzhlfWK+68nfyn1
Oz20LpXaeuZzWUnfnrq99vP24Kc+Rim3LOXikJmTEzT0fyCbht8S0p58XYkBtikK
vq+YuXtuFGiSIBKCZRXFAUeklSlQ52wjV/aWllBmn0oOQWhf81nCeRNliJiokkyS
+K7tA6hbgrU/Y4NMYViqe8uhr4VJGFgnWcpfd1UCNnqRcLQkRUnd+R5IIBVYLLvL
fHITFG8cQsVSh+v6U97uFfr0abSIdp0bAuIdwU3diLammutoiR/tLG5u1dzlZ7d1
6lHSEkMT3R/hDiQCnA9Q9OqqfmMaP09SG4VpDEZMjebMM2S+JFS00RmXpTncDKva
skIICXyboNUMU/Oa8qgEPXVvYxGJ2nkvpk+veDWvA4ufUZaLQHvcizycIrPWZW/p
MdrA+kUkucLER8zkosakIqRjbNRO8D0xkklbWCX9ZgGVoGMQOFpS33czReDxT/ac
ynJzUXdD2nPbQfe0C207jmAXVekFC22atrJGNh6d9ymnJtFrQM2Cmnlqv5pJ6KJR
J3aKTTqQqcIict6UDSRFVNzdaoaNZf+2/JFTxD074Wg9VC7eQYrV9fyLsCn5nHOg
3wiL1VL9PWRQlp5HqPhf5q01cxr9L1oICyI3e0DgbDALCIL18T+ZwqBiQGWJyM37
ITg/vF6eJdSws5bFyz1gd0DbBPTyM1/bGFy05j0GCaHF45zEWrZhAfGYse2vHLE9
DxvsUOBKuZz2W48esiBtRjrWDbVVFSyrln1MBLm+nT9yMcfQ9F2ZwHskWpiaf2lX
I+a4BryvDgqKWz6Kbz8RSugIe3zAGsB1tf3Q4xOpWVgzp10+Roz2idUxlJwzc31L
pPYS9YKft10yduxaW/UWR25zY/SwuHupwk7/ZrP5v1X2BuJFw7gkNKtIxX6HxK79
iIUXrVAltZY4qP3LWwfOCKt3s45TUgoFlxfZo99b8pEv7mzkABk0w7h/qyfbOM+g
24yKh5hjbdvINEt53a/c8uYalNVhK79cmTsCGS91g3xQjCVHGwCkKDVO6OKrRiXg
5OXKEObAGmaGxN3DsHBEadd71GP9D8jYRJ8MybAvgFg/G6jcWzO+sRDFN2U/PHoN
19/NF0CIYnVovOT9IKjOSwSN89yj14xDODocAQVfXATYq3iVkzPAzXNUsZRv8p9P
XQkll1T+M3sJ5gWHsAfQCCK424IPAtpHjAyRPyAvm1l+TPTk5lkkzk2zMD8tBXmM
40zBOE51okDQr4EWqk4cjFNmWheBCZ0Bjy1n4G6mD1p5t0Ja04DPvVjZljAdAwBn
Mbz54ocnTqkKEL6oYYsR/jTaC7EAxYLMx4V89gwBxmkmUXnISLsckVixOD9ya4Hf
rwZL5H0Tq+IqW/quWhjJjunQDN7Q/LMRmlILUOykZFcbzLkc/Zs1sGUSaYUNfrMn
/5Wn4eEgf2KDxq1YMUW/nFEyunLQtg368FktFENJSer5bcZrr1jwlVz4nkQ1kuf7
aASBcBw5Xc/7H2nZJD+TKG/LhsWb/xzstjDh3El0KnHSq179zacJ7XOZH2vQ4vy4
3w9b9iK14X0zJAhDM8Stku0KYBnzfcBj7UmvUnVbNAUdMJ7oQfxhOtJOkBz7NJXA
CKHBAtw8aVyRqCzC/f5cswPdA+DcKgMNno/vHb+0yI4SzDwCp3DNyi7gfkpNy3hG
o8Rs6QC+PPd8tokAcRmCG/iSDBQZiO1zQabINFL3kc6FIbXel1jLSiuipVZyRe8G
iAKQ1/+4LsWdUparVZ2iikU7YmwWxOb7W3PIrJDv0qsGUz17K3Q98yC/47vZ2iGn
mGDgz+dYFlBCPt+CnLRe285lIgeon3s7Mg52nxdvUu8HKaVTGzc/4nWMJqU/Vkyt
UaX0dsXhjagLDrFFrVx0oM4UPTOT+UOnLIcBdsHGDL3vfLXzXplLmiF+sl+oKf3h
oelG/SKSW2Shp1/n6rK8KcxYr9EHzfZxss6n3meFeVVn772VaPA+FAogEVjIve/Q
0m7JPnfut6v6Mg/NTLdiWrY96o9O0T3hpGD2zHWjNr8IXLwG2IKEKj+zmnlrisaw
Ldo9bDkA9WrZ7FUipsn7kg/8wAhnX2zSU/kWcivyS9QPMWKisQPwDqR/N20LPsSI
jcKnO6ZKVRgQ7AVP0jtEK+G718FQi3yy67/XoizBKJGfYajqGfG2q89Xplko9IPh
6FEbPl1lutLuprs8H+zHJamtxAB+oDjdZ9+UJf90s5UjoWgzRPsoRp+18uPBqCw7
glqdoY4cDUkgWFfaXIFNgzljPGwWxLMPu9/3A1pQlfW9vboNNsMk7eRk/fD2rrIG
/b+/2qDW6Rv/Stl81rfvM4OiauUARbPHzLz+pFFNxsTqQYdlUe9cPB/UI7lO52y1
ygq+HvZlHBZPAUNYMfb+yXfWnQh/um+i+m784BQR/jRBqDFxKM4iwOLbFtyVpp25
/8wzP6QtYjbh2lImTciwUEkeuUGVduSVefpt+SULXstCW0noh5J1Pt/TyJvgWyK5
zQS/BqNZRxVCShqVFdoY5yp2AGnyv8C1rvhPiTfyF3OTzu8QXVkicuZKi9kuXgQK
UrmLGbL1vpCa4qsPlX4hF3RvAk04TfbZ5Q4H5FkLQiWd+CfpwYXAy1sx52NrHRHD
yetpzxpvZ9WQdLXUKsDi8pfrCfQCNxcQ5T4/pwD5556vFcwTda+fERZQtnybdMQy
MP8+hbGAqQPDTJlmRhfCcYIccR8wTHtESkbY0OgjMXqBBVWQLVQjB0k5eP/jU/KX
KDfSSHtS47roaQckNQk9q4ZJQl25pOUjvim6ZSoIrAmPQiNtE3ya9kfouSnv2MVr
f5Tea5Cv9iRDu1jycgcsEoCXS4umcETmy/WJePmh0XnLa3LhFf3RLyAQkVTP+J2Y
Dkv6bs0Csr9Y/0whk3U2T9XoyK9jxpJHJl3iR5qtMMAhEA+gDAwkKFK4cpUnVPtC
G/EmpekB1JtVrJbNgW7xOP1+mEZhN9hFWyAv/mh5DHuSMgGgorxQwG0c6S3pwIVA
jgpR/CjQdtBIKU9F+Qznp8eNxnRGv4TntHLlgWp22yYNT1TvSnqyuiBD1ea07tt7
FSdkE/RnWCm60RbG42GpivtAnODSpWBs03eKHJcBMQ/zPvGCSysADo3L2bgAcOGH
yGHTOHUl1dfij2nmofDc6W1DF1oTLWcbPM/DFpp3v/Gr21TdECKfidajrz0CUwqK
32zhp/YZic8jQ/QwkwhJGY8USNvMLwrtQteHX5fyRvczXEVCaF2j6YumOhmqUCKQ
dyN9xlwi4y42mt2SNQ/7WI4i9pSkWNZ0phDX1masHHMGo61Wx7Q14SfbkxfNDevO
zPnFouBrMruFH2vfZYAK4R114HG2oeVIc2Dhd0h+PeCe0kosjBsu4H34KRPoeDXm
+IM1PyifmjmRQC0aGIg+c+OOuJUvoSqCufaTFRoAvVKetZnE7Ld+NVUDBoWSkRHM
CjR0zNM5SIlb2CR0k7dWfhdUi+R2oAL7FR67b001JFGkjKSlsTCg8iHuALBtp9ot
sq1LziU7iy8TXyLt+tYFVx2QIyIkz06FCqUtbQofpZ47LnfVHXHJ3ZR0MrdGTRu+
i5qDJzjJfITDXLGfdvTSZmqwBJMYyCLBYvukhfojNF4tb2baYel8BFbkTxkyCesO
zgCSPXt0C01pv47lpnYRnciqKiXbNl/bcHJwOuWzsm7PcAIEm23iApWTKbbAR9Da
jMLWEJ+uYbvDhBVLcpciVPQcDnteNPKoDt/JshgPca4ZqwTgTt0TOaNFw4MmnPPe
kCO4jSFY9ouoK9ECko+GIKHFYZ4hV/AwyiT1SEJLBK5kblmjEPieaL1gjuLdzSJO
CIbsRKTiNdgclqDa+Ghe/EevAeBPdDfktOR0JnT+0t1CytRNrD4/7OdQAukLwF2B
efjfIK7zqxz/Z1jmFj/7tv+SXgdAuPSsDCHdltDSTTZFnRquJ6dNJrIw/h1UvwC9
FfvoyJJuSOmDCJU9+x2YAPEVKGhSvhPXeTOQXu4WXEozoWnELPTDVCbYoKarSCO1
`protect END_PROTECTED
