`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xZw6Xls9ZEYj8AVlM+i2ZEyzEWR2EqH/+oTe8KAstay3MF3B+/rq5cYwQ6idgLUD
/AnZlf6DsSlYQhwxZga4xHfkcYSvl3pn2UEXQIoan7h91PjkH0xrWPv4w8ksYaGk
YM8iJApIWhgHJg2jFOS80nw03TvTIM+j51HZhUvxDSFHqKwdOkd4lZrPBYCX290u
BFHnoqMXh9mxNfaWGbfXCArIA3vBSa4I+uEiRLnus0XltFDOXB/fRM1E/55lvMS8
WS/pZJA7B1Nf1wplTReqaVfIaD3uK7gDOtnYcr2hHymiuDiYA8SUF5sZjCRjN4bN
jAvfIkdsg/OiPgLxgcgAEQ/42Wk2T1NNWkHqMMo5fqnkifvTJATH4r2uOvSde9gW
RzEUqcvoRDeoPjOaPmIjDA+D09v4QrhXT4CgexnzdURel9FMnGZhyIXIazAtXbsV
D6FIBAU8NBj+waV4hQHBphVdFjWTWPDUF1W3E49L1Ik/yh1CPqB1ayFu4sKIeU2Y
USyVwRYZlh/fdQdQlVCb9QBM+PrDgbvuYlZFpr0lmdMnX5jEza+s7QrKHFzI41vO
y6Fe1EbRlZB9S4MFZibhRL4xPsJbXb3WlvhN5ky6dX5gjXQZrBeHH8HFlZOe+CCm
5nwdecWKQnsmUR3vguZGAA==
`protect END_PROTECTED
