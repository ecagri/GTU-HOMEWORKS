`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bpZKzCtLngtnAXhSqZuvEaVKK74Nz9xlt+JCXjyXXFXsRiuWbxHRWaDidJWJq6VY
kdrM88Xkx6cypyNgcAM6WgdgOv9yF0IgnUNakAoXtsKhfqZ3qvI23uad69O9Sedc
5VcjlGwo7GVaXjzzuKGh5HrlJmBynB7TMs0jC6togtDQA/8P4HASwYI6q4330ZYE
ibKsr5u2ZT6UvV9N023Fm3YIn0AMDOeO6mcem6T7Iy5RGg9u1bIHdVJ/6IXiw2I+
y0/UUz6VyraWPPHK6w00Qi5rQy7Gvai1TGMYDFjgrwfy/gbuenkXbKRbOVC/d1rC
o/ZPhRi+4IxK76JW1H0w5+hGNWP8JQC2HyI5lem+TK2ILex0BrDtGv+Rb4f/pLzE
UEumKK2Dtjo5bQyG1ilW4l0yjTUfKVa2+m896Q9tsTSTp+wzJlqMsfvMvoFZ2e/I
o7+ZeIiumT+c7R/4fJO3r7DUTU3F28JgZ5vyCKjbX262fUIRswXoxvhp6KYQejNP
GpFzEmOdOKDfROs61x2iSvrclGcMd9wmaM0P+WLSRksneT1ZZNagccJv62KIzaYF
Sl3N+bwL0WalZRYe1VdohNQnFZMOfHLOZIbuaj3mUHWrbej9082PQtmNKdBASpI1
RaY4OOqhXSD6+SiEXqKwzyPe3MdF6RlVFNAyXxmI5LuVhGspDZwhmxu+uyDUBaFb
JmE9xduRkXzBpaNvOqQxXPsSZTNhZQFpJuhE5bTwuMTd6W9whY+s7pliiFqrUNBJ
N26ZeG6lnj4vhM/aqKK8v2uU0I3mkusBJVWYlQGbYbM=
`protect END_PROTECTED
