`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1BdScWTnVzY4dhFOzzw/8fVGO2m48T7dEEwo1nrgODYgyku61WqZ/b/wXOfBjNCO
pGOM+ShSWZV7cFkf/zPcZiudM6vgPlwYn18SgJtTaBgPxk+3BYXI+NSPhck/SSP0
bu9f2HMtm1TJVq9PVv8mmTHt64zrJ/GkE/wKAQduD5rGK5MzMvOFHwVkO2AtjlNi
xMgfuUIiZFnysvOJO13NU73okZ3+WPwye8nqZhWnUyUoXozuqGXUId/0mnRd2Eiy
p4CZ6Q4AHDGIzZnfba5u1FFfO9aOaqF/HhaUuwqxvQDkXZl5JKiUm2FXGwADmzOi
ZQ/w9W21ByliJVKJo5XeposuoIZIPyxBGbocVuaz2Tsq4QMnrGzQDKmjDFB5x9CH
VjqqOlLg/yQag6rkZGjSjTdCVM9JN/WLSdpFGrZe64q8hs+g8gkOii+iu5nxWRUp
r1LLfIlbSzSaaJuztcHYKzmZ5M09n5kv61FPjS2JzeICJJeMmMWvCK1vLcBR18C1
xxSYxcm2g6owqKPBtSn8OccF0xTFqfM64X+pajIc+WwOuuWeEMMCwt3JuMUE+evg
5zqpjNV+RKMfpuHL7srf1eJymIMYZ5zWCDs4wG0GpkXhi0HtDz8/L/AQRMo7MFsx
+xUi/7b9/2t1+s9P9/80Dh62FNFeSftNb5aJhu2N70QKFFJxDwfEOYv9V/aP2AJX
VcTRlT4ARmwv9F9xmmcdmrYDjZQO9q4bVKW8zHvn++Rm6QgvLu74dGZaOa7NkCHP
awN12rA9Zzy2HH3owHkXh8BP2P/bcQRW57nEfcJm1gInUgiVytNntKf4LlccFMeq
PmqwkADJ4uWvsvXqWL1SZ+dl4DGR5SMhChnMr9UxtlQk4ZE/P5/GfdRAgrng9oBn
IIVU1p/4z0z7C5Sas4YtR+n1724nH97uKnUh/LAxbcBPFRXFeI/Q+A1YwDCwy7Qd
q5Fh1jImyEKBABbptSwoUNB5IeL0bFLXHkxPFVD0t16ldULFBj87s6sAVXC3o6TP
zLgLekPWIcnN10GfV+kw17KOC6LDhe2RGLjvX/WxHK64pXGYZGlPXysl59rKV0XG
DjA4P0e7SMe6SlzMWQCodCFE/hljop+1e7+pyONbDQnnoOIWEUMs0N/f4soz1vQ/
`protect END_PROTECTED
