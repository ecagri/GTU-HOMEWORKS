`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zmTeaSj4iISZIEvuSZl2x/Xam4VNYEwt1BkzrIwQAC0ZMcdnccSbM0Dfr7qMO3So
4vBafMJJa1SR1I8yJAdeIb4VwPwxC6pMhHPo1kDOIKFVSXGbBAP+hHD4ooFesKcW
50uDSq0QBXUai8PoGolPIQ9UhoFce0a6/W2w0tTA2IZJ4o+39jutK4t2Y7SizAGY
89xlz5cmdC+gIH2dY1hfK5ucKZjGai96g32mYNtp9MJueloPhs4Y+7PI5CjQ56Di
I0uVk50vHAP5Y4UdBEZsETJp814su35IlIjq8/ETk2rFhtH+nyzZBdNsC/E+1ACi
MHQ9tx9611Yq1RAdJUzH1HR5B7ub6DG+/PvjZ6UYtpvOAyhPK9vjoRh/Lh8LLdLs
fSPQtA2yvc78sYDDP0eGOOq5ZQo4aBxkhoTU0ds82Yl9x0SyywLHOfpiPfCUFoJu
L8VTIWthDLzW5a98J1xMplZRfritWDDpe077sI40dOIFbZ52BbowON5najirI0i1
zqJO6k0mPbZf1NzZB9htm5zMR/42fWf9AwqazP3MhFxSD6uuhmyuoTpXke7qb5Fo
ewwYxYm+aNE/6U3CtlzRQY06zHX4TQxGDQla52jJESbHQJIJ8cOZUaRaMven4bsV
AnGIFjCbzMMMclfbg8Qxs2XPdBpQTbaPggj3TwTMEQLiqvAlT6xEWXubc5Vi1fVh
kWkXwvB2HWOE6e1K2501PpEkZ3Y3aksKPOUbTb0x7Mbwx87YDNKJIK01sBoHSPyc
uTMNf5UoyQKR2XQfpOI4+aiZctBgNEXGjiCzeelgsa4=
`protect END_PROTECTED
