`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4VtfdD4c0zLc5QkQP3m9dUiqODckPR+e2yG/YH3VmH4v/RfbHXzeVlxHjPPsSlNt
JqwlFsb0kOwqJibPp8Oa6jJRqf9FKElI/F5mHN4813wzOfEsFhfV9j2wshBaYV2t
yXgsXrecf2NT01Rt7N49BRs6kztO1JR1YldK9p3ELEgoE1LjF0tnVWDNEG4bvrNo
4IZpNqFQ9bQRBpxk0jWqCjReMMmBbFe/7D8bnqV/PE5Ju61gtamP5LG1LxlG0tWR
h5YRNHg18RsrTF11b/ycj4kexv3UaXrULyXQF9fG9t8fbZBtzHlgg3ZBzKcpFxK7
AOYfl+EqIztgVxK5XC6AiyyayDEvvfyvWUOdUxn1RjFTy9NWjgZ9g4i4aO5wUn/T
OX/RygrbZSjYhqRMLUSvu7QRKELujeR2wvz8vC7KBGDlav13KUVqnA1fx644ppo7
lJpXXSsAbyv6x1GKyfK9l6F/fmqDHFYXYmTaneOXDN6lq0AvX6Qa27FFqslAdPBV
UHxq+eB9QFmzIH7NeMen8+6rWWH9qy7jy8XMK/rpym1K0TJ7qU6T228khC6LC9j7
Q63zG89Lg4q4roBgZ3xQHA7ZL/rg60lBuBLXsHEmm1FBWJzjT+j7beGWJc7B3fx/
MH3isBxkUiP3FZTcnJx3z1dGamm/TFoxAPGS8T3O/Z/5HWgpGKCd1S793oy76TmF
0iiHOCdkZt46N0ShwIcv4FD+YDTwV2pTH4q9VVxZl14iRIuI20uo55/WNs2cgXsm
HpYJMw99yd4+ltFUh0aXc9zgUhIbFXLXilKus1wQIhRZ4dmtlk/tSuaqs/7t2Bzg
Ol18dENRzC7pUKxtFVPnUdUFUBO3faiKNyfxQficRMyLBgHKXGofsRRKYeJS9fBS
OLWg5uoV22rkoqCqFH8ycs5jHPN5x0fp4E+s5V4ArIiY9ml8/2cR4qkgXa0pjXaY
mB5DCvN0j4WqrP8sNsy/x9BjwQiEg5VOF6xXVEJtP0pmse78c6zThdqhqTUpNhRq
n1+hhSwaCrDAeO2WWfubhBKRz2wJG6yI7minhvhv8Rozg20XZfcJ9GBpfTmGhgJD
ACd/GbAjaf1yy3Cy7w5ruL0IN/y6k5WjgGpKz3nZcYCSg+saACYIK3oeYjhmLe6b
EA4ZIzhWr8szI/z8w51eBAIWwaSMGlTtaCuIM3db1LUsNHldY5CJP3IbI/rAgcqw
CBCtEt4sXrYlQyWmiXCKoLTUxQCSllU7Pw9nsN/ccYjesPbYjuxTsV7Yl0C+ymOu
TawpeTFkPAH+mHv513+ldS/tzVdCsBXZKV7jr68Y51cReHypORUNF1YZr1JoIx/V
hc+qd//fXoorPBslLeUxW29TJ3Pv6wm3oY63YMBRc8vHkTmJ2eA5KcsK0mJBy7tI
zMc2uJuBmsT7PW2g5d9lN8KumOlLSpV6GrHNNJUZc1KgBsOwj7PoPQLn4IFKnKz2
MxuYJeBq3qlUu4p3F4ftAifO+3hN5XPk4FG12AVi6ngCbrm7+OBzsUt4qWQr+oE0
mLHEC0PWLvzSPSlCIZmPJ1mOmr4MyvoHOfk/8bQomzXRikCHPKzW8MY6fEzv1fMx
hYmxx6ymRd9/BuIEObknNlE5lobHE8TzLzZ5a7lMwhRLd62qjTFv4pKlqPvCCAXp
CAfqAJf2mHtX5PyWWcKr15I+QaoDtCa+HQru9OaMbPLHYVlURBdt9APyPkT5kTCD
ypXh8YAS+1XVruoLSRcPa5ydXO+FsKdBpGp/OOJsKdzufcq+h3/dCVMqu+JWQHKD
bs7vj/fI53JN1Mt+4F8MzGES9ospdGU/FkSKiRlzxdXPu9t94iH+9wGb8ZwZBZX5
gmfQ3lf9MT6t8iLNVQkA8It+vtyf9HboPxaVBkDw5NcmqVPeBHSRHo/XkItVA1S0
NvWls97XngZL+wHwArotFI+YIQzbGs6rDh31Wv542/LezoxEb5cXN7YjUW9U8MXt
cko/GswAVZVkHIj/S+ZiqHR1K6dCzjQOXOsz+UyKFro3WnjmaCdHPKmwHUhC5Gh9
0+5IA7bRGP9aWCEaY/wwPGpPppdSoOUExPUXyxM8hfFaqa6q5IcJJ4fK0QjfZMnh
6rvagj+bx8IZvCLJqO7xT6VVk834/QVjm3PrQlmZAvM2/PjBN3/RXRDxEu6KdDse
t4DHPi94d57qXxlWL0AY7F9VHfDTmj1GlEBg0pd3/Vg2FfshjG2M3cM8sHdlrHBh
zP8sUrqocxo6/UpMHyUhjTUzglPRXVqYtIxb8+4fcqpjxvzXMbAiQOT3uF5eBfnB
DJuoiz/KCHp2swDvU9z6Jc2XBqUjKHBAZdhHWY+dFQu/PGD34hY99UDbumEYeWTS
gAoQ+DE9SxD4ZG4BeYv53MtEpSOPO+THdocgmFb2TA1wBqusrj9J+V3s8zBVX3Q2
rG4ajkoxPkVUUrLVpu+CpApZU3lzeojDbUsMytYYXvNNqp1v36lq1nH0D0UKj8f5
tm5ajh8693ij4jdy21SE8eDTgFUeQIQR+KhU7fGoHbFC+cNnd8hG0igltclBolp7
xXUx+bjjo/IRNWGgTA1526J9mdsfujCbxgoEswV8P8vmWthX0IqaLxIp1xxEqeOs
RIr+691CoBCkXbV7qkZG7QZTVkhC65vaZZUun6vywGoZkzoF2S2Nn/If95FGO9Ri
W2uWYOZtT8buoUkNflgNZmkZ2VF8Ki2dMMblU0CUc/wQc7WjeOumQ9M7DjXcUPhB
HE5XTAmYqwiHcWSsGc48bC/q7mniCtn2/Naha+FffkJ6Jve2q6GcNhaTZErveanK
noQZ1dkMeC+HxJ07pOXlL4Ij1zGcYxPNwAmLP/t7kHhKe2f3B9aVSrtxw2DoGdmp
1o0SsPp1YeNYDqDpCtnUTd/uWvaVTqilgTuiZlIjWA1uCgSbzcTVoMYaxYFv+asQ
mvGvyIxxA6ATIt1VngeUBamn7dBsnJeeBvlK7VLK8x62+FcErot02zMz6xMNkth1
h5JfZkzwIGn/lu0sfcD/Pd/pVmbW8VCDD/GtwmtAODj1GgvPbCAnrIfab9qzGZLQ
XxqKAsCvh1027bpDBBGP03INPSgnbGn50lcFqhQUmEP14EqIWMV0BYSW0Vq24jvA
5Lanw/zqx5INimjKNCU9idBVTEbtGlrmbpv1SwspolsT0+hkbh6RyFAvrzd8vGOx
vAOpMd+mcwQAFWOOxRWfN9nUuzeHBaZXUac/oaVO8I80+QjX3ZkAzfwEypMYUlaj
eu83WQwjC1rBE4A66NBY1iGuVD2vx1D3SHX28VoayFJUcGR5miC9qkogMwChBQjQ
l8fqb5lQFQSXBDq8zkkVUIaJL4X7s7Y8wp9HWACqPvSNJEa+Zz6lnEjjULlWVA46
bxDVhnW+jikqInFiL7g0+JKC2PhaUh7L3F/RNeM7wkVGdDSRSViPtiLsn4u4z1Z9
3hIvv25aINIgj7g9wdFTZRJNeDHcYEM1GfSfbhpAuILsnkEXjdgk3FsTifHDynOl
UWQ2Ns7ia/3xqwfMW7z9gqKPBqfcdvDpWSHGzwKlJAs5lAhsBDQKBIo5Cs1XDEH3
t4/hiBlC16zvrWfQuxbrm2MHGEkWu4enxZ+6drVgzaTOwnu736Dz7aQ5fFGgm+Ac
UhJcvDwQY6SwdkMZqjF8YwEW37N1xdzK6b/i8rAjGKaUuuztLMVGxS4yRpfjyr4/
Id6Oche6bi4E4kGfdKa44Sn9Skcf3zk6IPVRN9cnVkEmeX0audv3HK8KU7lGyQOW
J3CFxpB11Kk+QnQ53sETqnbG8pPlaD4EOYj3N22OcotNv/hiykrWJO3nn1ay1eir
7hf0Ek4PuWxKfjSrCE5NrhTu8uiU9VoNbX7A4mXAfrMLv6OvfJ/2lqDrpb1pzAij
LGtYQzm1MhZrosWDjvj59/a3JcffrKOp4SQvf+6gQyXzn90ugqmcLCtDw3dXtvJ/
RLL5XOJVBWaXkfdnedWIBv8fLcmr9zlV8LvQZlsqN8+zmfZnssxS0CNJINwBT7vW
EgB4MCaW+HETYSKmEGdmFL5/JDAcx9MMT4wv4IRURN+0XdFaCAc5vDl9AjjWJisi
zFlW/NoK1KmfEOnRS5eBQ5okMhxOoyQwX3lyMMvDimaAcvQWq1Jth36A5nFQTrcg
z1SOgPYI4uHaZbvwLLNlz88nnH/ordqyC2Y+aE/nn4NWRzmjbt7gTnCJ7SkTqd1b
piFeElCFey39wcy34VkNk6/46AYQwuOmf+8HEXBgN803EsbkwIfXCbhOHARAOvG3
o/EhOs3qYCEt7BW7MZP/OPfvcplTuRtxf+AOGe71kDvHoHinx9m5zoHRBmoPJOft
7Yp4t5AotAmnxISEZQrvPgpb7mUeyqIIwOPllnlra3mtEdTPS8JaxryJM0akCwi0
huGkPpgdecb7WcCiA9ZMcH9III/5jnvhQhjPu0nLWphe7VeFjD42SxOw7BDl0HTt
XfnFr3FcVmlqZ6r6SwUBkSXbd1PJuEE6B8aCZcZxK6hB8iVyg60y9uA6KIyix720
ruC5qmOx1nxtukwgbVbJaJb8sT+HtY24P29W9doZdoPgKWES8aoOTFlFOAFUPhcO
ZDIs3erKxQ2gBLP0JzZb+KWRVXtunIa7PS5O0ZDT4bFX9tQiznILPmmBW/3m79QT
4JWNkhuE+3w7JXaLijCxy8/ztUnluU1GUSdADuFLo5F4ZT0BU5JEG9k5jAkP09h9
2HS5h6u7gshmEmkO1pCZLNGViQESr6GlRM3Pugm7xbxj6n0GFLZgd1mYCaMft1z7
QGOmh8xMZD1dMUYthLUSuQxRsTIeTqaRgug5wdGivm0B1oCxKXfp9teIuVZVI5O+
SuaxtDM3SczZSwce6PMqmKVWqtdcEJv2ILqbrABCdrMOctap+vFIr9IhUkgpd19q
KPwNtz0Y6tsCTmBNki1/H8WvKzPogTIpH1t9vKxxisALeevNgHzDX3V+jR/laIEb
l4pOdKeqIo4yrH4udHKP8+L7x7TcLiVQgdbflXZ4L3dHIJJYGG679oejmX9cKlUU
iL2h4JnZMu0OWT1TnJV3LkCVeISQ6S/btsEHLrb0rIVQEUZDen3nYNJNphV2wW4w
TFY1Lu0OtABbGtPBean0LUinBMYm5hFnMj+lWSVMvAv0n6Ok6M5ZDHI5lB5r0ezn
47eeZzDGtXDngbqNrhGAJj+GySOrEQ6eUWQ/puNtibx8FlcD5V40max+OZro6pZx
wHxlMNLtLvGtE0MTEtuV2dlvxPKRlRvmqPCSjuJhe2jBBSxE0QQUCzFISVo9/wXt
2DjdGwQyGUDS8eYKu0GDI1NHLh0ZVXdQVjMv6u03qQhcMa8Do76SOY+yXa6VJNGf
rw1d4DYAlXZdGz0tIxOoHokcPYHZj/OF944wSaLNm1/budtTTd7wRWjI5osDxafE
trpZonSetmq2wIJcnBzvjx3Qx6xp6IXhto120AVy+2BJG5j5/9l3tlgq7GV1tvZC
DgVYmMvuqm/qtPDi8U2JaDhKXw6+in/RYutLxSj0pLngvmGiIMBUuPKiIVcy4dWi
RFx4+a5/UpGtHZ8hVupM1z4V47z8PdR61cXo8Wv6jaoDGJiuAB3Ro8N7ATxCzTZV
fCut+mLuzti7wZHP/nBVPq5HtsABbQ9vzs9ii0ul1wfv3nZdVI46zwQHdPmnzvRL
Kihaosn6K/lOuMuIgDUcqS50Vd/bYpgL++F2hYRU5l5HpOtROzex3qh2MEQ4bMR4
chUa5d37Dri6PENENjdeSc/qEtl7k7EsoWPRkmbLy050ZVxY0h+UmqaLm2udExM4
mcufg20EII/wmU9ZudQGA3ctbbV4SUtE2fb9okJEt0bslTIERY5ak6HuDO8qXILJ
ZVnx2mHCOJadZMSVPDzlKBowZpVTXPtX2oAinaVr5oCf8FdVDCU+o50csV1rzWgl
eMeGwqJVO9eSxqaz4ZZlV/UgQZ/7m1imr95/IDD5PncC6TKAHF+4ogJJD1aLfOGo
JUg7sPyS9Ej0qeOoE1Ih3QCn/PpD1AFE2L7Mozdrv0Nvlel+2V6fXqLzbQX4OZ/i
j8ts7h0oLtxy0oBtMafv63H8zAyevEXt9Q9E2uHjmKKMEo7jP9SQpvN1fNL5/gNT
7pnfM8fPCtEJZ2InK0JcJ0liezNg28TqRLfEX/aitetQ+TzkNfXCBihiKfJRqmR1
X3qjEhG6Hz4rIYiBBwTBtBcH+c+dH/oMWVQXMKmGG8ljSpgQtvao9r65P2sDMli5
lgtLn1jtTG7VU2OcLvmNUudECsJhwLTdr4Gbui+5Rm4E439XSmtLn40hvdojzlOS
NZydzdRdDMpfhlV5qjHD68zuNwyrtoxd2b1YJwRYkWYRdtjVt3d0ZodjYBVmBoFB
Ogf7kC/p01z0PidUvX0Krr+x41nikT1dtRVMA9O49XFcbWO5A3bLqJyjTDr0afqG
Tui3PgGSMvvfG/gLfoATik31AYV7abwqLEFxuhMttOvtjvDKQ5BMBFzKmkrp9AAC
Tei0flli2RkZXy5Mf42iLT4qo7cm1E4KUV7pby4WwuMCXde/v/LtlJwW01lwoIen
YvXukVeBfyHxH9omvLEqy6OwmGVGdlo9uEfWJc35rvsSlY0dCdDwa6NFziYjbQ4n
LJWh/O1OJJsY/6DecHR0Ql2CJovC2og0SQOuCczXqIc9rkDpcnPBZNtcENDb9xl0
mD4e3v/8DYDZ5zfPkwJgktZ5EJlRZfjAu1hjuyV0EmnczB9SNnCJx3UeypsHQvTS
aaC1xeYWHS6Y/aYILZJJK+r5wSMMAF9rl7qZk1kHkcnXWrSObFokX7LCJbUCpMr7
hc43WucSL+kIdFJ85WZ4/84JFKl2N1PrqFpcBEkeCYCCUHB9WHBsaEtR3PveGJXh
FJh2MGezMjISZzGnzxuRYgdc7x76T4psdwn1LuPdVC51gS+MOhIVWPaGk1dykXv3
+z1RgSrIZeRkMOYKewYj2/Q3nyD9Vxf+Ce6zqt7M1i2VUMtAS3do5GNNf+AtGQHH
JEa0tTocYd4JBPzZCGTlLlbVPRVk9evEOC4CXDT2o4a83jpNYnnD8o8ItOCeDlhe
XRUBLe3hyyzwt4ydGCCclH+a1+fKQjeMQjvNES6KLRmNpdBQCMqNUQlK0ytmazvd
9ktry3gQlc/xVomgUNLyDzw90xK17Y/6GUM7K1bmF+ZeO+ooadc92ZuRyRwgxvko
Ze+MpXifr/1Fr/Ojgu6SyKZTXjF+1jNyEw8zjOTCCv1VFtG8MWY0YZvDvu54RX69
TDvRZz5kXzip4B7x2uizBBo5q9GSpgo2l0R1X3BTyML1JkOJHPtyjD0AehdqrPc/
t+e3H/wkx0Unq1owPKRwXSS8MEhGpRTPzEd0+QtweI+yGefpjS9mG9RFzJH4qkyv
sA5ZPRiBa7KGdIduXfkzvlNu+pYh2fLFXMuZiJkm+DBx/hr6UrxvHTAd2vIrOuZB
gb04fIH5pUPm2hkWkEwAtC1XR96cqY7uwKrsDP4aE0Q3oXcnRHivD0g2iu9BlX2w
YTehHS/95EjAaWjToDJ12e2/X/QK+L8mKqUiBDifv26gr4mvuSLrexVSpK1+Vuj8
cZ/z14xV/BXmMR7f10sZhkTwsKEcP2NurkBa8RfaxbfkenGfdEwl+x3GAGAlBpUN
3dM3c7h6TVPHGxRPRyfHOBy3ghkDT5+SJhV/ICj2P0KZPR4VH1r2AXKO8arcxBk7
rbO/bl2yGWfeTOg/CZ4J/Qwu/+cVvHqQBSqPXc82sKiiJmwnpNrgJ0SJq97wNYZ5
WP6o8fTVyBk/ODXwkwDTnqgGnsVsyd3XVS/ALayF2tK45zbC6UiXq9OaNEC0MUti
FHAduF06MiX+HRhFfAMk8TwEQ2RhhvLZpsSKIzcjPlyzgAJp+48PMwuN6OUP6/Tr
c7rb2EAatZNF11vAJC1kaCwJTSQNYCs0/OjgDUPGBHtKqSg/VdtKQvm2Ybl+VWok
R/9KQTxjc8fc4jXQEyh9OWnBHTThyooyhwvQir/AWVsA6O2cYxN4QPJ2ldcVKtgT
tmHv+f6Qd697Yh5dt7ykeg56fOizqeMkoOR/srUnQ++7ck/5zy7fvVqMf2BCTvPH
G+CC//8Ytpz4pu714sAzrK428mvFv/05r+f1WS6jKRYxKl4hkM29k/wp+2oONrby
/KVtAR3oXLZ9SmRquCFyG9JrnUlH3x88oTeBmF1IXe77jiCPmBuMdr1CDmS8vdxC
Sa1RQaQKoST6oZPN2BM+zXQ4Hg08Ljf5KoAIy4Jf/HNK/azODzeSUbikId0612F6
qxNIBOvD4PubADrX/jIvKL5tVYcCYUYSi44i8BbXGUnq8p5DkNkzVwaTmKD0iLkr
l4N1a/8oj/Aydt+ovVwnstnN+5quk/gj4ERMp3egaKjWl8KDvII/cC9eZ2ws/PYT
ERYL9P/UAKDt7MA++Cqg0dUPi8x4Yh9pdWeDIo3lm1gReoAAN9qvstmQ9gTwCA5m
BMom53UA/XMI2tMqxkIlQ9VqaNl2AGcnTpfiEZ5dIKTqAmnL5gIWGSIVJrIMBz8O
WNDXxZT3UvBk0IvDWuHpEve/t4SSdrTNfLx9hDBoGqekvyXV5njSzDbX3Oc8w7Cw
3X71qfvG5c0ndk5efZcFnoM3e7/fLplPXY0vb+qD1zV+zlaHoQKY/HaZ7qXlT1pc
yQGxNzmxSpxcIq15nXPH2vTime4oa07duk3tGBXd+Ebb1QggrDZa1q73zCS03qGU
SU7sBuy1qyc6wsIexbIwrLuzKATre+Fn3eHHlBoU/hW0NKQQ7i+GPWvN0GBnqhN5
TISDXImd8fCV1zP6TEgN0v2pCc7iOk2OJAwv2vlKruq2emAPqQHD40GCIgN2LLFa
xl1kcrK/Ox+9ZNzt5erT5xcp8255g1ugg/3o3UKIM+U3OQUjfw8N3MHhWX9P8Gfe
hnhKaPi6dJbm7XNt9h8HDaD1WhlmqWXQU/wgCb9k32UpaxHX8Hg1pDMuhBpUAgKn
A7NkcTNoCtBH8IFi3FE9AJ2WwYxgtXa15HReSM8M+3tr+CUvGrjZWXRisYN3GTwj
DYrtjK3rd1EI2+gAIuXseFAWv3JyO4bkrilcBhWewObaHUurkpjLgqOfiW7uYO/6
t2+6wI8lJTKa9qCk+1GNBtfl4TukgSLUUipmQ5ZRg/vYjLUmVGpKnJ1Cpf15JLS8
tTMyb8GH3G29QlhBRnNv+vRjmiBe7s/ZCpdlE1S8O5OcJiqb5O0RzsPFanwgb14F
n69/Ho4OM6aA3lqZWo0+me/R7BLkfVR8l8BsHvME+FJRqzAvxDjNUA5qjIH46In/
qsd7PX9TpOFPbfC6vruHbe1ALfRmmXbo4/FyYVpvd0K3L90gHhPjbAVpev0GdYHk
VisHpWCTjCl8fcVZ7Q26H4My4Ss+vbhMFqFC7HL8dnDwxYBz8PUP9oCJ2awsH8sn
PmxXeUiYdfijkQbA3EN2gaQGIVZm2xye5Pvk+qAUr/rjtdaeC+BfrOVnn9717hHO
j2K6UzMjWKajWasyIopYKzv+zwo4rYPpGCPY/7+AI3uEko9MX80Z63Ao+adg89XB
Ctn54uxiKn6HE0kzzzoI/GGy2Iz9z2/c8xYkQMdDtOdalx8Mrv5fYm50HMw5PCJz
AFWJJiXEMYuGt8FW4fciSm5qWeJLhH5jBBOneEGUFp6ZaME5uFLaEpEhO4BcvmbP
Vb3wJWf2l6RddMGf/j4n29SG6uHgMkuum28oi/GBCauEeM2sYGApWEFIPiENHZs1
HXKksfNXYdyGGyNCLfw3zz1a9R4VcwNp1xHJVknnA5M/X3/t3uEwet2oQnK3wOQZ
xGZN264yCb7YRVY+9H2fVWCXcj3bnNLDjMbgO5FxIRIFWxlW+S/aBWTxtvnQ76My
SeR/hRJ0pWm8i1T7PTGJTvySFCLiXb/wiKdqin22huGeY7b2V0M3RC7hs80UOF5y
oeo9lcWZuX8DqELywFB2Tox7Rimxz0AKj6m8xr8IAn5MpxfZMJhpqqwGLnzW/3Vg
DmT1FsTXN93YnXOrjzhlj3HZitxkP5THALmf6tQ0ZgGNhfe/1DGYUStejHSjSQT2
FDgaPO9pP5EdU5MhH5xwYZ1rjx0FtK89N/Hd74QNzLAi53Z0xM7zAxtq686Dul3d
niFhKPnnRYWoqgezHu091DxOi7e1uaAHrPOTNOcEOjaWRqH3jGfKdTO88mdokArt
5GTolZ3ViEhYtVqlrXAv8U3eEobqm2zRN8ww/4vDwB7GP3FCLAw9Ma1pS3FnPrlu
rIk5eQSt+IUNx2PkK3HfotH8dFiRbUsTo/K0Prv+uOSPMmBwa2I3z8Ea4C9i/A93
OPSADefchQtjz7Ho1QNW6e9yGO/QV7ty2iaQ3kPBChssTGNw45VXn1nMoH09v9G2
/7ffak2oiZxSBpG/o4JsAaANKorueLnEpv6VFZ/Lme63GcPdSjk2I1qoHF/Kdnc3
1FoHNvGGtJ/6TMUu1V+penuGkTzPC/rbwBhGGrDfozf44fw+VDIYc7IIDMO1G2Ml
0PxVUD7jD90OhoZL1MImHQ1dHv5wri5afH40/bnyYijVT16mBKXLqPUfic4obvmO
159/NWqxzIw+a9BUGmrqLwZUy275WRa65Mb12xpMFKVuqwy0yS1JGVTogzOs84rr
YBVr9KRa1iO2cib/lIx2A3U2Lvia39yK3fhiDG9i8DpKv8hL/6wHkpHfMv1aoMVL
kO8V827DtVkfPiJhcILKFSQZMdxi4Vs2nJnaGzPZigmyIh7xOGgeAlv3lsn+c3+R
KWSAijV6gbLAAepAuXkMPmwwgo0hQ7Fr5rS2D7BL9Ql6QtHCz7pPahVNev06ZNhc
yOGPiEzLexJAoxjsLezjybBlEZfZx26hpB2PATJxJ1XrPshE/zI2WIM6ZwwBwYga
713FUZYc9YIg0mnS3pAR3HZJWNPKKFAt6WubcWSTUJanlbBQzpcd2jPimPThkSlZ
84r4DHPbjgB68g6BG7NILG0PfrrsnT6aPCG8jBitGhD/zVlXfq/whaME/ipSqFIn
86PqhuWLiU4zqVT0xk/yQjXZk42kDk5qcpPvKs1E6AL3RtNIBPq1DEnD+Rxy+pQ5
jRP9rxprpGdZzkWCDln116mLogviD/5zcBgBSv8X00wuhtLeDk2iFe54JljiJoht
j0kmxRI0cxGCQgQmlK6LrQbr3vlgx0xTZZGrgtS/8reRPBAFmQ7Sy5W4RR8pkCOE
ZZI5Rr89ASo2b1iUvDlOZd9i0bm56Urmf0PJz2dXLp5q/jg4CSWsGypXvBoXSecL
vCU4tqT8Ly+uyo/NFXh5MYB8lsRLaEpGqvZDQNngHwBvlyIzM8yldIcLQl9lJ414
/20L3MJxqjycxHeZG9PTOphnZoFqWa363WWPb1iy67r7RZ5Y18cs8rUNKQ9xpbaF
Gj6si6jDRsf2FUz5h31H4iRwOCx7ZUBBcivrQiyHm9gzpp8Slni5l4LGF854GSSH
5I05Eop6z0JwkUywJSv24dUc1zuKaXdXWtCqeYUN+po1k33wl5vtR9QARihbhcDO
XTCr4TZ6Icnp/crd67h1o1/eGxpmjenn7MwrJ+qvDa2es/zNB17c8xkbhE8H2ak4
vzvYY2AGwOKP3FHiDpIdHLDoK7yah8ezFjT1sZRQb2Ca7oCfaXeq8FvsqaHMxElD
GjBiTpiWZsP9e9IEJFE0N4qu6nuERo+1gosCmm6FK1V0Ntj3v3U8QoJDA7rLJDLw
kUV3Rv6puj+3sCKpUOqtuWapwekjrwHWOhLu/6Jp2pgazp5yz/dDv+5A11ubry+Q
vaCxTaY9SCTTkNfegExU/864ZAsjWPfiMn+pNlPsX9y3t/npk0sLxR5oFFpl3xQv
MXuYKHdd3DomCHiQWqhTv3q0012Uc949TJZiJzqWBh//h/cw3gOTSMHU/lULkHQt
tTAxCAyYR6KuOgKRHMJzrbfbUhIKvjuC511P8T6rdE2IsnKa8t/52VjyFsTUhlIk
Yxt0gyL6xOzLat7/z1YRorYIXjHpIv96wwqouyUYYmI5KokBSOCqYd7Cx4KJAUZW
G3s52EhXlcftu3Y0//iz5QI1dQHDb9Z2sGsoQnAm2rRMLa51MP69MZYsAHyc4MND
ouVa7fGTkevGCnCSSa8tBeXnnPQaTl95F928DxvzdpPOIASRPV9IIM8vnYEryW5o
u7rcSNOFdY6LHls0357h48xrJizzUV9/UvESOelakYlSj/oaGBFz6/NhadqwSuP3
Jpo7DAu44ikTHZMe1o+LccFEzthCj5XhAmp1vznC9N8QyCRR3PPM8w6RAKjcJ3Xn
owCDUxoXdn4dE/KVYuS6R5/XyUvlsModnc/t0ZyJWlreVRysqj2Ut8R/1NeRg2A+
qjZk4E5Q58LddGKnakMMlR8Hpi9v4mhWcWUNcxv8lFLQGLX1CfPUL1PhO0PEEqRR
+zUsOMO5FpT1ONjri4IwSjmoBkv6RajdIWj0wV9hHy4Bz3Ipc68s1oxKU7q3YxsC
inO3gldsw5rckOAS8KtG5KgrcgUVTndcIPu+MAY74qHMi/kw0uPW1m18WCHQuSk9
e2yu/KE6lZ34QZbmtFY5hYbdVwURY+isEFpIEpeJpV0PsHBXCDKxgOaUQ8nRQOcF
vQM5viYV1sGs2M34bz2M7Z6zk8grSRXxFEMQABZRWNpe14F7pD7AgDea4d9HMAIz
2f4VAKW5izIORk0JOqcIGQo/NrQLOod0zr2UOnsDTPc9Ctr9G3UDjNcmTBPYs6tM
YK0Zk5qIa1jEP7Ki9DnjeTQWuT9GIbuT9TIriQ6EksAhBoctyYeo9CzndHg7bLhn
FJ+YCS+A26ZXuFHDGNmMLiCbar3pgBbKTb86cs/Bycg3WQTebblLJemZH3i4kA38
ipifhDkq3q2YII+n8opmTGTbJrDP0HqJH+UyzutrO9TKHEVKCC0lW5ROdSxUTlVf
s8jYn5my1NMMFjs7u127UCLd8NmnWkhbCIwmsrbiuuKxqlUX6V4itm8AsVB2lRkS
mdpBOkHJdBukU8Hx1AmhfrB//i4dSe3n3haFCMZBcsHbnJUu6PV7KqCQ3qZ1U7xg
jlYnu0TXgLpcHbKy3/XOEpm5RuZGgIkKXgYkYeiSjtUrRL2NRI8xI9tzYXPB+xhW
RuSZkKzRKmSkopYZ1GS1/MZZb1kkdbRhmUDTn4f13wgSTchyvhx3NbDN3wWK/v1Z
DoBMPNz2m9ujBSfEt3hkNRYzyM5RgXMd6YnR27KnVNWpSraubQLPKEsSEyXU7izN
xRS6KPXe30l2pHzah0Pmz/fWaaYdI/cmugfnpXUcG3/L2MdwMZfCcTDIkHfw9jBP
Tqb4wKnMCjZSWgV/KrUYd9omjT8wiSyPNimrneyWx2egGIzQD2l6XaHvADATV8yD
0GpGgdR1vA6+1ldYjLcadnP7hf5ls7gLX9EXxPFzrWB23FnY35CLZz5zFaKTO9o5
0d06/b7mjsnYoAvToS/tFiUIR5TqpaRTT7Nkxc5iJO+wnxPBpbUe9TWBml4RrStQ
xpEr9ClZkKnP5xYEwooIAfhE/3G9N0PaapUOZsTwcKfAbRKrba9mCJOw7LFionJb
/qmqjDv+iiXAgAcZNkIM6nCv1gjbDLWAZncTTca2fPbeQF3Y1WRIO1+a0OAgZpdY
vXQeVnsc7cJyWzzNKxsKbg+Gxu8b5T1881diqKxSOnThw+GNjgziEro5jAgTBHPo
eMruq8ngAWjYEHpvlQsGATHC+YXz+yZixF76tcadPiMUmX8jM6/w7E+QLlUyZB2b
YACdiCoAO6jU81ZqaiKE1LWPezvscm38OOJMFCcJ+UCXOnCZhjAHccvgRMD8OPIt
Oj6fvux4Zywlnit9ISnkfcpCHaQ0LafzlGNDJqMvRt63kzwm5ZrMl6XOiJ3NiYIz
8LklAfK0iXn7oB+7yI0aIa/1k2+ZIAPbrSIIxFQQs35BrkCFfAaK5EZp1ZsI3hCp
DsXYD5Cu5ys2CxXZgbODSjbEILdgMK+YjdHd15mxFmkIS603gYhS1GcJz85lP+tr
BqKlSzkRwFl3hfDUZICsxrLLm0keEbzdsW63K4NCPeWIHSiKlQkhBauVSKZ+hvJz
9rzFetLKD/pVl5F4DC60vax7RdljA/FR2h5u7nqOHQkdnggdRXsSdhQvgetM43Z6
CQFMh9P+QEuqSIvU+Fe6uNJogocg6K6C7r9r//9gmMr7ZIsI9R/xqAOY15Hoy3Gf
HUy0/5XOp/taCfItgc+iU7AZJ1jBVPW96G1eMPcSjTZMfnlNIbfEl6xGaqqweLZ1
POgVp+L/PCqQoV9w5Aqhl4lfFiZsYdkslXXYnNKvRLI9DcEYt82UADmCoX02KcdK
/sYyU7PsMeJHZjzgU44CvRlY+IrB+pT3QIm/+8qRadMS5tSHvFrGgWRtgSOdjIVA
zZA/QS24e3w3fyTwBdXkBFEO40Ahv3UMl4U8vpyr9wS1iaEjLp/GA/7p2BZBwihh
4aXbKwSmgwlxJQQdVI7yWUSW7VNjhGGO/dYOsDfbWUgPIrpynFHhtQdmlLC/etX7
o1Xk2ILa531u2xhz4wmJ1xBBQSxf4XkLnYtQPR9SlimKtucdSfGsKyVYmIvfjaUQ
jLSFDiNqYB7m2pQC+v5sVKxjm9RuJc3SpTm6y+2CfJt0KxvCpvIetKPjtnLmQvsa
Bo0eM63Hqab5eO9KqlVS1bEk7f+0/unKaUZ1hQntWWBYjFVXHDVn11dqvvcb/Txm
BScVVHWK++TMZIiIg0gEBD4/b0sbWLg7xzGDNSSkCbiqN5KEFDXhC61tYi9OJB1U
Aw3GK2KLcEDqqhAFp+IMGwuN4giFvloJKQr1W9wkOZwUDc6n1Jq/aLTp1jcOBXTd
FH+Sp4ETHzfwZ6+xWZl0D8rC1K/aTuJVis825FzI1dz0JD12ZOkkmHnO0MzgIg5b
m2r5SM36+cUVBphmIMy5K4DfPVTA1Eo5Hsy7l/v2kvcRmLrQ5J0e/XVbVKcyoQDX
3Fq6OknVG69xBL3uRYoLEGLX576vqjTaa8z5rWdCXLEeU6ehCxoHEE8x+aJodX8h
xfkS4BYn988Mvwqn1+psJNIjxW/68e4tyE3w7UuqsSWurDydIsBVPTknEMS1+eQA
ng8OW2ybIBkQC6lTtgmoiKb+BzXXLLw4s7i7ufKBgZZ8H3oGfG5JYvtrrGu0uGer
0kfihoUfUT3dCtPEIe6q8KL8XSHoBZroc9YK3hvUY9YUiwn0P2zPnbXd0JmX1Wgd
jt5wx6LBfsJCcGljnoHrk5IeVDInVsPfNypiJ1iE1U2DMq7et20vre0gA8ncCjzb
3K9oWDBSFFmPCL/O43qYk6lCMf04Aga2u+XuchqPupIumKZQkHert3pmMPJK0Av/
kNdHTkGBvoLCHedfM7u3J55w+wOtCneHyqc7zBlgSHzXN4fnRM3F1zR28+NmUI1G
AfutSMcLAx1FfPp4Zw9+w53HfQzEJgPLgCLDITULZ7M9FDUHwOnVLQQZP7Sxk2tU
lGlt3rZeetvHvtXo41sCJax1c7TJmNNxkcXy5jDpDE/QQ9UAA949Lycba3lUYQZ+
zJmeLlGigXPtfNyccRfA0liMpGri9lsnQlV3AibJ8AyXh+uhGv15HPj94RQs+r5I
2vDssZTC8Sf3uoHNPsoWbWBKL6W5gdL4+DhTsc4kPkt49jRVCKBxqX0WL02Kspn8
RhQwIfOMW3Ms/j1c+F9h/TT9g5gFIKjn2xeTqU0uXdin8LXX4mXC7d6lxuO2cG00
BxYGx13P+YBM9xsHzq2wlXjKr94CKAdHXBMEamafpTkbnAOmtcY7AJfSt/aqzbdQ
bP1s1BVvQj2yjipwLoqS/J1YhAd7VTY57mzO0g6WM2ItzNAPyL38Kb7HkxfX+hGb
EJG2myDjufzmPBBcC7mCRVmMPKLULfEpvChDV3ie54VmJ6hAoECVm9MsJkBSeRWR
l5vNEWFyNY4k3cphiTre933Tx4Dd0Xm2YqCOQo/syXxt3WJn9NRcJC/vAnYAVWZ3
AP9O5RvvUuEu5C97nNg1AZv8G2638A/bWMCaYrDXNA3+jGHuZim6EfNFXEIUgqHD
triN06fGmOLRLv7A+m1ByHl3J3dLsd1PVNtFXQyKabYc7lx+q0orKmDgpPLPmdl7
C9XaljLpL5HlX5bSl84dUwvbpv7pG0Wff5B9cDocIjvNZpIdeZ8GJvPzv4S2bURr
+uCxMT18SEnA9cRPn2kLd4ael3ms08o+hV2WEXLVAU8T4lDnZ3biv9R9c7WPjQ4C
f3L5szNi7u075OZraCQ6cdC8plte6n40yi3r6STcKhu/8IyiM4ZvIsJv9DprK2YJ
vO14CU1fm5rG3/+CiolmRfzMG/9/5m6vSzsUxolfLladoA8wWpxmB8KmfmIL0nHO
LsXYb+ZAzBgtRaSHechrmedpAT/uP2m66Wv4SSM0An+fMIKMwzbecZqFILhoYU/K
VXnkDvlySs36ofJufs+2Ok7Y1pcyiU94zLBh017XrQQGQlocYhxaBQugxuRchBM7
cTILIc7ZSEJK09RumNFQIL27L6tzLVxcPvmNYnPTNMb9vxsbvUUswUNuxVKXKT6y
6dMlmp2T/JqE+6+HZOM06kPP02IW7RSBTUXQJ/c9RWglFlDI06nqedkvT/8yqTo3
0UKkDRquMRvsBquNSSFXRCU/JDsdtRtI+/KiSXPgF3dJRKVk5YYqwBobd/F9EX8j
bSwjtSO6cvAlIwhpMocPWNrDneClILSRsaOuotLGkMEi2tL3hsYq9w5om1QmiOhF
RMGhmLQ73T+dlqXLdqAoiRag6X3LsmLce204k8LUzR97hRvyJt88hT0W/8fHeW1Q
bVYgE4rk+VtqHcNTTrtSBIWE6NK3Ft+7uM3UtHKcTOccqyEGhyvd4+7Pxhs6PDGU
pxdJjibvgSSbA2DhdfjXS6mLcbis2yl+5Pntf9E/joak5q6XNyX/ZEuqDGdb615a
TGKRyORHdeV4NmbvvkphWn6MNC9cSbT9ElHyp+cQkCI3DQ2VyfGQZcofhF8kW0Oy
VVLGz+ctwel9XB3JRy8YW9p6nQ7OQr2ac421/7YQMnyj394pOHaIpg8fPZFZva2T
xfIKhsbmmyNMpTA/mBv6Ta0cexhSVGLQYj1MSi7k2ClNU8WZMrm7edSB7iG1DuxS
5olw5YAL1Io7xr8TK3uoqVNDs7V8XduWmAiBkIC1XSjQwCo/aflz3tltqU5ksDCy
GXq+7tHqMpikR2oxpmXYLlP1ggjApfzBbjyuXVwrn0G/h9bdGgMDPDACt/wNx7m8
c0Wm5AUJob6cnb9RVTc/9cQaIhm3TnpdLXsTXmiM+StcuxjbREgyd6Ry71pYv1t5
FL/GWN1fccXnD2Qw8TQ/yJ2k3thaUy0SOZPbO5rAqp26RFzaw7R/2nh19ud80OwS
v/le6bo6yriW4htG/nZLhn6+TwElLVz0jfRYd4MukUawr8L1zUP9pnxgzpQdXHHZ
DXZ85XZ+QrCAI0z1L6IKo1gOc6blRy8MRZZ4EtyedbnYtZ/SMsqEVtb+cUJOv6Ma
ZG7tRwU4Tiv2mMm+1Z/PyruF3xhqr3rW+nK60NKaY4QEL2c7K6EBvYxd80sEK2HE
8Eu23dQG8Qa1gDNQxy9LYsLZyL1ylEujvTX+ZNcgc3aT3bZ9gCcdfQdUz8C/bow3
uQqPFd1cMiZg+CIiPIxrD4YdRjGE6L28zfxyfi0sCBBHqWwScvB174kCK2DJyVg9
YWPy1OI8j0HPD5YgdmicOhlD8+JsTLSrb1pDMQuKqVeZtzOOvNi4KPMhnbfHTDsZ
t8VF4WMdCGklGktIHDVjxVBhTc5aL3M7tSAfMcv/UfIfvV5tH342SIzD2nteBkOD
n4pdiHPOJLf2LSzJLW6ef9EAtKwNS9UXIsXO6eIOuo2MXokcQqz5xNeczhpF356o
2OI7v+V4aTassHDdyRk5SR8g6efzQxp3Rh+5YU2OAJePfLwqvTHGgqr+naruigv0
85XEVCW7sErkKoNiANAF4EMeN9lMmVRLd/F4FWsJYuTYa3WWGsz8eETu9U25RRpZ
pYuEP+caL28AqMDhe9Kp+JQKXY5EL6NKIzvWuO9E6HCFpYvwM05ISabUhZRm8NJ2
9h/5+ahr4/73gOeR2DhrvHZL+IaUHl8yIPdprEOBZUgFZN/RF5jNjQhLmXpeHAQ5
NhoCal24DApE5RIM6FHSdgAbJrGFviXxNkNiZzNCJzkmLnddojQTq0U7Lhjl8yvt
1rgdFan9PA7TFfTAvfHwPzQfTPdQglnLirP0/LnZmM5ssM83i3KHr++dDwDPGzLG
w3YF3lOAVUaQ+kL4bs7Ben5OliEEqeL1ga8jtjicKF8lZuLamBfTtj8S6PhgfqAQ
UKP4pmUurgtToINST3ZbgJObShLv94UXb7Dl8umyLNCzoiEItBb+FMcMSN3qQhei
VSA1+xVN4XX6vcCdarbSv7VO+btzYVYYs+L/jN5A9WIxFVEC7A5mnJepO1Z9kVvv
setLc3QIizjkMUef8YvYkDZadNSztM6MnDyHWsFWzXWaJtgWRvknRMz9wT+5dpgK
ehJC3hvAODQr2fFd7CbAA2QxkP31BEqmivUymsQffTEFWtqwEi3kQdvTlRCCPo7K
UreA1U4gV0j4OiT10jcOtvE/zyGXiTcnS9Yn0Jdn98dEF32Fm1lzAmKmhA0/T5iZ
qRzkMWmHKm7reTqEEDid8GzbYWUFHewFys8V1UHTH2ptIKK1ScRwCdT/5RR8Pmxd
sYtMn4zcohoaLZ7Enf5AS3xMNbvWwhgBLifT/D1If31jJwKAy9L7UzxdQmDAJlXg
UrbKi5lWIxOwjuoF0vMGqfJ7//xTabS7QYI9jZRZKNaFalINayS6vLAX0wUg8g0j
Mt8rQPebEK1JaiG9Lh70XCsRKT5wZWaBnMi7o/qAwwFUxavxgYuG0nEfRbSq59l2
ZRJuWgOrLKZiQMIxT94KFbRVOjEmHy+83YJBXng1cwyDnEnZQmo4E6oYXOhPop7S
HidMUf+wey0tVd0VElsW/ezkjZ6PbaNscMyod+VJFJ+PKHSLsNmOkN2nY0sYJMnm
SPxyar97eOZ5Fl9PXEPbUhIgrac90Y17B0Tca7cg7O4pe0cqYJuwMbyKWJKqak4D
dpNMyFuPz4nZjimcKvJPdmOhs5GVZGTD88dN+HKlPUl9d5umO9apH9lsTupmShyf
Z7Di+doCmhR8mBseXRtKYSI2aiulG/SKoucXcSdSbVkV/xkRzqu8/+4vOuiNOBwO
W4VKaBfuAjl/B5R1GuMnYa3ifhM0Iu+/2UqNZXG9rgN/zT5kPSucfkiw/dIRfNBW
tw0IuEfG3hTv3fayJRI/OdzgdrhLwpFSd/11vrsMqpx4cxFBtcmi3gyG46kmnVRq
SYi78ywovVSOnkK7Mc1NsCBOVg68q7ZcC76xR7jW/zrOz6cSFGOBpjB1qGxDRp3O
dBwrPC8mifkmy8KGSi++sJoagBMBsziO6isr+XZtyB3+pinnB+mvBG5ytAL94oUC
HwEB+wrBRRsLvsegByJIohdEd1Xc7zDnrylcoKtKxHb/cQuN1C18OqZqEUbhHoog
QD5Le3+95magddelOCoKoMeVwKapDB4aLPhBR/5RbC0oS+81TUeY6Wh9LQ83tAxb
npCWuDvCz2qr00ybetriRdqYduANKJUeRpbEXdb9AvNDw6cRQeS/OezWMD9wWNCH
DyswDt88wDTRevFNGUqcTFkfpxIpFhXfSNOA71qDYbZCl2pMp2CBE/ltUPAm496A
SfxeqxEgKcUtAaP54Gy6Tg2JPRICNchFHgP/osuE1DqNJd+jLO62Jy9uRE+giR/k
bkNmZVoseOtLxHl+Q7CzyurvGU9JwdG4/Xwys6BxuQlD6GBsqyNVPCAiyMMvo1Ly
oiPlpz9tDpeFxaV6p1l4JCW1mOzKOZ8GfJcYdgp+ZwIxue02nAxaZ/ZN8oGwu3IM
No9V30vaJohcCEdhS9/91/V1AFGraCfsa/qG4e0qNJqHIku8iyg2+/gTOrqDyeRO
CG9JA+jCk09QcNwXxlLraFcO+uWnrVwKjI+3Aa/aiI65v7nAWXWNNHGIio1twtG2
FKkvHlmfeRR3xsOcdAgiftWc5Kqop0XuUww0swUaFHcFvg2nhgptMWDwfDfKwRtC
5GgNj0MdkXfGNZQ5vvEVuVT+k5amAH/vKkvzvVEuZi3efX2T/3gz7MPUa82Ic9RU
ajXIEysrrFo8ZhIBiBtj5asEhwpD0dr9uP2i3pMEpR+6yF6cq/Fqp4xeEgnnMlsr
4XFgsxaRNlQk/rW720M8/o3Y5jE0YCgLaLfTb9CoPYKMrD3Ewcsco9jruVaLcpa6
lvkGKBzqupD+a9NVdJDv8z4CUULD19vYHvu+93FcA0oVu1eKvov2k2S3mBkQmJFI
znnKWNmzLLaEXx7mVTpgvfCGrImvD3sxDjveGi1Pzk+dZTNAtG+pJiMjDSG3gKGY
LZJzuuhHLJMuxJdCrHny7kq4U22Hqct4agQOoITVGGrd1OE4N3UXduM7I/de5dyV
vBIP6vVB9FD+cPFKgfW9v7yTzrZkNsu6My+oc4crpx9gvZDR+lUwzmTy7ke7tI6v
erbz4OTlmuqsgKWsWNzawUfpVFDJuppBNn+szAZEgXY4BBeFKonJdOGYFPI3+ssQ
/8wLO0YUA7SFWRsyUfVuJFWMB88OIELJROQYL8N/1RVzrrFlZczZd/benQvmAfjq
6AVjv/4ZkAJZFmsGzHiUuoE9hVt1F0b1kkbjIQtzdP8K72K4Zw28o5XyyAehg6td
kUvKKLl0OMpoMgGQPqx8f2lxLnbYJdUMuqyXQydMMN1KYhY56gL7aFV6UCQyz9JB
ECq2WbjBioyJnJBBz55kqcTEPcInZPExTf2nUYXjrFdE5dc14L9hUk9OHAYxpDHV
8wJi0oAS3WRgbAeLOBM3tPX0QzshzNGTKUeGDK0H/UxIGNocfq6D8mbBuZLA0I+Q
d/M/PszOV+2LRESRNnc5XVh1TIQasKM+bF0QaNsnELvcI90uIbgqgOnBxiGv4/Iw
PhDnlZQSVkJl+YJu/i3iliMydfh6ohNP6wMZhVta3dcmUfHMiCP/DwRuFiLL0SQV
ysu0sXJcI3r9hBz4tucYuw6iRjkj5Aj4xzdN8rhNFmgfBHm/OXOEPtdNTy6SWQJV
goCLaNcb77TW0S9imfF1dpD3nXMbGFqXskqNLDmyYjE=
`protect END_PROTECTED
