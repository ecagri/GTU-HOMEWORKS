`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ERpY8hMTQUN0vTA+cFKzGh1X3sooEdFPV8/kBUHjCMxwq1uZGHaBM7VcZLNQH+il
1naffdVAyvp6HvH0p3gVNYhGj3MbTq0XpA/uS8ixyd0KK+JAI9SdRlBTCNNQ6ka4
5VlFafQYzRDfpdV/5Ki7pA6vORaGivFxz/7vEY0ofqhNSISEGixUIp7deNqGv5XJ
gucC0gbwUTksqaRnD5c6tTJ7yeEKLooua753HTiXtKAESMdzwiqxg+ONjlMm+9nY
tw970KDMvUN6EIbbRywSlCQytvbW5aYGoqYxUBLvJWahUElixwELK6m9Sp7bXNLJ
Ib0bIcw4OfDy5ebEunIj85kLVHmLyeb1cKVPkJ9AQJ/hX94B+OKAGIN/UkXTMgeR
hl1iX9zuGgAAS402bxby/un3kWFb8Ca3j7F4elbuydh41b3ImgOivZ9P8Vh8aKBS
bAGdeQAp9TVI8kbIGOLwa/Wr3QxtO6G5nxtzg3KQ5bsros5gA4W47al5ruYRlSKt
DNTLV78bp67+b6opw1iDweeTYnamkeRVKIo1tLKuez+m/BZVmRcvbJXhEp9PzW0H
2Rkn2dgBwTh8yPNdjA5JLA==
`protect END_PROTECTED
