`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GianacEQybXuENvxKv9PxL+0Gqb2gCIqZrlneXbcrFsPt6aLvr4Jzhmu/C9FJEWh
93bnpKvT7UWh7iFNxEYMiKwundL1I+4uQyq/mpfQNQl4N3DILc3eJ9aTxvwrIZAf
nQNmbnVVisGIP4ldZ+8btMGjkmaO3hCy68qiFKEk62Wil92f/6Pzh+zI0dSSiLeg
9XMg4VbcCBah3h+S5zgZl+QFlmWAsg6Xbpc4OVPs/wMrJfKrbSVUMmETvktsXKxF
j4wFn4Tz6LWjOk9x684X31aIQqFDoYuaYtUs54zXxgB+TwG3FSA7AqUcQVdRdETB
2n/q9dCKOEdMh6L+TsMAoRR5LaqxVxHwZYPvO+occY2kfQl99jk5esq6cGVfUZ13
99vn6djTnvPW5gb3Joe/EUJzW8jvDBXqheMJdNOVWzKkSv0A4kXNEsczkZ1lzRXR
c8JfWLWvLnjZnctxwpVT7XR8nKSRfIb4tBNIimx1urj+X/yazBvx2v3F4BLR7kFb
5OVxpsDBnXe4qf6poGntbtPFXlOdg0JQiZIa/FJfCYk4MEeixUcG/iu0tE3yYpld
7liXBwPuxTjGMbEtIN0eFpljbCN11HckcHieZEl4/AFRLmqvtxywEF/yHdH5Pr9C
ae5NRLDJBA2hbKLoqhr+F5UBY8FpriuWUyuUMLse9qVrw3cw2JtmlzKkvBgpZsb/
zG7S+0Zkbq7lcNRUn7Werdl6eenfl4ucxBvdKyWRuHIRb347hzSL/bjQhJOgc/p1
WTSpvH5nIPVLUqCQ8FnL975ouorgw3iLfrGjacA8tUHESG5oq3eG3j9RXwleVRD0
6V69rLWYm4SwIf+OBsf7oh4OPWrTQqBg/8vLA2hA5HGUnJZag9DN+vQAR9mNAz3R
/9WJM119mVqeexufTf2tmY4XlFkiEAC9YLECVaPypeZAv87c5ZgQuhKBgvQsvGy9
nq2aVT76wgtBU8CuuhLAR9qA0D4W6rtG+gEUh3nT9PM=
`protect END_PROTECTED
