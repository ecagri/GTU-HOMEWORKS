`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
doabQlJKwKckxMR1yIjhpIc39TVBsndV0Cse5NCN5PYjvttM7d3qB4fCQJSHzuKh
Shv4wa5ceSsiQmjezAe+4jIBu2joX0miDIh4IZBQoBfvcMD72osYDwMuXXeAaKyj
+1CG+qkc1tKDd+VPU+LCVbG1whBOELRaYcZypdqhbb6nX4Zsh0oYC6OkPEe/d2pM
hui4QraAPmfi7TkqNJGUtIU263dsdmOK1FmvJ9fkvI7leES5L4V1BSxA/8oeAOBs
VpmSSvd1yjW4PnaTFazCD/yDe0eGdxWoHdl5hGxW9kZs63qqny4MKRbM1oIXND/0
AzY0pX4BrwfMItiJDrIhVc5n/iguhENusZU+Dt/8a75UeNwsrYRwXzX3U54BjmNW
OmtZY99lVgID08NS5PZyq+Trr95vPDkuziCXw/v7RU7v/3oBriuNlDR4hRi54j3D
jNsT6Fn+0IkgLMFQlGvVm7OPzZ1HR/nfNZau9QsJOowtm5nUgBRLDUd5HgrjBNp3
egNm9djbUCH5PmR8aupvVJFlEBYP4aO/H+vh9MQXuaRtGp+k/7EgojQhUJ6kLRKR
MeVAAyKxjmyo0phPYo+S0LjgiYdX4nd1QXc0wxKrEzaX63B29KHgYuEGgfmE1fE8
93sA8gxjgfB1D35U9dnwfGNt8iJgsIeF7nJnqfDp//7vKjUWJyiYfypHRmOn9sdH
15X4OvcARs54vl/IF7/Lub45mYlVBcFWmcg5hthBH/jss9Rdm454hDNLkLN5IFFn
94htIDzoMWId3n8n1V4RZrXATg+dPa0sxSKSk879UmWIyUJYy/WpqwrAkTrhSP5/
GAmJ7Ovd2pKQk9+MKavzLBJC0SncrEgASPEIh+VRYJ6PScQGTpHalsCWCg1yAXP6
SWucKVqstdZ+oEDI0u6yPcXetRkyw/knNnYsHJ2EddR1wdVmbyg9k633Wpjb0KUp
yBuEMQbvQJXxfLZJDH7Jmw915xpMvi0QeoDWrddOmliAVHDfQnEIfpiSWlgDbgcL
4Me4mZ/wtJ7+T9KjIwxe8LLls0cjd1T1Hwa/z0PhR1wkitjyaVyRIInCvuHSEDFu
Ku8n0iqnPqzKNFmH4SZ13I7D2cP837tT1hTkbtozpt6mKZ7khAKYLMzR37bLpjZU
wV8NZiUSrL2tsElEt3gmofamkMw3WSFhidLDDZQsluOdgvTvAXWqVtoCHLISQaMz
wkRdYuhItfBLsyWxZPJxpqJOcxLu/0xrJ6Ds0SnpR0SjY9mf0T12XIU5t0hgXSb6
zeuA+XQJDxNoT+antKgPnnv7WeN2Kbo8/eQs8gRST6sz+6meEBnr6STo0cGvZmOX
AKUKc8NbV+/QI3ryUwxRaV1dvr+/rHB02qjT9ZX8i5v1d/AFlTogLP/j8yXXeCk1
MpL0g0B8bSX4BJSUGl7HLj9802Ka5FsMdXMybmqIWn/BIL63HNq8jbS2GCcX4Hcp
QzLCuUdibRL+sugw0gJ1ZungNveXaIstwDleu1FRT5+2/D1vIZXKwAE9zz9zqfzt
Ojm/MI61CrZJNPLvFhTmf7VF3nPU6yFosy2LNY/Tis5e/0BzkwQg8VDRQLU4Kith
CYKjqJc87FIeXkXNiQuJBl5wkAFZoVQLsYlTYACHS7/s22yzXT/jkAZ2C/NFYnjv
jXWx/hMZHl9nGgINjvXmC56Qh+a3ISQgKsHrbJ8nTutogcJSsBzZYRr0KOnZz+k9
fvVswFbszvQfunLucQCwHyahJMnbsA8tvJStTcFo+46kcrBi67seDRCrZ6CbRxMk
0uwIbIEH1qQMFIiqXxljX5ukHCvhZmPrcgimDGIMUEGjuqJxeFj6t+ZGFEsQKVA2
+Ls7n2vYI3K3RWbuRSbdOssILxQL2Xhu+y4OLIjuuX6jnHQdvyTo4BFq4t36UtZT
NGSenuMhpbHlicPkNmy28YyhL6dWrMaMZRZRnONeepnZi3h/RzVgd5AI/LJ04Ehq
ETFd3BSzdWh99Fl6ZJb5k06clLcu4T1PykdYXynrEPag7zjDzYA/tAq3k1vj9tcq
xoOXYkQHv3UXUXxYkeoBThA/j7oqdU4hkycs1vtfwkunrNyuCjkOwYctBEM8pNjr
6QNwD4ALYvtAdRGhFQzKJSfSU+48tSZ4tkw7j1u/tjGNXA12vaRmc9kn3g6TgOZ/
D6jaw4c590lZFD9bO2s7ttW+ISAf2y9rjLjYEt3dSOnRkL+E/NQmYdRFqlJdDoIm
7TsqYI31MpXHWnCBKaijqTy/4Tk4jBTNJPs0pIbcQNT+DTYgzuQuKC/MqaZv4r4d
bKkt6dznbOj7HzgUZyyVaxZPZta7cAqVng0E5RxgoWTpVmMgIcbN13+r09MmKx0z
oncK5iJibbboFPqpL3FWkV1Qq25HBHmxlVG/K2zyq5bCEycw86zQAtAEG6N2cnLC
DZ2CPxXQHA0GYDcmu061d3TD3aXgVxW9wEy4JO9r5q/7XCLbOQXJqHXh/D/CuEH6
IyhKZx8/zVnZxPrCco6c95SNDDZWcOtQ82yXBH3A4SsPbbJtRlFis0EVw8iDgLaI
Z9fRiit9baccHAi23PVshM8TobmCZezRi7LJosz3B3NcSgphNmdvPJkpBd70Qgf4
P+OoV3VBPsgST1u/OCa5KkOfCJz67teJLB6Ao7ox2HXyEojePg+sGzFXwSRlt3mw
FuuoRJL8yDpKDiBRSINrcZRTlv7+DX0GserrURHhKBu8V1YHxr7GbH8NPzx41uNp
wlfPaCOe2NfM2Nc4/2g1nWv+SY6QUw9yr1+edRMjyQpVnSaeBSaaxrS1jhTJRYk5
o+TvOwu8JrF4p/RJ/X1PaYh214SBI/PHP2FIq26S7GRedEw3lBQIDepTZFXulPVS
jWMO5gxInpDhO4zk6g4Ea+pfk3uLtSOQ+7tkFhwNaGfiQFxzwTwEVhsulPSoLjgB
YlaPx7uj16/6p7WVJiXJJpgyA3C3jbhexWJMpUlkHSdpctq5jV1u7N+vOYzUX4VW
4m4TJBT2u6vpS4LPwZFkZXw58sYSf+Ue2I/T0aNNXBoRdoyzQekffvVT25uDuHHe
294+rupmT3MJ/mBoXCqo9V2ufHa1Fa0alYSoro+/k1fApLwtcficV3uPFqCScN7e
rDt5zOljF5o/GQffmo/svCg7q24EuFIWqKpUZgeNletT507C6YYrbtfW702tzHPC
RiP9nf80pSWYs1Ie6VBmsddftN17Y0nwuuNq8ehl//IbjtsS2B7JU1EGnhO0pGe+
VSBAybldFYLvTx2VWitxXHEcC0too2zByJld8ukINXqIxpUtfO57pQt4xke1J2M6
1Glux5EzchH5Twvt9xqIzeO4EzxxS2kRhouf3LBoo9/rIf1Tvaq0/ydL3gCPQAN6
Ak30ZmXL6DJP9TkHS5Jhk4eNpJXZNgs8idCO12FKP7uSvi1fBR2oL6vA0Z5ZzBsB
kagGn9GnI7014Iy0dTPIs9qTiZrS9+r8BIRUO81Qh7Dt8piLqLRpez6ga9Y5XwsW
ZBsHiE0XsFlKhcR32o6GOBWT+umFRQhH4m1rxbplu/0IMdK6ToapUEuzvNOKUntl
CT/+eXbWqXAf+DZkiGPL8m7zugbIgYnGALucOJixT0oie5G7jhcmchJVCwOHz/ld
YL93kwtzR91GC8nSRveZj7+PRRQCp+iAQXZyCdTgosMnyXJDWqzF+Lwrljb9WfdU
YZTNYEvigZ3+Iwkej5QgeEFEhvJUM75Zl7/iq2NfbGHxed0dP1sMA1nyztbfWOXz
bwjAPmcBK9wu/HDGMENnfoLofJWgp5Gy7DHRm/l7QwXM3l/jOd2QwNf6pNHHx0Md
+1TfjaKyfPHSs/Cztt9uMKo4g1+1rkrkwKyaCUp5ot3PL82pWBUGalUAv/a43j2D
u3DM1SjOwcmCxDaR+c0uZ8ggp1uXRBgagd05uQ79ZB5j0ZpaV9aSTdxf2l4Vj35x
OmEpu2yOSGqbMHeCVLqkqo8OQm7Jl+f5hfxEABrV4hfN6UK/QigaRG7cOE/grn1a
hijgSt7tssSfev64ydeCIUJjbUt85+JyqD6HnryPrWD853ABq904RhFDawCKYap8
BodZ9yHWSi3TVM51WapYR4rq10VPlngDEtYyrb1uWUyDj5PNV8gD6pskfmxdZ93Z
FI22uFfwFWE9iLUgbgt3Bi6bJ3ueXB0hixsnou8dI16X2WQyu9Ghnlvbn4te5/P6
xHG4kP06Rc0BRNRqLNADp3AnBR4XvkWKTiw2us27PQiWuPeDGHqraijerqUFUqq0
0r8HqvJzrB6uFnv0LPH39s8fjF+epButZWlQOqqSLtCFWuqFowbAxRcIit6pikZ+
3TfAcdMco776AlMvwpvUhRLjXiv2yhWqCCmnIZGDEdX8DjDF1q8iGitT3xt3vbiv
fUdV/J5tDPHGuoZuYW6GkkZdKI78UfXVPQja0xdP3ATWHEM5eu8TpD5sFvFFg2HN
SH8Pm+PEVU+dKo0qaq8tG/ZhmsYmUtCN37J8AG70vUb95K2MKzBNNSFvUIUorHVM
Jdt3Y7HWA5Ekw6nkNpazkO3y8PMUbk/QIkrgLBv3Ef2uieFDmN0pjM3FBNrK9PiG
wFuX4WJMUlcGmpR09cUpB0NisMlJfEKn5sWVMtHxpR1/k3Jd1Nqz91BYyfIUZliZ
ShshNM1TRBczpdQnG/MEyoMWe8sWs2ECIdfPquNPCibhXH2sdthGdvMjIKLqwY44
SZc+rTWU6+X2GiUNPEbbB1Y24P8Hst1FnFSrAXz82SRw/NLlogOY6gN15K8DzUyM
a2bjPgJJVgIsTl8nnasGSMXXDHvkht3LPW4GN0WBUySnGQQjBTPG140IidMUeeKf
iovp/VBOGzhLQWqgI9AlJr2Uxc/QxeRNPqlYkQpDEK8QLpaGtvKR4d195DTWa3Yl
kgMCAvgx6joNvVZwf/MzBICtuGw0WBJupZ7krezFynDIvGkvq7cuWLwGFGQWIK5A
z0nZDwHTrcXpeEygb7ap0iwRxC81eDAlBTpf7zIUr3R7/bSTFQA5XClfua1kmwMC
Mdg6jJemohoWTmWntrlnog==
`protect END_PROTECTED
