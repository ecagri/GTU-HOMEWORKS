`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qAXo7PNqvlbt2l+L/Mp3jGMZAhcaAc2nZ7z9t1XVYJrl4Yga6uIu2Z051NCvzKEH
5XU7TGvfTrDiQ/jixLM51kOdbR+zawQHkad/ZbxPlwtZDrL4nrR21E2XwOhWI5gi
5wHvO4Z3/fDUdRtbvuHM627rrc/Ti7hPCYWkIs7j2sLm2bML48DF94pLs79E46qO
OzGtWFIQ0uHKPdr1aonTCPr9EbWeBau5TRK/dy/l6LwlOLFL8Xr7utE3pGakpzw6
GgrYB7gYcEMAVXP0qV7aLdXYaY4yTUz+g210RieiVRlYAdEDeormZsfKFH0feQa8
HVuKmhMyU6BqRAhhLUw9dBZ72/VSgLKjiEB4dbUDDvVZFVOvaTHJMhcsU9vrzFUs
awWSjLgeguhW55eU9OC2ql8yIkPOZGfC03IyqsTf+ugUWtglSvIWwBZRoaNy4pDa
DDr6YhXV3JdRfMkObbRHJ7FLLA7+PKmZtxTZbIxTcr3ZD1BdnGQ2xBgUjWl0kkxj
HdvB+hx6ZHgLdc9MmIxLP8pqa4GCIlEEWjMtmXy+e7ajRd7Tyeq9zbqJWdl6W30i
B96pvfvavzbNxwzyAFqI3tkarUEuV3pWoHAilgmICaTtnvhKWJ5qJsWmIQrUFUPY
LnlW36Xkj2WOiqakuSWwCnjQelJ0RbPkHfYRAx6Oh3nx/CvhkX+WgplC8HnVwM+2
DciAXKa3gV8CQlB0u+1lG8Vdlo4L18YJO7xx5beHwO+rUoUKNwWrEFb+gG+mR/36
UcDWr6Jw3x0BYJywy4s8OA5j+o8kB3o0t4dSIhMxBjEvD0vQENKd57yRjh0yTYQj
fksigH2A06Pt8cp1r+66MqxKQHN4LqKNycuIg6dL0ovuH/BQUiOT7J8I7eJbp2FK
FA24W49aEZ54CZOTYlXbBSmrXyg9wuJbUk6ZzjwgN/50KabaUFcTWbmnpsX09TOJ
mlhZQnvyqFYXi+9GeUDUu32RHGyUxqUx97VgZRfPhCiJfKLUSgrI6P2nh7tR0Jj4
0FJckuC8hqvOSxTVlfiEA5vnB6uVfjbakBVjDcnipbJJzBRtJpebCFsFgYlJleLW
jP8/k9Is3F5Wrxe4s2b/5vkkHfkEIJIa8cmPPd+BtkLAH+lq8QA4t/UtO101Cpfw
V/vwa/Rbrlql2M+CVsUkuUsgsskGS3uK8f/3dK0bbvIrLimpRoJjvO4bCgQOkOsY
Dl1XA3UJSIf56M9Yo1eKmxwqH27cA7NizKR6mEjLD+rQYuA/dK6R5zyJ8Fb1SrmH
t0ELpv2WUkj8tCvRyo821pC5kX4cHguDX8Q7CkxpzQJExGAmD8YdtW3p5wsEDZ31
iEZjrNnmL5Bd3mJmwUjNuEjWMjm5FHH9OSQ4CfQHV+n8g5Xb1uluXETgKiPBFISB
72rHToCDYAD/IkpeNSCbAHcj2Yu7Pjk1EzVgpR3qlsdoTNcEMlG0rSIetPKwVI94
664bz/0Wm/azwczg5ZNDRm6wXSObLBFm13/i8bnPPgc7V+2JtFAyW+Ekrm/epEHZ
ExnxLHRVomioSKfrHu8WBdFkqPxTyqTmQxPq1fZhK5ohw+rJvQSgf9xFTzw9jhYW
nRvk6nnULTtCuJ9XHiSC3wcRCdVq5fXg/9W7TRl2efHKMRhU7BEbbOyXJ0bbYfT9
mjyYE0zFJXST+lAJBQqfqqQoGxl4nfFdTN9UjkO00zzwCfhB7Sjoh9P9AHUWy51O
VuvPiiODhzimIt74LGzHDgDIoHTKuTyTVKQtpGf0UOfu6ODE0c5QnM5W+q4B29ks
ec5W3qr8/FdLIJABiDFEKlKSTIDwluMtDuQsdmgus0LoA2l3zSVO1VsxPLoIW91w
yWrFMNOypEUiHPBjACgbgR0ap2bBHl3ovy6KkQbrY795Y41E4WQm7GMhKNzIWR04
oB9aQVoQ3xlfevEabAmnRNfy+5Imzxg5tbs/CUgVtPatfhO3kIEquKECEAdHC6DH
AkOv0kk9ZSnrFoULXT5MApKJ6Ar321XJvGwyov0pZpq59RJq9Xl7lna/s+yYnKno
hkeXzsY/dnbHDxSIaWdpx0PjeJuGNAl1IEVqtk7HOVQRVBvmO5GydO9MBDY24aoq
HV8kORe+KPb1T3Zh0uwrx5IpHnMIeNp984wc2zMcpvwVFW6PVmGDmk4VTlXnbeGZ
CFQ5ICSZbcU85tUGsYAnk3+KLuv+nJfAcNMXiILSygB0bZ2uUP2H6kmrZmd7zBxq
1fy1APstk6sZd480F/QaZLT0FptIg/GZayVJTV42B0uMpD05NhUo6N6zL0K/qS+0
8CdMbOtzZbBOxWtiYbKFuVzN7xef1LTNsCundTvwmw4HX7Z1sipPms5aGoKuiJeD
HUNBQAGBNM7jJLFo2/lhntTp29lOW3bReYJUxYletaUwbINYDZMYK0JyJ9s5mSuX
aw8lplxB1ylL37rU1hAmvm7E9QF9dUxTAzhY4rL+nQq1pJnHapHUFIDfW+RIO1CB
gzf23IMtCVZuMU5bVsHa23TJqWAlhVA9nS9ew3O5hyVIA9rfFf7Vpo2bSFJJ1F6P
1NCqMzvo/ttxIbp2vWtMTMuRXT82JF9FoOhjgNmZwnjMlMiphx/pS3pND5E9cdA/
Y5Pm48C6HgRZCu3hOdhYkLcCflOileyYQf1RJe0dD0c8sZrGtjkLG0B6qaDT2T+e
2ECv3FbCpbtRTsInMgdO9vkwiqGDJNLvQaDZgfWbmXCFjDr0Kft8KMeoaxymrdao
kzZIFBLnpt2UWOSBxSmK9ZapnlvQC/hOf5O1ZL3DC5ja9uTQpIWLMcs9BLFrpSG8
w3JEbrXzYgX5H/M2Xo4wDLCIARsuN5o8Vbw9WmnzpMN62x3JAD5WceiczuYOfFVT
2GwFv8Oh4LV8JtzHfQL0vY2y9Lea5fPs1AT6kLUqznI5GgiQTiaSsPx4NJZxZHAM
0uAhtmVIPea/2BsomVz7f3fQxZnIIa/XWZew048fuMHV/0Vmj//Y1BOb5F3bQB1b
Dt+nlI8vPs3B0pnhw9Ff6hS+K0UNyu+6CLogCF65n0AOxBuC0HNQmHqq20dfwk8K
HMLf+Je4HygCGzDDgEZ4+deH8JMaobtvJkyMEQ/jsETT4O2G8plYbvyCwV5F4iGg
hzzlNHVhBqiLQAVAgGzCgtC+xB8YEJxfJ3t0/S8N5HtrNZm1oNlvsmu2I9zyKHvZ
bRjWYQcOOAT4PLTnLHpsaK5Bx6qvivKTG5P2I4jLr5zGRlFQ37hqM0Eh3XP+SSHs
CRp3dX0Lg295Szwo0UCX63/shqIXzaOvbEB5YPAbrVFl5DM+bXGme+/cq5C97WWQ
Pc4aTukfRpvNlc+brskPks7RsINw/AZcueB96JSpLJQOHJMOLhuaToroCvG8yoHU
NjlYhbPaULz3djSwWg/C4Qg164ywRb1te+WTDFzk9+ihZIOGcbP1QwpKMIdZZwHG
ABoW89cE9bDct+4r/F1ViN8ou4fccVB0Sf1027vysmJ3CknqqR2+J+fcjldLiGNv
0yv412XlOWZ2GfhMiXnX56VvSfa6NAyRbFP4ztqgC43gU3y/k9Fm4NTd2DEovrZG
HuNqE/bLsxXTE5PQ/Cv2Ui4yvu8bAapAUixwCsE+UB70MsuQuoJOEZ1ZW+5nF9/c
hjCtUEfuyOwX2zXk8i2xKRFSvLs8e7L5ByFUxyx5GOXlCV+9H+hjWadwYMYUJEzD
R52Vzewd0uN7YBQ5a0eO/vktwBckbzQVwvaZwcw8sE5JmkrbzCO0lYIqf5+LJY/N
0g0WO04yysT1/X0Ohyc+njl3CWAvKuOnRkb6dlcQXIS1MAm195oLbVHJk5BB2k1h
imfvKErp+Gtb0D2xqxtkfhYir4VboKCA4z9o2eJ4G1ZvasiN6fsIYcUCZ3N7WhTu
2V7pktWa+Wh37GQff9qsnaI+BLmEcvRrsg6iiEYcxGGlqHOFPn2xvPaE4uAw9sPE
wSQ0p3Dr+KrUip5kcaxSeh/x2Siyu9yxYyon44QdD9JQpK+Aqnwp29nE80ZX9MJD
g9gWt9/UEKGaAtwPB6+/H6jQ+p2OkX+4MShSThsXhxKS1TBS8xAIteUjtOvfs2Tu
u1EHWEZ5f3gENsQOVJ5a2k0UObdmkxB4siML4HPIqXOFZoPFJ4eApRPpmmH5H+Vk
y2sh1qM7rqPalf7SV5HFxDOrfm4GB/77A497PCGfF/MM017NaLnen51ANk0EydY5
j/N6CvKF8LZsvsZ8EhVKy56sj+cKLwMBcFKakNzRz1QY6ieR0NF5DQg5MGzR3/ac
sRBGbRaveXQ2Nb63QaJnPEWrlo8pW19mOLIJK0pYJjRkrfqKmN6tbL5jp6iEhwds
sHb2QxX5Z7tX7o84ZLJTv5p4OArDo5egLCeKuvrEGXTkcJSmnT1ukRQhvz3980Kx
qdLwEAlNTRa6M50v06Oal875H/ILaoywY56KJJJkSGDpnsOAcZnMGWkmieSuo+RB
6KIGJK3kwCZGBo3CjAkPAVshXXdLi65VP3cX2me43HfLdmckgKANSF66CFox++qT
q2RcOGLf8US3ze1Rvx8DOWeQjajOscS1QnCp2POxwUusP0irlYYkGL5rhDZFGkvN
LMeof9XhXl1MQ9Qdo9rfjEeUHbwCa9PSfu3nJ0uR6bxuqXrDFyiuj43XDZ56VKkP
pp6XOGT4oJtVYlMNlCmzguDVv7TZ4Jv1bF9lZKWHsoRF0RJPQ/UztCw/uJ+Z3dmY
mA9MmLh9FHZ0wBZ73AEHqYRajihlJgaf3nBjgrX3HpB5CCy3F8b4fn2nNtk3gmK7
f7sRpAr7Rxj12QxLW9X1KM+qBiu8klcOOBQ8/gBshVpiFP2iky52BUgtLXODKs+c
6xbsdXjnZzX1xEmSlHmaiz6P5f+4dycDVeWWdQOKWNlPfs8IDsvNIcikNq2HTxLs
hHZpBKTYSa8LMX85wit8F8H84tPI/TJWw1LoZ8inoQc9Xwh+K0qEOh5awcgzjaVU
lir4yYEwkpLaCVKSjI9raF+ygtAP4mvplEXZ/wfMN5bzHMmFNjV1gtetvH33oVV5
V/Eboz5Da8rfvOA+Sk6RjLC5eBHieFuemWcTMsdA0i/PRWJCZ5ASQghbNyJvbAq+
H8t1G3ILO9rDHzT65ALZLIS85u5PWMHN75SO/IoeX51pJWi4E8HsZk+1wHa7GzEd
Hz448XM+03GzGW/ZQM3EV4au0zi+Pv/Xc0H/miTCinOc/U+Ni09fFzp6dqksiDTl
sG35QrqH0KaR1KzACsIdWK0NnfRPyehciw4I2y1Y4sjaYv72x3Qa94rJmUGII9Rc
NOSVv32f81VA2098sD6Q4CKm3Kiirj/RsYPv5dq9j24eQw5MpkLNYpFbBYTrQqkS
RT1ScOrSfppJVe/tDEFFX2T5CcJKibrR8XFsEzOn3UQJzP9v8fkABKg8jhh0Mg5t
y7HMUaoGBKbrvmRcHdWFSegezsHF8Yrs8bWXCd6c1OC53u+I7tnB+hLDObkwhvYQ
nILCJjVtNPw9c+UR9rFkpVt6KwT8f/egjaiMxuBV6eI1LDbnen/cYGzcCXFCzD3A
SNwujopTeKcRd3wzp3rDzke48doE+h26RmdUjvHPn170GeB2CRHh+Qwx/Ph2wTmf
Q3OCUuv27BqEXVO9szOj7buMn9AfDmv1UUcHlgS/Q/NeK9whvSitd697/8bcNLOT
pHBItgzJD0oXwgdbDBKUWNgKVkbgO4hI03BtGv2GIOM2DQWPFEn5Rdh3rb9L0d1r
yVG5GG8loeckKco801W7sIRK4J99vXKBeB+Yf2id2jDR4bbXl2PB24X4AmzQtHw0
3+qsQl0it1+12zzKeuFkRPik+YZ2FkQ/8qtYZrudXMpzPpd2iqi7SOse685WyEuz
xkcyUcEVtp6WM0OrdBwh2I3dcfiyMPYntC3lyC182HYBY59mB8n7SSlsP7plCaAg
dZeQ1PGeHF7KG4oIolpKx7Hb/L3cHIfUehmfsEfMt48LHomowp2OsMKOC4cOR5iW
+ywKnR1tZkCMHDApTmEw3x8oK4sYpk+BE97SRPsIcihb0o/qKskg52pLzNJ5KFFV
izIKDvxHKXpEFlBCIGhiTB66MpqyRIoaHPuPWEtqdGC5K6Kn8OW7duyxzoPfjNXE
DR2AD3l1/52CkmtFweaHy4qbo/rBtm7wJFa8Kd5lOg5fBi8mtHfhcwIeFKvMWKoS
audSVLJKk4wmmRCrJc9Q5ItBRJkP4i57GZu3sgeHq5nFUYpKdi6GwKDWdJFFQe05
rlthk3+kiOTLj1b6Bwz4eNxut1KTptYgRqicHpGmWGWZEHIVJ4LZ15riRGPJitea
0c4u8312mI+R20bBdtL2YtcQjVx8cpDn3F2uMw8NDTCcSR4tNNAMzRV54aTeVisQ
ku4AlHkKpO+Zu5NXU7VQWwb4z8UfYjTLlkaGkLXg6c0i2A0be0zPbLHele7jp3U2
1pzj0BXPsu7NehxVHmg5kKw5GYYwf+4krKbdZxqpcpx7YlTUTuic+g5V3vKBS+nW
sNdecKk0pFglM3sRh2ZInhyMPKjG0B9vWLpbDrz4z+5YvWw2WWnaYEdSi45qoRZ5
cfmIrVLwMahzLPjm71lyTz6DcwJ9OY5wGkPGilN3SjQKPmEvArRcLMOx5Mb86nol
J19/P0La1nHU2k6TWhv0zeM8duHXl/z8KcsYzBCdzIRUzia+5UAf6JLzPOomF9XH
fysMR/x6IZ8Y+2tWCoNw60pjC1/DvwdSeqhhL4Opy7m5WbrRw8a93EFDNScr8lBl
d6IaZkTDhDJ1IfDv2L7grk6ge8JCdL9HLcfDCcvJWQVO3+544mGeMV+bkSi24sF9
NLsKeCza9OzE8Vzblgx2EaXz48f2qc6kXM522ENPPtk1aWwTHeoFV/5nkGaV6YcT
TPYToFfZgKdNvpyQAKKasK9JHUe5afZJAnFg7G6TckyaFIkUKKOeX6/e85g1t5eJ
WI9gk0SrC5qMPxwixaKATN7ZGpD25p0ToAkrUGVTDoueOb/HI+r2W4GJzblpCPAN
t81+PDaQbVurNkAE9WqlmNLJRGMDm+eYPX2AyulUoKaFdmeIl9KHE2qQicvrE0Yd
O0yiGsMs+S0TgTY9/5lMVeJReHgdzaSRryCkHdC7xgZRXxBOvBsdXOVA0lj09PMN
2RAjytXIO6V1WkoYNGUUAZ9uh7rkeoffSIW4HjmJjcvMmpvZmCF73hLGgkiEeUXt
ukb3HmXscgZyvIvsoP5AFvI/6FPLgLCHgBarUPKLGypEv8Aiyb0SUqaYDWGRN90u
HFNBeXSFtbYhiRsxR+8cHhsMvIICBtvMvzxvudztk+BksfeM4qDbRnwETGD0E6VF
lR3uPreToECq2vzCJhtN8a/bd9y8ZjAg2aj12JBshQcxTrLOxmf6ZT4tIZhZJdeo
QsTNijTl3pUDXQbgBDW8q8tfZ8ecsLAmVbGqmsESD58W+gpHl1+aXfWvyp8ZRmtY
5M4mnxwSVJ9soMuuM8uDgR6FXVwDcUqerGwnLd1Fr7BAX0vot2koaLa4URD/5Z11
TEJrPPUuIkm7Ia6zaFPP85OVfPvGsvowGTCe49LvwuBGtmBmzURqW5+InTfXLiVj
uQDqyuCtjJ8BJwBJLFlgj5Vb09TFC/jmRHrYzWzuMuDfpmZ4fksqwEvlEYboft4Z
PzWNe19LM0S2hOszICooU5nyCXEAJ2llBZCXLYPI0X6bi3Hc5KmDowEJ45RV6lr4
lcOVjKm9o29RrQ737gHIkDujPvfXQKM6NSzxEaH4MNrAOMFFxngjoKSW7EGRqK+K
TaJcTY9LYfM4OWU7HkropXex4IUpMpn9BkMsjRMpPbtsvmMgi0ZcCHWg+7bxN/+0
VsG2kkTEComHagb0yLcO/Crem6AoGURo04cIGqlSKEogoxyC/sIdxYSk/LXIHqMf
JR5NokT3pq0tcmCKh3rWpz3XESZkawZ3sFGaAMrDHxRiRqjFQ01eL2zAV+FIS/PH
tjrpmp7qaApmhLdstmBlJJXq4c+AdAhjH1ODfsVAReVllF51CRyrfDY9r2jazK5F
iYq93KUwgd3sxm3GPkTQEVr+WZQEJhMFwB2HpQPd1j6y7eQ0fjbEqbiB2V0BE61U
a5R54kAl3H4fa/JCiNgFTXfK27avsodbog9fSgs0jRpiYfh/o/kQzESxkmqsRHwE
AeoCZ03M2RWLecG/ge3A4CvFbdbh4OS0ETEU5FOfQSX7kTeTzvCs3KF6LaSULMkm
6IPEwoSOR9ddFrjM8rzp99K0cSqyLQs2BRBnGooLJF6NtP+0kjDzovuBDkZBfFFd
JAUfdhKYi9Ydx7Z8+JVivP4Yw4ehXPyMFQT/I6QpYKB3EWG/pnkGwn/ftiGrirzG
aUcBMxNqPsFjVJb6DYq/+CeZ6cs67TzULH+D+Z6k4bDPWlF/dLLdMl7JbjM6vGR/
E2qPIQRfhqC927wZg0a+ClAcuwshElrAPz8C1tXIdVztAeJF83+h2D18smIfGbqY
bCh8QdETlB+y7NgMJg7B4PUrt2eGY2PySyNRmAdKqYZClmzSDmvSKuI9RJTD0JVE
+lv5EyI/LW/EjE7PtXyVEeqEsIDYSVOoZQIh8R1QO2yUn+mrANJmda6TocQgXdh/
WPvvmtslbbpGEn6WrAUVXEtlaflH+Iwi7QRtF84g+gxjWgjyR6+TnA+ow+JUMSv/
6dcgTsQIKOnzVmXbOTf8jSddetwFEK+7yj6HGNm7eV+6X0gZZvfQ7oi7/xBIlJna
PTJo2jjECnrBpm1HWOE4bkZAHjNngnTTKTNJLj+gIU0KwIjgx0IxVFJUu7SbbUUy
MH5/nyj1g4Xy64ACWVaOR3vFf8vqmfu9zbtBhnuMyEJOEa7GCeaetcGvH0tSK4x3
y5owfy0oTt+lLXDfD3PRYeKNmUMA0pWW2H+yOw7xxeyh5ifiSqrvXSJnT0DB9sYA
SAbQstCmRl8nCBsyaW3CqDLnWIITxGtfaezFFHx4sr6QpmnNQZy3fBxMUzDvjON5
AetyM47uDE1MoxJNrbOP/0qsn70ijf/kwIQxdomeX2r7K1PriqQ76P0HabJa348d
9D9hol/kpPa6VOGvkr3lbz7lKpKBYFNGuvajA8eogphoAJQMJlwfI61fI70vie0G
QCg148zlI0Mdl48G2BwI4RKURgpOah9rgqdzSJbGQNhdVDOKHvgiUyiAErEXnpF+
nEqSN6l4h18PO/2SkOtcAuaStxFKtWmC4GiQZyhJO/gBkJr6LYbvW54dzTDT0zMu
dQiTGvKRyf5Tz1Q21aUUXfY1dwyu4jQfLOY2tNITZDDtDHE6Kp0mZ+AsPeM4lWOQ
sWLpjqeH+kg6NAJ6ILVOyoLre5XzNTuFTB0MI7yewvOweqzjFw7tAFuMRjEjTYfw
dlMyYgUK/luWsy1fYudts9ufbu4qlbs0/h6LzBS5lz4Myl+9+6Iigfiarwvn5JSa
pvBA8m64dfJmnLbRp9Nb6hndO6Okt1Y21wAtKFek7I+5fwV37gtYs6XbrTtjfByx
VjId2izitxxpJVHQRVui6hYR77ALFrc/vAUudqwMJiM8LWovgswnh1xFhlHdkBd7
/Tlp84X79bGc8S1suubTeh3OAzWL+tSE9FmZI7D13P3DrDoZN1oHklFv6etbICNe
GWjwlG6s9MvfTS95uEBZsZQ/QHNoFFFHDw7cjNkFEPQKaZ49WKblwX+/xCipe8X5
NwohKaaIRbYOwpIIho/Z2bjkig6fcQS5NsSiwiZJCRK6vkDZdU65z2fgSDXfH7bI
st7aXK1pvDNz8wGPE6toSir6zbET7YbCLZn3fZ1YWH2W5MaXor5a0eEZYmPFHh3G
X6ry9NshNyJde4dAOVze3V2Ms+LCRKzH4Z139wFgjm3LqbEe3ZoAgAPjbRi6+4wF
/WEO9brsUhXJ/Em8CJ+D6pYioyufsYNG0AF80rflbgNceROKEQ+D6v7Qqb7mqwHa
FYfe4VXzzWb7ADZrrZA34jrnHCiTCd2R6vnpoYCblocNtHvjmMxo7Q4T3KkXTKoV
LEF95UGbo4VLeOzS/npNqFTJWR2pWIbwYExGLhcKk8kA0GKAWeOYz+At4p3hKA0G
KfnhIFDZ+B6zqb+VWezjHSDEwulC0yfHFL3385qbbrLhZ9JB6EVS/o9sQve77MM/
Z6sTnMnSuwL7nerCAJOvLGWVW+csvwKEHB19GFEaU7IjsB6N/cQKhlRIQeupJ8oL
4/Fr39QDq6QuzWt6Vvs1UH3GW3RXjzOeY5W31mmEl2iGDvlIhuTNLIBFuP+25GGL
50eV5OC/9TzONcWYZr93tXLX5Rt2/pXevPR/USlRhVW+4e7ac76/uB6qcjJCuvcN
mVdxz3InMyEklQJv9//0clNkDymlQ+NrWwg7VvbmAsi51Xf2c+fztr1V6Gdd8I9I
cFg/Eik9iIw6jNOK0NCkXxBvJR061xZ+v5XlvPUefluS9/MGsyOoeuNG+/L5e6tq
OQHpRnpB7bNTB2N4Q/BP49vEvqY4bugDTKH9zbwaAJkOtGLTBqag272F922igIbJ
vmTKl6Jw94sdn+7NLyaX0vhZVjnDFSRIfyuEzbTVgywiSmH+4rvGElKvc0vJWk+z
J2zHkCJQYq7nVw03uCwIop8YxbAuGBX61etbOy7VggVB5rrc0JsYQ7JbDg2YT6FC
6GJn7nbvvzHh6pdLz2uxsJ0HuvmxiS9ELUb92jmmZ0eAJcsnYWM47obh5yRdOS4Q
SnhRNuxF0F91P0I0Yw5g3rg0ljtQ93A2SqjWvzngW3bKCWurbqzZZQsM8P6r9HYH
E2EOTSY4Y9UpFf0egRnuFMnG+60Vs2rPSinaa9FSdiAuxgZRMKFg8c78LwSXXQb9
28vBzrfN+6CrECK6nx1auZRSTefabABiHNuY8gKvxzJwkdlYOuYI8F4GAFOsU79j
/KEnnRGZ8pxUfGB8OCvjRAiJUoCF072DpVhLLY5syueG1WgzCqpaheY8Dlcj0NFW
1KPLHOGnSy6dAcFJYY8/UzLzSlFqQb1ErucHPVFLYDISs6sxASpsuceTI2n2dGh/
fHsEBOSimno7AtzDQCHpEP0O4t2HBU6bYyXhwbKJ0SZ3+TW+f3BW8W/f4zQdASPB
SmkzTStvgzON5YfidrOBlo3xCIdjtUZ0iXlMfrSMwdZvb6k0CZ7/URFWXCpyPum8
ej1X3boYpGj2hYOiyoAN4l8YF0dGeidHOOdzjKUjruyHICLCEiUWQmXPVY3CD86/
yZfUrCV77lwSR3vbKZxfo7rOtyeM7DBZfWzr2QLqyazMCYwAJhkDsMAxV/O/42/L
eIl8f9GE8ETtS2BPxiNtJO1OFgQyYNLDCAK04lJOldR8hpMhmMDWbAg5YGFiMSM+
vY1xqVWAw3zqL9jMOaqxKsESGqQBVGr3gnzNP3VqexbuBI+Pyqg0a4yp5e7LyN1l
HeGtK9YgSe0HzVWLaubQ9gMnFasLh/tftv15mu0JvFIsWibDCbpJ1gcOUeAneghy
OM++ckgxCrUrV9UJBivV8SCO70QrGqXjkNyofu23Lr9/E32T5+BMjFWGRECN3Pi7
rbEUI5XLWij357oUOvrt4apuu/YdFgTXjo5rkhCHlLRjV1uyt8EOq14MuhVXffKI
tcB8DbwEptqQBqv6fS3C1xavDQAdV6YuGPc+6IT1HuRBg2ZSCaKW/6CttXPoHjLA
m9TIWAowqEjDZTyi2UJ5qwzuCd0jHytJq17zhTpf0vO/KZF23wNBlnewhwtthxs3
y3lwI+O3TKsovJdw3eK8d9I6feJn5cSRP51CTL/lyEwTlifabH4wQ3o41B5T+3cC
CSdt9bReZdEOe5ECUuJ1a73JUB2hvQgALLi6psQD7aDAKwuM9UbqPKy8rKGjs1Zh
iy1VbI1+EtvumDuBY0FF/aBTQQ++wzmCgDHvugiBZL3t6UHwF7oiiJTY/jZHnDbU
qE2u3FkbNrDTDRvm96z2iZcq6xLdJcYz2zEgRyasK5LRSmC59Gk8kPfOO/CVOL+0
3Tyj2KQd+taLGBbdv3FuOGf/h2JufB6A/iGhVON2pTtM5MfrsNPvW4cLnK0xc/Dw
a4dHyV7/9InfNb9HfoSkHZhP5PJ8dqS1dQJFucSqdVWApbCAqP3Q8SLztL4Xb/zp
XeRZWgJLvdHOxsd2/lIUoDvH9NJq1BbS1Ju4vSyoWXDHe/ZhLmn3mtrPNBUOOXQr
UzB+QzMC6W7NXw5MmIDGu6BUI7EwtQbmhHZfiTJikW/OoEAebHLd2O0L5OKC5uGn
k7J9bfYd9xYZF5vmMRAMVB9FYGDHM1I/4uMeeCpxfnYkvqNeZU3wa8B8XfuEAKVM
J52G+i8OwNQCRkG3hkqFFWYGZav0MtMJeKcToOFCiu9uvo8VSn5bDLDHEgPbq67n
9FNRFfiHYnd/6yENo5MAoJH0lI/KiiNA4F7qBqLEdFwcP5QHDTZjhUb6P4wwwgce
8tfcdMvpZrnZHUj8ZKvjrfaJoQKJcOXDT61Auf8A2MPUCVEKJEErHjM/mk+/07f/
dBMUljaWQ8aDXyBZWXR5jJ+BnM/3QoMOVtmyLPBeeXSCf7Wh1SXdo5WDk0IIH8Vb
jTYyzUK24jfVED74CDODmt1pRX5MGvwFmp/GcPrxrap/oaybjPjwUuC+G5wW3/Yh
RttSdXHrAo/Eeg9ZJhcBUO+1J5TB3M185JwyZQwPDWuf807XpcbVIhQQcF1+T/ne
i1SlTQKe82pRz25HqwQkHq7kDJlwtMXeygZxiCjZDgyV/TIHXKUVorOvJfh8ysfA
yE7hXnYOGdbNPQEmXSpkDYA4I7TOuYuD6InfYaIWT1FOlYa3C8DXJQkyCD+5bLFD
sp0T66V3RBYq8fbPSZV0wS0JyvxmPo6WppiA/iVYh3w/Fb/HienGBSK4s8sJGHyy
5SBFBdEQMHIli8d+XX7LMXuHcV9aROEVNvl/ELdmlBkkuoHEB7VmjnncvMyL7EuD
bLQY/VBS/ld0f2AYAo31Dn1ce5bvQ9g36ypNhSVfbFqR2mPxmjPVIVGuGRNpTmHR
JKk6b3oe0d2hG2wI8Dl+cq8eTKVYTrcP5XLqYvLobcIJB9LLgtaFV7b+p5+KV7Hx
eOFxBYa+WPSiXBn7EhbRwARp07rwPcavku2H11pEyVfsgY2shvj2yWewXwZR5b5j
pUX4+JapT2MH3hIptjONsMA/ekEABqFOJ/dzlf06u1V2hEOaUEdB/t9GxDhCZ/81
PxZEAyUKP47SAh54GVwzRlqqsM/epgpvmkUT8TsmurCZZm8kQp5iVI1qpxicWEiv
VzS1O1OJ8xMwzPLhur+wDIl9JHuqL0a0vi8IMxcEdQ+nXbS+8J5fmM3p5bLCBtDx
/dqyuAvEhW2GWj+1aTQRCOkJG0Etpkajs1+S8vGe3bQGM7yW/WlP23OLIL+dVBrf
x7ndEt2o/UtA1Dgp4UBxwsZLaBg0sINZAAiBNckTMJ0YQ07QO2oSuZ6QoCZ9fXTp
6hQhOv7IlV1W57xQGdlrjwfiOfXqvKdvfpQJVk4si39SrdOSZbvvwlH5Kxz4QiOv
O7pZzSxkLxxdbldnKwBIv4pc7sPNDVFB4ZieswdD/NkogYocCbGwD+2Mke6GU7rr
Z6UKW0W51t3adYcpCZ+GUPsa+UCT0hNgOPb1/xGHQDgbVRcpZmtvtcVTGvHuOWt5
T5S/vtNKRFcLqWXKukDF2B9cNO/fI2eNXoNTmWd1xmfXcRsHqCGws3kXo8tR/GnM
C80ZxzJCKifUzo9Vz3TUcEgBmaJIGLl/bpVyeN4YKq7YZ9mKQBanwssCtatM3tej
r2WOG8D+45+8Vpd7XM+Hbg==
`protect END_PROTECTED
