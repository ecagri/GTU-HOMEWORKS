`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
844KbQMhRbe9NnFNEzO4w68wfMm9DPSXccNlYtVne6XGHSltLO4P9JD4VfSIbDlK
PWFzXKO1d162e6tDT1oo3Za3NYN16isC+C16YQsPUXbM4yGcwOlF9XoD8JUTPOPG
QnU2oYC5HcoM9NiI8FAFcSYn8aemUa5oHeNumr3MChuyKggih0rCaQIbYWse3HqI
dpNwhj0gJCF6u3yiFlFUjv5Jm8Q/38hqxMYyG87PKedwF/zzHrVtGQ8TIru0iGaW
D4cchJ8yYQ8dAODGLMjHtVS1/Kxa5zo4ld22Kb5EmsRVnBBaKp5JCAdLJpHDCVkf
ITCZq6hXlEXtA3EDF+L5Db9bfkqQ1Rm5k/5TN5TySow8wurfOQp7eI8AulJGg8jE
rwSJHsHb+jr5WfnP2+UOGQBJ+nyVlZS51tRneAG4jNBKjjJb1kCk/B6KzzTARm0+
4RBL4etp8wLZHHHJITrXcCnNCZxFRG1S9SER32VghZOyAgOMfd16X07ZIJ6ts0Eq
NovQI0R0qHPa/cOhbFbQOp9UDbw43Iq+zv7CCP3wA5hmtb35QPXFe47r7jvqArcA
wVyu1DV6bYnwT/RzyET4MX6tYSBRyrKOPxMeDXOk45Kq5cWVU2UlT8vo91ko8LSs
BNONAfzak7vASZ0oXReM8SdYRD+/1aTJmJCAfBEbh+DCfB/yBEcn2twKrTLMTKg6
oV2hC1iqqpGhnYtk/zUmJKKxC/PXvjNEM/OSH6KKEYTAF0prdU9BDnk3kTYyn58I
VGltGB2X7hEP0Bha9InwNIHvY+QbJ8t3fbWM83/58xIY9CkCJP/ijXofPPPAB7kc
trR27YjsoTu+yld57kN3BXsqgKmazE716zD0dnSVFrmcKl48+znjsMYkk8WmW4Gi
xbozyfuu7V5GxCASSvXtpkvqMRT0sR2fFhDmsJBDsXsnEvbmZDIiVHX6EwEjCsFH
bGrD6do6MoqfFrIIGqaR7kSX15ERmbcoXd8gx5cRgI4u3Fm6TeyRiVQGbaXNteec
T/BoiFMTkNmDSDplLYfFJz9yC946yJOtt0YeMJ2OGGOsjyxYyLcJiCK9IGvRxoan
P+WzT7gxwFPZrVcxSlZdDdVvOcpoW0X1QP83dkbpG7vMojB7qxWpTSjfJ+qkQDra
8qCgwONCvhHcoCmasRd1FVmCiR2k9Fy7riDzqCZuU63o4DP+0+/1dr2jbLbaKeQa
vSwRC8rbDfWIRmsaTe5hWtPTKXtNVJgXkMWSNQRZ19WDgGm8UPldzusTvFIhO/Jn
AAvE7XFEzvVAvODnz2pgYqToGcCJ8pv14NZuFU/ASwHrEAKJw0JlFLlffLUigFBf
tY9ZAeQPiQtGJWc3llUgTd7tZea2NiamPF3V/Gvz0vuXPnc7f3s/8kvJLfvFQz1V
/6TgO6KJaS+ygvxzmVCFDkjpJvUdfn0gxoVX757N1PuVq8dtA85XDINHLwxskaKH
8YfMLpg13AgPoQl6aCNM+z/ohE8aUvqDSQ50JspO2l+mHlW/Bcm+29oDNZ12QTu+
w9E7Q3zA0T9i5lXnxP357KJ3a8TwO6iHFFiMdylnIDwpls0NiAg17Pdmm2KHZWRd
1ZG73SzBx7Li18ppNk1agA5R7pldyAsl06fF7y6VSxsvk/h6xnoq5/b4UcFNQCa6
IY1bE+QFg3colRtPC5Fe1FXLno84d6mHQgpmaCJfIX1zbms/jtsYdz11ZbSd9oO9
Kth0TJBiKUM73iKRxEg6/ymbcEWS2XWrBCXEzGFKCtRnm7CcmkKQfl3Zr8TSXhYh
CuIrmuylbx4fAJ3ZYzKIRMj8hpGmlEnPV4mP4D9IPlenT9xjGcqYoYkkaGRgY3xE
uWJIP5UHWfsODtJwJ4b6e90k7QUotH+hcOejVLKRhF/MNdipTeM++8yoRSOrsAna
H/1cW2uY3QPHWmOiJm9UilS8JjYay2PBIR/f+TWkzYepyQJpOIWr4U7wQGb6G9wK
1MypamYTGllADO7bSAZNmxt9n/HEbLwJNJIhdKoNldBg1N5hX84w16mMrWfY6e5V
8jPQ50Dip4w31gdfTPHxYlU85D1istKuf0R3+EocT7mIn0w8CasBdbZeHa9vUC8D
Cur+iqwolXnqBlIvvpT3sk2pjlHCbPBzRiW1OeNnyzd7+jjCOXYzM+bZGQst37Yt
Xzwj4Nwxqc4XRIFYcZwUwVNJw9Wf6wUjjttG2VZgxcIYFYbzILlm1ydeVKNHT5Xy
ZyuMX80trg+YFsDs80vaOjKcM4eNsdOzXHsvY4QZ9sdiONzQeJWew+ncdsTwkLPv
gCto6+W1wnCN3/9dqTV+zS2KLh53vhT6QdYSmkURUju1veMVCz0dDQyUdCl1iklV
Iwzt5+OTDDhz7SUXwLdg+3XW98XFhWWZc2KLgg+iI2a4CResOXmX2o94vygp6hH2
`protect END_PROTECTED
