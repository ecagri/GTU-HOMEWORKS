`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VzdkcgpBuBGxljsl63cSG1ppqYMHfpqA4crb9tx6O0Uz7ml2UrovV/FP4rwArPjf
rLSxBrJsTUjP3nTsvLK8/rPyISZDTKNpEFkfvsT9uedBfLCLgEmxJD2lGpepahpP
HDw8gUTbmZu8w3rIJaCguv3TrPrfWKlf2XgWgpiWGrfjqhh98ma9mpBvEWCEKCbV
a8mwPMBoWY+ZyGu5uyDFwvc/AsUxpeXhNIL9/Zgj0iNm1Thz0lJLcE4NLLFPd10x
VnpBXO5pAml/lMGkTMgw5lc2sChTsVh1hDRj4VrixDj2YtGLTfGH1L1N7yqFyhQ3
iDToM0srw9DYr45D6zY27JCaPE1z7QbB8UwWzN3StLTMsjfWygAtu3XoMAgbBSa/
OeU46UBmD/rdroHNpBAqrPaJGEs3B1X0pxYqomPsVmisEfrp1xokCkRXLpfVbPGe
l3k9a4HyX0BEyLeZRKgtnpPQ6bkgaDHjSiKHjCt0Vtt5VF5lnUCJS2uWJGg5WtFh
WOFgMyhU+Fo8pS5bicpQBbz27ny5Fpg2TWBjPF3n4iVjx22w90AvIU5BVpLOlqS/
PmOkAOdEcTNYA/e3syEIqpNsEfLPonr6801CrzebKXtvyhFbad6sbTjULekn5wxM
yqXnxGXDLci4rZNiTVMWwimQqjpHWvOFmVzArv8dHw94eCWarUXGJNeKqRJUgCZM
92OYHaziAsnM6WCrPsp4rUbw8DisMOgNpQB93B8jGhf9MthYxYgKSWRDguuZZ9tX
Kvd59OAXKnt8A6HMKBeGCrtAuOXW2++4fqf20j83O7G6CuRCcqmv/+NSQXUlDDa6
YomNh3Yzt6UOf+lXwGTVSo4Jkbf52bec7DfDMi53oGATwFpoKwLPKLeTl7B8PVrt
bTSfO7l1pT2dNn0ERODgLO+1v4c0bWhOlvcGSKg0aRAdhMp+fRIEIn+M0hxuvUWv
1JIdw8FAN/hq2kLpeBbuP/leW9pWlrTdbOkCrfzLyjeHCNdZgLNPPRm0rkjj6fkp
BwxkPVTMo3EUnyzqdEPoRUDZ7zBU9YzMD4UG8BJDUWTqoXgE48p9Eiuw+vDj4KLI
YMh18iWQY4GeocAQyMKgWgm5GhH6CM0w1+KTLFQTBQwvbNv2httUIFSZnTHdPCOq
sDtyzGoQ/ZozyVc85i3uMMrSBeSgWU/thbkhP0LWS0NW2iTuWnQzoumznzeA3ln6
4fZj/kCiy5B0N911dE+schOgmNO88uQZ8d96E9rIolbfxA4SBx6+zriM3Yo78biM
BXxYpjA7vynX7nuOGSqw88GBYcmvVYaozxjPD/FxfZWwlM1B+PZdxZOq0VqK2Cd+
OReodJozP8itnsLUECtd/iZOSqxoIwE7ZQJGh1wkL2ZmxubSH9wwNhrz5IayTUJ6
tr0aiuSat5XS8x6z4YBzIkZkQR/CNamUboMZ0qV7qFrpN34f4LGxPB0vbapbiw+8
fvfjeR7BfikMdykWDP0Lnt9RF1+0GSyWIpCvpRBC3EylVE5lfqZxrOwvPmxh+3AI
v0qYX+VNEcfJ9sSqFbl77RE1YS5Ugd6D92EHIfigM9rUQoCZm5zmpnIMRhyEWSh8
iv9o0HwOEOHT4FKaFbbvC+xva9IK4afRANY0/1A1XyZ0+azrbQPll6iLna+UyPtk
COdPMAhxL4i0QX9eO3yVu9v4z+vatlGeSmb+4KX3yLKozg9NfRjIK678F1HcijUk
a1q3yVs9bvAb+TJyDmkHFeoMvkRwT5F+J9YBdHUppqjOSHCRAqEYMLQzVf/e2JEB
ieOjEkNWOzAqegWglXz/uTFnGO4Vbzp4StlE0iFZvEO1PYLHKHrXl3IES4Bh+8X0
lynvjlyJxOa97UR1WgDqdEHfNkNYKarH24xRX5Nt6X6exeF91v6hYgEp/41n9Txd
IR+r86SaaOizKCPnwsI4MXCoULQvJV/NpoxhNxPPj3tMjwPykZd2lexq/6aQM3GN
JTFL/wc4JAkftTt/orIxoe0weA2rg5HpHa+3iI2FtdNBjFn8Z0gk7Mjv2wkkVLC1
Eml6RhDSXKfXdjEejOVCm826nSmUxRDUTEKhgr/rceBILYSs1JmNcKS8mPLPChCA
9m9v0okcymt7SVjgxLJt7VZmAvSoTOWiC+pJB1VcGvIzCi9xFcLxZ3xBoxRFPpPU
WW0FwuUcrlltm4zlIQmhSom+8+Ebuy1sTA2klFsrWQ1t2cl7eir9RWsTARp/Tksn
c1vl8tGI2pyqrbq1JyIgSIy3LTLe9S3wRa8fR4R1NGygLaG/n38u4G/EWeklY3oq
r1bONI9hL/aG8/yR4tFd6PDisSdR9C+lbH8/+E5yO2MQh+kqA+ERAGl+DGlbodMV
6gFbcuzdDPxrmV4b/j7aynA+XP0KzZrjgAtMQQ9JHayfZxTEDMeQWXHgHn5s7JKQ
kvVVik9aVvIflLeRtA1EVVJNn93iZULQujLBswvd0RnytJTR4lMuigH5DM6c56ix
L92yh8L5+Xup3s5cB5r79zC598BV/BTDitcDvPjYOr/TsQ57/DTXdzhloCz3qKNY
UKt7CVWDET8BRvcOF9UEpdT6s1yr/UwoC5WMbxQc8PyeOjw20UkvWVfazwrwpR1V
lJPMAo67d+G7Uar5Je4Tk8/F+m/mSHPDd+J4zGypYZCqFazLdVOk2DJXQw6EQbbQ
UnPY2eYw6uKGhvuCvUTitq3h2tCX9v5xyYkt/gU0sT5XxmZseGhOfWBmqoVxKfyb
AHcPFk/bM0t3nXxLsYZ7NOeqmsoHvN/8csq/zDIkEnTCxXwolre04t101Hle0sVX
s0hf9qJ9CIDkEh0xpGGdYNPW6Y2Ta+jF8ei6S6keHSCc7xxAAESbkU94ae3fGzCm
M49J3QlXCWgl1pywlqc18etfBEqg0m8FJfz+xYT/SbBkHXAVXa5AUy5o3QNaQ688
jcQSmTn1Wd+f5GZbRtqbqoMrcp6TcZo0Po1DsGS6zc/HVvqx3TpH0q19JaLfEdp6
vEk6OJfM5vDA69dlE9p1+hReyWbzY6YE1O5kESY2oNpXnTcUQ71kGliyjjtKi3DJ
AkpZTW54VicQ3WOE/QyoRIBXO9cDX6GY6HF4ZMHNzqppfr20ZsQzGzpxeb6XutLp
5TbKjH1slOLexNixeceUv3Rfo0Hz2kaROpcBBnbUyjk0KkB/+T7jS8W1FZYOFB7A
9M88Y6MB5XmHAhYF3lUEmOLLGOsvb3E5GIT8jsp6rJZpNtTVwCiPFvWIiOx4wXEv
tXDl0GimZfeCqWv38atAWfgbmNRGmzKjMBeJdFrwbP3pT97GmBGZIvsjGa/2Ugxq
/rnVMryxrZRYGlYQ+/lHC/PebuKdoXQm630X2jZmqvQuzTq6P06xKdXmYYh6+et5
WRMflzYcHiRy0J7ugYv6fOIPhpgqQxGe9IVP3dEYpuxfmP4RKveeaDrOb1CPv4mq
8o6zSXkyRc2rh8X52PNEDse0mI0CvE2vcxYEhYIUSd4arOeOajvlLqlkCzZgvjKc
IfKXWg3MJMBxlD0A2EGhdVBmkWeHbG62UPITIe8Lrj6mtl/Y15yImC00sdMaDmy8
0yjlAolM1sGaJBb9wYWLNBuSnPfQvPcJIT5039tvOnUA5GeSfW6mS7qFh6hmRnMa
8IVfXc0249v44DMENMx5P4hMJdz6S+03Z/XZIr8Z9oppral8YBHqQGv6rgNCbRCN
WfNp7KzE7M3Uu5x/29lEPg63F0tSMpaAsozqOABD0cg76PdLZGgUFKB1/ZZkLm17
9i7ZKzVS3Fq8FrYBtza4nb4JrWl3wLcVxhoL1Zv2LWYrOL2qOixC6QHRkHJqLK9B
pUdUSysTwueb9snE5iTiCuBRodQKxTT1UsfbR5KA2aQoH/iD8WAh0aUB1madg8Qq
Qm2ATOy/gAmkgSCvtqpAz+QKjpjU23nfhc3u6IKrGC3Q50iSdMSXWSNWu3T1zo6C
WXOuU60ihXexxYzEG1ALdGX7uMEwIpppmkqJKMd2mMP0gvYPsq4n2aJDgLpruNEc
tft7Q9EVmXvCMexHJYm8t9OyUrDyibeD4yovzTX6xdbSK5OHELsQGXEMj+VM9/x0
xqQJLrd2sEtIqTb5nlQaAl02yyeevXY/jprD7kGFNiAFcAzJYCADAFSbZNEDxVsm
+yre/wLY7AbwaZuZ7am11p8ZC73/3I9KJEU5bNTkjoA2F6hhx8T9RTkg7DE72fst
+ifg4N6+6LViBgEMUCesqn+Os7UcNUvFs460Rn0GOlfxBOc6zyQQ5+TloovozAkV
sj6dkwt8JYAZCyCReT4RvlI1CEPkWAyOeN2tFW6P3RWuDtoF0+/6Q7B9HoBCFJmV
SogwqEIrVw/SjgK3ssGR1mIWEct+b2YQTrdJ+lPQny6/z+P/kQKyt81Yb6Qjea2J
I+XhwNQE0DK7jB/XoBooy8jgn8eKTFh48m05oK2uuiu9rV2TTUh1xztTse1rkuvW
mD8JwTT7cnVayQEkTWs2hR0kWBaVmV0yX5BUYLT/X6r9hGMCJP2LWOgi1mvv1Xcg
9mpa14Mz8yehsDF4QaBHQR3njzEw1O/7NIvNhC+qdKXSEb78gK6EN5PUe0FopWAG
xdwi+YqzDJz9h//Va+BKjzNMXOBdnnN/yEVvEFqAu+bcdaaulYk93915movrKwOS
E3UlDGrKbWMp+gHS4t5wJKVCeVrbDomec6pmW/ikGbN9Za7TZp9ClCK2vkiITpJE
bVfjhOqhgN9y/yqUt1n8uhqQ9vXlAeyhJPQm7rQkoSNXQzFjnr0WoBSBuX/0ugAE
JLb2/boJ6cOCND4tjPLeFgD8QArTNjf300vmgSBsnwSEvHXGN9CXGByPkD/2zgV5
uQxbfMkMJhi4AgHex9fdFAXuqwmA5J02JRfLhHvZ7hGSt47dWJwssXLCtIlZzOy+
ULpt/hluJCsTVDf8SZ+eHqIn+B8yVfhoEvkh6Q6QiN8RVdBMn8jgnNZ2oA0WiEZh
NwVLhHttrpF2BxKqxFGBJfn9dGpZ+eQ5pyR9dbyhSIhDymaFQPTS3zZan9f/xhAc
OVUeE+BPoff9mAtLBUEsew6YISMZ/cC5zI9cpxW5YODOFSUknTz2Ta0SLL3qOW+R
i+x2fF93UE6rINituofZ18ba+yZKjm0zACRXHZj/RMJ6trBBRsp2UCU496f3+Wzx
muPskRAtSw/+Sofwmrt74UgSjji6sopDPI8rJ+Im6rsJ9Kr93vE+7L72sA3yRrN6
cc2L1tDWtFJicIbm9YfyNkPnp8yOLnn33gG/oY/vfNqOWEfMjRnlFEfgeFJQCudp
GDssm/KK4bLuIqWSRWNlh5DzqKk065nIHK40Cb6KRn/AdLc9XmHRu536E62Nw24B
Lt2/HM5RmRUccwrhtFm64g9XwL4ZbjIc1lKVsqxid1khEoQULfq16y60S5SAcY45
VxXjEoGxO7XUKWT9qyex5fouI04yQq2e6YxnrvcVttynSaEIODPWFvQ3+BwcyKwX
+RB5hNdVEjb51YsqENvTrNs1WYQviWyUiTi2VUMsX+PjoC2EGL/5eeVmJ8j/vkaM
SlPJne5Jx1Xn706AqdwCk2BNNX46JvLe5YHpjo8bKURGWb6bMpjdaTaFPPhjsKem
JneVY4gKm6oTdXjTAr2SGunlh+Nw6n85Ee57tCdZINgjM6szYSjBs49E3re4zVCf
0kX3qUFhije/Zy1nV1oVoDCpp7YS1IEosYtYR2G40y+hh+JCHbqfTEasXlZKEqE3
uZKdFVZtLdg7tco4v2vec7d8/YVeDcasRKKmTaZDlHn8KS1qREh5P8ByeouVxVPw
TLbYCDscSZHij6ALGykGKDw+l52WsoE4Ed4/aVMKh3cyT8OUHmQwQviChj7HK9P2
8rjCKlHog0W3DyadRq7iS4bSLAfnCuoi4+gQFilEpelfzucXRNwqSPpyRQtb4TIR
LbpfLeXJcoASvagytFUZxQ92AhKL/3BC4PKx52bs8f4I2BTjm9f/fFN3pl3XTmpP
yj/RhdaMrEfKk6LS+e00WYUsos9oBUcOIWLm+QxCW6WaycP8Ymhbq9GGJR5Rq6S5
t4ihB8o3iaE8+GymmDIlsjvy1M7mWI48b06aAYiIziGF5B095xDI0cyN+mkoryxl
AdfuiNv891U1uiLg2lPlNXEt41AOLmQ0yZZ+zerJPa+ksI63F9LhwuXaaohW8+se
hgMPPjwnHwb2cOrgx4QVv6cex7DxueGb39B8EbG88On1znQeRstIDQdJoxqzTOo8
QEColvrQz6CbAYGcpuKYPyiDW1iEdO8blwOwlmngn3pDk0U6wt3FXaTK2vWyoDKy
M8ZSctEcgw3DRR5HOnfK2sDBjvxg+I9hSOQZayvFlyqBTtApQcLq3sC2dwpn/1I6
KoNDxGedCcpNFGK6hGuPYnfFRKvNWbIG/Nafdh4hvDen7CRLML+bV/bjAdUW8bC4
7B7nL6HxAjjOP2iw033zcpekGdQ2QBXd3ZTG3N4eg9yidkvQsHWU5CJCdBK/Fx+X
V5fdmRHMpCEc25K6o4N3vwcfpWT3Lr+77BnQpZEppLqOW8ux7WtLwasOgRM7SP9z
byJCeiXPJSoIKbmsRPMPtLkB75fyr4PMdz4MnG3tXUJnUi7F2IlhmAgHmxa5oz/u
9KlvSZ8csQik/Rn4kfZvpkqJdRX8K4F+BnTZNKZM30DJXbLGxPcfpd0S1zgvSCoR
IdEnp+Q9ulmz5g7w7rzJXZ8lYdQFU7UrD5Aor/dHd1PswSHZE55VyCl1wmJA7r94
nsKT/JzQVHeIM+QoY/07M+Pj5lleW42g7owHdM3zBhf0/VdvkRC/DAuKsYSkqUJX
PspKfaq63XuylJ3GOUVxyWrFYJ+FbQS7xeD+cbgco3SqA1x4Z0jxGpQjJGeGYTaH
NUPbefp6wxozWtpPQCq67ZVtTuHj46Kowb6GYNS+QI7pQQPi3b27HiO5ZTOPWu2k
C3VQTDeEAxKpbYsSvgi3WR9w/uZ9khZ51pIEumMabePmrCluMIEN6QHmk0E8wu8G
6WtiNhvrSclqrficlv7yii7Xsxp/6dvgPf7E5369OHmRKknAejjpggM8OfAF436G
8x501RgqsGlV3TVky+9+2xwclzovVrDiPyCf7QdfucgS5CG/NNraVMjvvqGpWzZC
nkTip73Qwle8Tn1rnKOZs0CyO1FNqyZpFZWE3hWx0ce33JwKby+cCl6A3lRmECKC
R8xXiTxQGx4A08rhI0kyrHMtQjelTvryum6uJzisnbCBnGHvpjUO4mUW6WB5Qakr
2cglP1srOc1Kz4F5BqWZ+t50Cwy6jsfqUVVrYu2On0mUkT+oGrSogGEjkIJYcsCh
69A/TokVlAbuQeGHCFHydsZspd8hACYgK93fysqDQCdQ9TEGE/Uon6qcx6jF++Wb
Dw6sCcdRtEjZdPFFuTOqLg==
`protect END_PROTECTED
