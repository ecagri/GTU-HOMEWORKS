`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5pd+iOZ5qzVM+iMqMoH6zRWDW86fiddGGeggPxLj24sj6yiUVe8rxj/aRmol9jJf
bku73hasYo2zfKOrqO51bukfjl57h0Rupyua0A7Wvl3jLhruAAGREsXzvSjUiEis
cBv42o1Bi3zx/vJCD0FVoayqeFusrcm1zIQAZEOAZwSPCzGJZWn7b4Rl0FvI+1R2
wWcmSQZby1ewQ5xtQGM1HCmns3Lx4BpHc4CwXmWGnmqpOTduwCXWEH7j21eb54xZ
mrd/n9Nr/jlrL9/wSSVwQkNd1d7LqFjBv0F/UvwPT21cHg041eG4BbnXUpVn3XMf
kNIwe72vWLwH46naxECzN4JGU8DxkP8h1Mz+z3+yv1uynts5o3NqAZNnksmIJk0w
OSu3kqzLUi1mkRJLS/iBv1Rk3n38AUDNNNbMEd7d1KPI/XA49JLW9ke2Kh9Gck8G
X1h4Ht2gMxH1WiL6PWSCe69V8QKOHICkLQv2zmep4aKB4qXD5iluqYLxbikZByTZ
2FdgD++Un3qb6OcoewkPd1p7oMqddBIRMl4yBOYwG3LTGdmXAjC7LzwjXZlu+Ziy
zQC4UYoScxe1OwL9c/pNcMD0RMpofPzYCw8XPvQb0PYoAHFx4GYrdJ4sB9gpxZ54
zZk/H5bd83ZmAI41bzFNsXCNwat8nCp/wdg8imFR5HLfGsXrbWldR1Jl/mIY/i60
jd/kOHlc9TemF7c8OPBYdVa6pbutxpgz1dnJRfO05F0tRBeTZ8+cF2qhzwKXXi1N
ISBO/V3LHk626LeeuUOROyj4HJtutnpbV2fAkS8GoI2Y6XJSo+7m+PDwSyBRbGxp
wWDvlalaFyEtCR7/8rlZ9PZJvAymggpcmFmaitku2d3qlffty+ZgILeV4mxKdtLN
+IDubDQiNmvx3+0gJDYysH73Ux5o60ALYC4JsCitgOOcLKUss9yjMcNCOnHBClXD
ckmusZyuBTpRlEq3IiI9NCZNFuZMyCX1yad6JMG3+sU5NkDwRGKGmBxbm/uyCkx4
5Wx3AL88T+KeKzLgj36wNC6UYM39njF0kFJX5Fr0SbSePAzSEJDetEj2w0gu+v5o
GZb1KhTGUOgy42gG9PITYItDrOEPPtbPw60mHaixysKIPTTtHiSZ1cECLtzFoWSQ
L7oEFxiPJC3I7AKk5ToyT/WYvl3LMOxmS2u2BnEofswPJAOtWojJIgyLql4SdgAp
HdKQAQvPqzkzSfP+cTSo0p9Kfz20S40II2kz6p316ScCSWO3MJuNjAlYyQhjaArM
JqSptmqRe+gecb44+cJBCLWmJBJQ9yjwlK02vOeNWgWpekNr7ERtmZgbeT/yfSOE
QQQiFKBOX40xFE1Se2lqxFjsXPbS50MeFmfBv2hQZQhvWVCcYOGBK6um/ftHsAUZ
yPypdAiYmwxJMM7bM5sT0XnnM8tqx5zAleHl6uAOj025CcwvjcG5tBPlwF6vEQGf
inVSHY+ASviCfcDO5mPi0AsluXo1Ygjg+XrJdF+zcoOV1IlBAZXl5M3oe/R7/mAz
nf++Uct7fRXaNSTuqXYzGKHGHzDRI145F2n8WlbaqRec/l0Y+LgFG1OFxd+BYsMH
vvyBV/0u6bWNXEwWBvCKiJD1lQMcEillTABLlvrfs+uFO1M4b8iMnPyCOTX0cA4V
0+Xcp8m3iPNgTETZdhlGAO27LYlH0g9oWrcMks9DhK2bmuO2GhBlzLs2MqOp62ZP
0V+RwdryaJLOohenwHZ4G7BWxI5s47gyHdFJGerLjQf20bLnaDsdyOnx+vQyEtON
ExNp3k6Vvtn90rLKYP0PRrjgwkiiCaDY3FJJ0mFW1s2uhZlU4xUGmm7SD4IauYEI
YNE+doybU/swkaDMJKD37c8FsFRRwkL822nJyY1f6XekK0u2RKkfRX9gs/rtgJVW
yuSU93hv9EDx6FHKmq698C1MHIsGfNK28a99JVCTZJlNGEa9e1t8+ApqcByXC+xb
7KnMvJUQIPUUE17WwwMWwCm3COly0Z2a/hs6154EXri1Qx+1Rjyq9Esm73Xy4kx0
SXwYr2uo4U9tSRKVv9tc5F+vdlWjK0bF1jHcm9v73V3J+GJAh9GH0O8ZFHKUvXsj
6IFujOLHKF0RU76rM6fZFnxNqot4GyoDrEwdZ8I1r8kdYkWHLGVAEHYcl4LiEcjt
QV1HYDMwc2X7cFXxd38AHm1aMhNLmYvKpauVYMNvJtui4s9u65vnsDTnRYEdMvEJ
m4u/lRJXd6Huuwn4muvzxX6Bxco5KSw8riIQuyCyApU3iUrRQy/RtYHRB6aI10nM
Yphsx6lGQtrD8nYypWw+42QABYDfGYM2PmfO5pYSEphfHk7aJ/Zt0Wx9WAarIhto
iffTA9erL4XRJrX5h81avhr9rXJjDNYOKyyOPyz9I2CZGTYK2XEQn66uWzx6A97k
weaBnwiDhyUwwGglXlr9i9yILA3BQeUBa199wPFwe+tgFZaBkCKhGCv3oAm0zkbq
pFJV9Jw6QzP1+tAFIGn6qukbM6zKObzUyub8RbxlP65I63ZS0OmFmCUXsILLV1Zf
KrhEy4IhWjw0nU3ZxhVVmd/U0p0DPn1ubbXU/kHwvPtpkj925674NxMHfIfb2Cpc
nbqrqBs2SHjOgmDyGZGI3K7J0iUIhsMLL8FZmue0JwSkDA3GOlBxpa8uz8AFcolO
vOhjDRlFnMvfKmRhr9oBQgX++N5onW6aSAlTdxExgs3NHEys4Zmdl6SBAk1AUcJL
A9nibCNoiUwnPkHJ7jdUMI1X/9x/aUcSYwWqEafuAjjPNqkWfM7Le/SkVDGNksCI
vphiDhCblg9Mnnb7Rz7NO0fDK7W0buF3gJ+ojrFdJNl/QU/fxFxreQinoIi4cplx
HAGXtF/PLlzpBxf5XsllEeMvez710AEyPdar+oiiXwtcYKhJAuJDE0p14oLeD4kL
CqKaouwyHzzSMTYHgM5xHWO7lEIUseAzDJPCk3unEGY+r1P3fUxyEkHZzMwFwoRW
uajEmd2HcKeWusNTatsP0QHUhFkSpaxvEyxuj7NFeN7WqYS9HINs0SzMneFkAQzp
I1Q/CSzdvjkFTTFL0Dh1VUCFZFPZMW4hZEQ3cOcuQebWOAmCg46w8JsemFJv2WXv
EGC/n6/Pgd1mh7bM+niPj656xdXfxH9F3eKd6y+XSxoygEIx8R5DSWuTkmsGDD6P
7bVrMUHg+XduB2gxOloEccB4Q3Ew3GkxobGpogz85KS5uKVomlcbTZ/t1Ma2Y/vd
l8HtlmiPmAsckpSWO+qxEcTEvJFbWZ1vFivRHmzZEJgq+W8yhfdVX2ktPeT/8+YM
PHt5Xb2mfYqsD4CcXt2ifywdJc9kxLJlH03zHzd65cdQBUBqJNaQbw+aG1qpYl0a
6zBW/9D6OJG+J/oLfB09gYGtLS1lxo8jBEfkayvE0t6lE1w9w/MG4C7+El7R6ebB
6EHpSqAkd9g/VwzxarzoK1dRy7BPWeK8bzYA1YGzMrCzsSzzYyFE1J4Dxm1Rii/L
jjr+1dnIiw0HBN6ORTl/6RR+f8melzP4DPnibUc0Xc5omVAEZDDf9g1fYjKIzAdy
hPTQdjHySYyj+/HKtIJ94I5JfGBcAN4tT7qw3QQGaqq5EUYzhukbVyGoVCWM3cv7
vom84OMl7RHa6I13xbl73VoKJbPKvdmE/tfvqgynPNSA6tIH/Hx4jvrk0tN7YU6q
1BymjyOyDo4GzkzKDtxNvX9DSGpzQk2OAnTbicWr2H6F/MqPUE1FuHnmkZoEkt14
TQtapFifarDHwcKnsfDkFfxkW2zn+svpk7XSHqC9R5HE0m3CZfYleStJPd9sXJkJ
p1tGT9FfR95EJcAJL9kqMUNnEPlX3k9qTIjU12LyR5Csx9zn5bwRauhUGbMBJT3h
9KlQvKy7783T5kHkZ41FIi+xK32LzLUb2NAna2ot9scReOnHLLFSti6Ygjba+O0d
WT9M/4bSgjcy0lQPcufcLL+A+Oaf3zMtvZABb7emOpSNwWxN5MtZH18+9Zbp9Lsa
rcID/ilJ2JM+5CkG7z3UsNCq1VMOJE0NJP108XmKO+BVMUSPMHVA2NDpmzTqZG8D
Qii4o4XbHosgNpl2MNlhVR+2owfqSWs3zRNkjnnhM2VvUqSPvYXU7YrUxPwx/Pf+
tE3SQuDHEQQ9TsiH/fmi2p0mt81EPHlmSCjRd9lBx8nA02Taa4Ms7owVCQD1NBhf
dnwLw9pqnw8sUxdH3BCCifmjQ3XWh+36E3EgyJwXkU8zeMjpaSBqibxvnH6NfHUb
UuK4D/Qfuql92kU1R0yV7z+Kzbcp8KigyJ77k15OxqXgNEEZy0ID/wi/mBl6lrog
JkxDQWtaqNB18GhmhWf7jlPNU/xauto3glt8xgeDfB6Va9Xr7LHIAMSGxX6rSyjQ
MMYDFCXqOu+7pB8fpEufhmpBF04RWBFkodgX4PE/Qw3zCHadGo80kbG+6rboZE0H
kxu5lN6t0AQoHyN4/tQBZ8CvuaaFtuLLhXJ3mIkGvvG1PIZ4hn9YtZh6H856u88m
qXadY+QQi65CWbZOEXoUXDFdX2EpNO2NBSG7+uoH54k/y0l1NWbvJ9swHYwTjPyS
NuNS+5ejitc5YIGKXkjBjJG4qQ6Z3IUSmI4RnyO1rnTciN0wSnZ0/CZjO/RwYGuk
xPHaerXknNcmrJmLPG9NVnvCFq+238hFGx2P8ipAAZ5cNjVLC35QkSq7SIb2r8H4
xuMDUtdCJ2of9R1AxjH2T94043wx561OG7gi2rs4tfE2SOgXjAD1JjlJcNPd5kHy
1HxLtSjdN25cwGZebw/3OwXcSY/ehYdaHzzUkXawobGwCuANQDQFiDgqgn+5h/fc
y48x9jJExyow5JzWYnOLwLeQwbGyizOdEcg+XZTS63uTXifk5h8LbkGQFOBQoJK8
pGhjJJjDwloemHLA4XhGfDcrY/RN26sCFksJeYZkyzMSRD6PjZWkYMe2cBB0CRd4
1+2JuX1xvl28cno2oKv2i9nXEMp2AZFuqTuMOsc7p018eaeORCbBnqJwTMJq7934
2B9VxS/+uvbK7Vtqaz4OdmXCu+SOXh/agzqLvCl960m42lNyzlmZUiHFjF7kMvIW
vJPA7wxtUgEfkQwUTw4oaXXdokwygat6gGkAmSF0mwr90Reiqp0BuyxGVMFilXpV
Hi8daQpqN1yUFPWfNq4twNcwtiwHKS9Hn7lLT7eG5qrNfC3cpmpwPrTMkZT++xFl
ZMkgklf11SrNCZi38rdSJbvezXBNd9+FnuR6Bu82Yt1ZAsTnBaw3Jn3LhZsQ8M4H
R8nKx9gc4tgzOjNduX5iQlisXqr4Y2u7Xvo0ULZcLLOTo8TSF8ZJCthuLk+8tlhx
8G6q7IqIh8YFe6+ijRpF9HxkVS+x630Kzzid7bOaHce1dsey/gftWFQw4hx7eGVv
9ZMak2kfMSdzkEOlpzur2b26goXSlR8wx+FXhxuUlVkQvSG3D7G2Msov+f5B0viR
hKYJYc6yaW7aRL0pmYUMKCy4ritFbRKLINgd4Dn7Ywf1LXTiWEPzt2TF94LAayyV
li4gkN9gPDdjKVEkQ3bLv87O/ipYuP+o4m4SbFHXbbE7iTWGQ47GvFrnBpuTbax4
PFoRA+bJ6HqR5uT5a0MKF6lcQX91PRFLn/W/FbRE7CoDURdb4bs8nG31JiKJ7yC7
2Nane52GL7ZoqobS3L/y9FJ3uO382MfP3A26K98TxqiQH9h5+6Dm76EHUfK/jdNy
FtmFQo6hNp9rByXKyK2Yay5LTSepqhdTaILBWMxolvdzW60WrSn/zMUZLUrMyZC+
TE8GVXX5TyjN3S9UG8+JpFdPYHzcAawNVaijbZlD5dOcMmgbgriwiFPzjm7nRV+Z
iOqUN0gyvoBJmxg9rkuk8LvCpvk0uIKWK7PDvNgXgc+GbISCxNm8wgqMBqnsbgUW
5BxfbuCI58hDIios6Ed0VWZ7Gq8xbjThfwvw6+oWsmtZNHse5YJrVxrV9wjve2fv
pGQeJKmP8tA4c40O7NkJowRKbumBlWfnBbsRa6++GCt9n1Q2W6M4AP5oiRR7WbzB
XF7TFpBTHuFh5k6RJFNg65dSQM6Bm1E+aEdE9NcoXwP9tcU/PFtLtO1yng+N1vDd
l5dVTO328UTdMNM9SwzvKJ9tkG/GPRZ7oBne8qMZrfthNHnMiTBfL4MJPhz4iv55
cDzSokmw7GmeSWZcLuIqHdHMqdCJenjvxsYcfVgBJ0Gp5KstZa9aMkBTuItaeGFx
aUTynKe0O4ZwFE/t3KASICbvov1+Y4Ww3CAs0+ZmvTWQ8eaHt1axs2cI0x20gB51
YwBNPuVvXSpEmSI2LbNIwgQcfIn90xO05FBlNhk0I2fyxlLgq9DNWfMFEPhOSn+X
im1RC7VBjpg8Mq32v7FXtID8KDF2v6coLUwrz/SfNM9h7DSlauiJN18FeOqFlN3z
868Ihehuu2sUml5fp4ITtzRqjooj4moNlpclbTj6u1usrYxksfcDemLzoGtJvC/4
yjLKtIBTX84fOXTPtpqPDzKhmXs3rGAhGCf6Ma9r+m6fE+tINFdYwrPtkjg3a80O
MOdSXAlWcYAFXO6dNAGr11g6r01D33xGYsnvZVIuNmodPcK4chV6uLi8/jufqwvN
jS5sG9tXRdLacG4UYVAnQD10MiGNgQ6bUpmXF4VD1ei4L6YpvPy75zN8Hcqx+gPQ
rK4cRs9Ng9xb+s7jwh+ohHBuaLvoS9ref3jMsAzoubst5gtCVUCXDCHMkVAmea8M
vkfWSK7FU8UUv6uMOu4IhcOzrYscpoStksK243rqD3wrH/WA4DO302dXnzLSUU0Y
CQe1+SysIgmf34N8WBAFwXXaPgGz79V7toH8jTz144b7MNhn/fa7nknUHajEJcwo
NXCsgNVEnsc3HjgYhNi/fIMZwV8xJ5o93E8mkioZ6hE2q2a17UDlhffS1lGSLbtE
K0Y/NzRbAYiiLLSfx7FXBmhFZZ2dVo0G35o9MmJZ0mNhQLJDWAXSljcD/XWgwDXc
+tSW3Vyux/L6VOaYP1kkUT+rsvBkz4sSHmPyy2qXOgEyk7IQxpj/L0ZPgBwfIzPK
LvC7ZQZwp0REzCjFl5fd4Ha3HqZW/lrVV1nnwC/OkdhK8L8xCNYY8II+nUTdS/Aq
eJjGDvleXYJmPgr2rRKghg8DeGtJr+wmMktWPgelh7PGtgqCWCS1OEGB9sOZtEEz
aemaJGQgMQaHDV5/ECCu6JLW16enWBy2w/G2/SXmPgQnVjsgfuO7LO0Vq+WFLO7v
npcTCfyrJZZu5jzCOGALWiqgAfL+/LzO7hzetuJnJ0atgywabAyfpBKECmJGXg15
+phbB280jKMH7Mqj7ePZDV0I5+clp/rP82vXOE3+QfiteJLnSuOuBK6ATk8fQhss
n2YVCZ9kh+FvKLnySy8LK9XNIcGvymWJImh7JJGL5YQnjNab+I8ykaS1XPm6aaC6
i+rLyeLASgmaASpGXDJ9b7Fnm228P1QiFau5A4UN1dxQaTnq/rszQRqBR3wqxvq+
8cJcYkD0SR4N4Kti/mn+8sunQq8oerl6B8Md9KuZXeNsPJlc3FIRxNTKEviQu060
xQdCfnSKpg3MuVUMZPHsAc7mQoA5LsOvMb+mgnQ4IOSXVxyviEPiyYWb9s+ei7TA
1kE2EDk04K14sBfSRzK43JA6sE4hQDqrOZGypAPKFYC3ykeOID36QrSIeu3Do/qi
0h+5ySzaYxjRJf9hXJAAMT2vt7idUdmUkF8CWj0r+59Z/fmQ58TWzC7EUoSXOZux
LMPsS1/KG/nEqQ+eerJqKgUttWoJM0fU9HiEfKeRD1MxnenyQgzHR5FyaG87j8QE
KwYPQr586hmBrwMKWp3KwJ9C7PZl0jFk52YMkPoYBs+IpfPtEHnQ+UMTU3s2GylP
Xx022h3WHqX16ElnAl6klV08l3nl81n75naUqEXAiHSJTDPRjLg4WK89Ddo9D4VT
jr2t6yO9SLIZoS2kQkLsa4osAjIdXetVyL1fqlRzAxv49CXu2zH+EJdxsdQZl5KR
gt+9eG+PRa1tXiCPM6lO/FKhiYDOatC3ibnHTLxwcGL6kE2LmST68Tgozl4eEQzf
hKbMf/NrPJkD0ScU1ezAZf4IQzyCJ4ZHsVWKTQpFWz+2Fr/zz6NICFMk1BydPrfG
Y3wGmOEfGQpphyMKUIB/pD3SkFV0N+uGh30D9ZfSJpd2/7oxtM9l+IRDjOsV3LWz
kvrh/ZJgcZhVzObxKQLQ2ZCPuYBPh9c5cpwCqQtTz6wA9BGhb0QrlH7A78x/Kal6
N+lGjQp02SK40Hsi07LgQPtpV3ymQKtHnFL5FgXgnp9QPG3bS0oZcIe3xvQUUrQw
L/M7kkBepyYN/LdZP+Di+XtapWsGpOrmcwzQD1sxfWOJ40OQTgitwiQig6grIRi1
gbjGO/f0PAMMaL+7KF4DEWGvJJOOkiSPp8h7vAhraqu9c245jF6BQTOWf7IUa0Rn
hRh8mXLodD33P2kxC4fcv3Tl2CoeRvcneiM6tNJM/H9tItRM8b2Iluh3iHy7vtdF
l0VrWLGjP/QXHjpcC+OAw6LwUbWQunbnQ4NQjlgRq7ZVPlUw+nyOdhYuniBDEupF
J7UIcXfLkesloxuPdI1NU+uQ2Xkcf41Mb+td83mHEmjCep+18z96HajdsZTEjv64
UbLGferqV/mAaVxy4bQhyya1XKMhx/kC722AHXQArFwXwSt2jHS6bEaaeHa+PnoW
q5oNAvgpLcqrIca2PJMtgfLgjwXtaRb0DHR3DIWXwsDRZpgE2RwfaPAAnYkWcEJq
PoEMrag6FBHvy2/GtHNHtsPfjaBJwurQRw1RdSBnaK2SUUE0QWmQ6JfNzQkTadqZ
kSCEmjuER0ClP3v4d8BypiPqX0/zN6Yy7gzoBa6hApuugrTUjaTZUGnAFXumCvym
Ojxo1FfUBosiHsS226RtZ/mc8dnagsxGapf/G4rj1Ja0V+BHWZB9V/xoniosH7oP
6QM3wdutFPsecIatLRZSC6gzouBomj3uGI9HPfNBBLYe0fm+K2PMc7u11Yh7abe3
w9XBD3iQUdZAxdat17Jy6j0nnJbQN13Wzt23UXFegNgfKEvDq3TCEeXPbp9mMEmW
jrK6SNVBUmPLqq4MQ0wDjmzsTovutYB8RJxBcxuXvckiD78hAaX4mUjDplAra6Cq
e4/7qRD0kp8bw3mqih2H7eXuIhXe5ePUx6p+DBLwwvkDjPq0RM76JuqYe7EDUJNl
mFLwV77rfqTbiqSz1sCD8SrZwGmUlzKMrdKyeuXhCEjigUr1rtEKW0VrseQJ+Zfs
zuO54qlXHb2TwXYQeIC4n+GgqcT5m2Z2tEI7adefay7bteSy7SEV7ZX9I9H7w0t7
+/ExLjA8Z6l7ugKBIK/JLyHfQ+sJ4nQV9CpeOQIlF6ow+RT2FVhymdmRvxbAp2u4
`protect END_PROTECTED
