`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SCl5upKHkoqZBxE2o1Oq4Fe/5J3kvBdxRi6zzWYpiNEYDrKy5jwKo6p21kxsIjnJ
UuEzXsa7mF7Df5rS1REk/IBDHFM1wPar0Gw5g3osuuG7tGeKnbi2+kc/CZNl9Ktl
HoZZT5q8pssPGUAegY5zjx255QqfgDR+01ZjLiewziadyaLcZrmuDqbVjkqJMQi7
qB+5KtQTl7xp2EUNk9WhFKAYgZ/DAch1uQmu1Hl+nwfNaQI3IQdxsU4nzPE9naqx
dq/EFDDEyL7SlFsiOYu6HjwwGXwkwpan3v1LV0SSooymFqWwBnt9AaTuLYCu76JO
HARZXcUsBuLL3fic9CQ03ZyB0xIdKlQSpwZ5b2aXJMFqK+ATJRndBRKSJqMfi1CG
FJ0xSaBmEW8zoRAQDckmaaU8iCgIureGROgEMTKZrpvZIR5awAEU8Eqt+4jCiggM
fdYtiCIfMMo6LL9ty87Dt7J3i8VTyF10JEme1IWrVN/r8++lWUp2KuIEBuEbVgpu
hTqavjcBfNCkk2+KCG8PJbJNn1RdaiHosmbMadKFG6pr17RAF16xFVnCx4wTLE7M
PS8ws22PR1yBnkzPwTYLRc+/RWQw9EiK+SCdHBafIFlTIAQYQUSqyoVThzNVHlTi
6sHMRC+24miLeLrTf7JR4VQmN2Xo9qsemQGWgTrMfSRekQQky3w2DzC9rXP9Ay4v
ZAmEnB1zoeY74cUejMpRzNNEGR85F8XkVsByOSZcK3f+34j0080Cp6YqlcP3yeyu
0O4bBVztEMPOfrOjj/Q/bW5XEPPSRXzH/lDG8tlgI01b7ggZfIc/sc0uUhfwIUyo
XW6LYZz81N+qQ7n+nmDX0bDH/q5kYlm8ZYhWbxKnuxgtPA19GtJ6sgOv0Nj4mlXd
IsLCUB1zsgh1f7qI0uHEz1hd00UUItHtxMXYdta9zQvsi8X9wHtc45M2wWxYbwid
aPaRxu9A/V7iKfLL9MNaBsaKx3qVPJ1SGx8IZrG9nimDJSVVYFNIfFp1Q4Z8Kgd8
IqSLmTSXDFYOfVjtJ5rFlcvnfAR0j6hVExVGcmADMOVsuubGiN45psUQbaX2RXkU
cDXJlJpe0bl5wZOsn25TWqlkdwKVlxp+mJIcCUR6HtuCoFeKsNf4u4yaBRYshJQs
7JLea5QrpxN1ysWpuHmEsfUREiRQ/SoKA1OqDHA2cPq1ADOjPtiu+hUmyENR3VFK
bxnyvf1nrTU6MyNhdt1t77ljdanVSwCK1I6jS6Rb7eYw9cSwChv5w4H3mmZTSwVi
hgQbGxnC8ZFdyx3RgrEfuyuQ1BpfdUanlwGBTgwjclMfaBBvKJR8p4whypZ/urLS
++JAf5o30bF2N0qxc8OURUvqaOSAlZ5cYU9gmya1uGU0LurgrutAdmAJAMTLOsh1
0ZLcXqF9sg7aAf8NsE3rsV2O1+e7neGao0WrpTSda1P44eh4JvKdq4c+sqZh+XSe
HVQRIAO3xWAIGbdBRyhhIPut6XNIHmQHGbEIfzNMzSoHpw0fbuWfmAA/OTQpraVL
yL693056W+lZJWzHpmlCIj3m1pvaQVqK9k/EY/d8fyQXCGYjqo8luOOV0FssQmLt
MrD+bZD7P4Uni8PlVhkRBnlH//3uw8MnjISvyz1O2XS8I2WT25rW20X+L8cwEv07
PGGhfLnpzw0QPJ8UY8NWAFPJLn5y6qhqigpTCEYdy/VMsQVrZ1nYJVGhWs7j7poC
WqQZl4wQxvd2knEpf/dSMIwfmpuisfkaOXywP2JSQp3lT24ELoysuozqEo8fgLsy
hg743GsW3qq46Ajc4WYatA==
`protect END_PROTECTED
