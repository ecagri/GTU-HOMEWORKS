`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EDdWyD3gb7YIM6XXNVVc1A9wYWklxsCHHn2F6uMzBFINiO1yk46lwpJzCRGyth7H
UaDre6dQJDPgvgEdns+rjwIk3RHkiTuiZj2mcLIo/9MSs3ZAGcDaIMaPjjSNOcUp
jrojcJYhqqhivxbRvEIYG9maVZdx1TcluWQD2xmvWdcKVgMO59SWOzG46Zh0Zbfu
/nMZle4iRyXOTRbL2zQ24Tn0/ibRUy/woR9GxdHpN0BpO1WAtpt7WXs+FnEPsNoN
2fL7BUb/mh723wCfI3GOw98SvyBeDeSqFFTEDy23mHib1zRhYB0lzLkbw1i1DVdr
j3Tu8tS2OixcjyED0m05qEABSh8fEA57hfhMX2YQfM/crEXWIUKUf0eG7jxkg/Tg
2+bdp//isXdRji5fRx2WkqSIK3X+QB3xEh/Pk6KgQH/0VIMGcYBxtlwOyxKUdgaL
hetSbh7FXs/D0Dkks2W5TkKTnw+8TAZQeBdga5MTtP+tdh4//XueCjs0g2tKTgBY
OsEsmLUQxCG7Rzp/0ASB/7+3cw+30LSjVAlyM5+ZIh0WbLabTgOKY2trnH8f2Hod
qu1cerOl4qzOgkFvZ9haGyRjZsp5SayhQTpFjrPFnqsuSkNnKP5TehKOIiDbZc3n
0NbVECRl+s/6D/ATkkToK++ny2WOsA5UB/djTG8ypVSXPMFupw6fQfi/yawfPEbZ
wiHEqyIWX6BQ95Zwp1e3hCsUK0CppbXf9W9PoSVu7bhmuTF35ng9umdbcX7t0W3f
Ea+9u/oLntiaJ0NYqXKrJkxxy86qnCg9rhvlploHpYlKxReDoUBGeRYTCArBTBn6
wvKxhKC50DkS0zVCJlkEiYQsO1q1ko5a3Yv4iTAvi4Mj5tgYlVt4o050Glbx/YFI
GlcUL9pHkIudI5SxGb4M++fp2drlVPhsy2l0M3wImxhBX6BfqoEc0127cvUgvvC0
YLRYksPznbrscmSlcyz14Q0I2YWyBm+zLU53/mXCfkFJVvO0wMaCOQghhnSuobYF
KThlD4Nt6lrkcvV2lIQmzcZMy+on7tG1shO3Qal1/Azgvml570nw7tKw4tBmVSAH
8d0A3EpgmKfWe2n4vz2PDnr+Q9ZEdA4AJgPvruDmzeJwPRRcpaAiG+eDGxKp0OxQ
6eR5X3r4FmoHfuZNKUK2bVIr74Tkipv6rX9OqZzWvAIMTpsOn+qjr1OU/RkY/boN
28WQGsl5QpafQH6pxkdIaILfTB001pmVAPCvkFL+iE4i/rOx9pfpZ8AHQzVbmJmZ
uFn0Hf2+WnAlK6GEEQMLTnZGinqAsn6+ZzVlEjcHYeEGskKUX4lTGSy8FX8lz4Hw
cZGqBMBIxHxWl2OEpE6llA==
`protect END_PROTECTED
