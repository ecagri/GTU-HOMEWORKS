`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l70ec9mTf8TwJTRQCEAchKKcFdKJ2U/mk60GJ5fIR0zN9btQ3uhaJ1NpjkW+euC4
9mz0KEPFemdFLPzkZuHH05GJJ7NnLqPwOYjQ/F0nyh/mopnMoxXr/vv91/bXBRco
OGn2zeHxTP9YW0hxZ46S1px10SHCqCDQAYD3cpjS5IAA/3JQLlyceOuuo2bnl1Ql
K+9WnhthfQkW6Mic0QCGYM8ntrxQcvilaPnLNndNr2BYb4wMHJEDpwGYsouH2RWH
jjctLXi9Y4nW522goVXahh4m75v/3q2lJ0rKO5ngf/pj1ndUu9ElQMT6iLq06/Rj
+Bpir35IyyUwnyFQYLIfaH/bYflll2r4t2ziQXU6j5jybPBDbUGXcRZ58DSzbgZX
68+bC0YZQ0vR9Cjyo4u9KAu1sJ3oDSiB1jDAIkZXrwUDXaZqwF89dofKaETRGsSA
4JdZpdwateUWk5XoYjLPRu27dHergwmQzZDG1qbEEN1dHu8XqgAtyfXZYpG0FsFA
DmtY7ntwkfTci1XSvMbEACV0hWTlue4bw0sVwaB+YiBgfgNjR56td7UFTwWMuKA4
3PTBCnvqm3LQlvUj6Ev7Cmq/u3FOPAZBRlAv1uXEiEbWX1CYlHGY51JxHBoMDhIB
XogkjHQE5ssjiX6vmzD4jSHPiMYe0D/PlOuBYJmMyYQZmq7tmofyjllPxC2Jw4+Q
+IB4ZPbkVa0SLKcGel08sVywaxkSja4nVGNS9Dup7fSzMAycGz3hXdLFBtXWUkLe
gWtGY2WS3Ko4NNLkRekJ71Rh96uWaEkDr8p+0FHvLz0=
`protect END_PROTECTED
