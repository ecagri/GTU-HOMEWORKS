`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vv9ZZyK+S+SpYPOY2NK36eeeo+A4+ZOrOF2KWQIFHvV5WeaSndRiX1dnlxXnQxTH
N4LYq/NLk1sPDrGN8q1rc7kXFTZVt0FyPgNe0veHNl+yYZeB85ahPU3z+u8GDrOO
xZqvAuZtz2i1wyh77NFuRmIVcyGYOmGTfljwBFea+6FZGMnb6SQ+fD/P9Jz+8Mzv
3DPiu3YnNaWFDSFFdx4H3onCYY1h+vEXemXNcEP7QCw8UWOlOqCXVqNBBfXYihFG
RLkZ1ZA2qyhDT6queW8mMiUkeWV4ua9QPOIzG7YBLCHWSBLOGzF0GxyZxb37rSpj
XI2IFxqp/EKwetfsaE4NBJA1gYJyXvDeCUHDuZS9U3WZdaF5XS3G+xpJRmIwk6tM
`protect END_PROTECTED
