`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qKAQzYTBUPiXSAgmS+VT9hpaU+cVpMgjJCaDonswKVKpEc4Lrt8f1zJmcwW5gMfq
zhg3iFGgd4n4NCW1x8n8J8048kslstM3wN7QcWAOSR4/EHd9zF6ufGjy327WcCuN
3gYHuoCJdW8SMzIVIoSQUsJVDe68pugLhy6rxOB9vUai4ajHoAUvBxCMfZbmiRPy
nSMh6airVtiXxNI96ED7MohWMC+sWf8h7qvmG06bbUbhD+vqhGC5Y7raYM8LiD2V
e9E9zk6o9T2EJmEP7cFxtCFPWxZidnnVHGT+f53qHDBJxYi4sxw14VeAhxKdLKd0
7BibwQHxwDrmthAlDzZc53+UA2bDtjMz5OxOLGd7RUFWEq6A9b3f7crsVrGOvGTV
oEdvhA75m05TXo8tS8Tm4LE/tjn2VBPywd4Oyz1D2QsWAYXjpdfMc3U999NgtaVi
ND5gGXtO7AahoSxKbn1V3DnB6zXKufthEtk7TXqBzaIPHI4Tf4w6JNkqsMhVClaJ
m/TCYljF49I2wMmLOTxpesBRF2oaeSO7Maz3IhKQEfpT3Ph75GvYnY18ki+vDx16
n8GyU3XxpVCo4El4gRgbZAu7apv0V7cGDjQ5N9C6Sa5wA5+vV/Ob+bjZUdK5xGjF
MV5R3tYSvjSA6hPYuJ0FZoTk1YMNpnJFCdBgo29AKOZnMQduTjpXPQccQ8VGENtq
zro85ogaPq3IIqAMMhTEz25VcmFxZ66NKWGNW5+ouOyJ76+fXuVcMVjXLuxBA2WO
aJdszfkVagprDzNpkh6zowo0kPR7htljbGPjTqiff6jTZxPjyRkb9lG7m2qWvplr
8IwLJwxOKRPN+W8u1OJyNyb/xK3rXnwoYhcFRgDnDqzyf+tHQGl4xsuEHNkNcVLa
I809RaCP1BKWtl6W6pqMDo8jgsyjqu4PDPQJT0p7DfhXEiCT2eineqM47jcGTzc/
+z7aV9yYxymbgjrTNTbtClzs/ngeiiwFwZx6xcPi7gEN+Ad9wHLtSAMA1TNBB7Hl
Alzm6mUFIyfrfz+zoA+SvOMJRf4ehNVM5yX69DgwOtLQEFQ3bDYNxoSM7LNy2XRE
gpIqvlRn4eNQzKzFJnusgSjF1VCEaOwmDs28F2z7zD0h81VZDrx2qsqwCxVs9yuK
TU9cqxtgdcKyatemRBRkznlz2vwo5BAXy4VCAd6dul2VwArFWLfQE34DHrAv/E9h
Ttd+DTSzVwcE6m0i95jSMTgfkutCTnhJkrzkk98/pQixSiVPA66YbSTUX79+KM60
dQJMNKVHX8ge0FrKC1pAt0xcuL1XotgdJOA3GLnYkH9Typ1/HjiKra3Ikcvv4PWv
AzkgLegACi/wkQeA1L+h79+dFUcf8EvjXrWaNHs3QO0rLpXBZifXFUPOrkGGojpF
3YcGtKgkzso87WbSOWHextxLzIqBCHIHS3YXHoY2hpQP0XRNk4yNvsiH00V2O+JO
w1DHfOsHitCELWPhowOgaNXMxtujkom3XZKC6N2ytjI/grisqfB50AMja5DeDWxT
/W/W/QlUwhaGqumspUvR/6NA4gzcEk74WOSUEbTgvGw+t8utdR9NrQdTEfZDS5AN
d7AG4rm5ObxtaUQVEhhCFUerr2f6gJkuTlmnCFZQ/W6x5nwc7icRCg0VcxH81AMX
mIZW14uj35qErrihrz1bjp3ssB19WR6J6Ogz3zS6vxpJcDYSMNuBlvkK3TtrwiT8
9zjs2otbwOeRNgX9OtGrkacLUogNWPGMqTcx5NhrJu+/tbUzKLCzKxMFI49O5W+x
taYqNtXQPQ7K5A9DNQJ8WM1cwqaJ/uDdS7qNFTW9JUF/KCCpEfdQmQ660xhEVN6q
5FyWeReO5yhzkVFcMG5RAp09u3Y3tQjRhCoxGNLDC+qtWa3nJdsRVKh0qcrOYiol
6XdZBwZFmkruagE0HCCRUwWFtgSvoS9FtXVwArlt2uOmXTeHjiXIpbPBk06+rD1M
SsIsaWvHpriwDvNXMZNrxHaHfKEmQFIksX2Bs1vQgMNhyP0i+Qwbwdg8nNKaI9la
116xGr4e8csR0Zudlv509b/K57NR4u23B22QEsChT7KLlYAfYh0LfAZJNnBExi9i
XhZYx9ExTD84gec15gB37RRITozC897dZUggpJ71wOcQzywJDnZ134scL3FeRrHW
y3knzTAE1skflsM8rx1wNrwqmsytnZuKfO1iJzTSbStTTShOl21Re7eAC1oIs7Wv
2fR9viu2++SvMY9zvLfCmvEXpJsxnLu/lkkTpepQBeb9v6obLK6e5dcOKofI3QeA
g41kcT0Wm98wy1d/usT0nFSPqLaSPFk5NbHzMlZWubVQp3u5tNb/ffb6rAX8tEsR
DjEQ//1fY3AcwDgbQdwVsRgDQaOCZqw+BoXwkZu+CZjNuqIsSH4039dEoVV7xL6u
WwTdgaIo80Ac24Ro++Kx0X0u2FkFo94IevpJoVW8AS6SCv6hnYs45rcaqkJmiC9h
SsAE30D75k7NZVlxhMhWYAgKevUcAoh3iH/s5F8VcFkO2xiaRVqPCTkLyagxcbwU
9RplByrfXFF8zXWkBbz5huBOo+1SvFehlLib+bvU6xAZpJIhBNFWgCTMsCUlTtRt
Cb+QNT0PkbhikCyAjbK5QI8o6f6JTUkv2JVzM6bzLS8lm7UNWSNkt7E6pw4b5OOl
QSxUyW5WhW3Tv7bQin1dUQetGbjKW3R3odmND5sBpyM/u+ViOYhLg2OXbW6M8me0
vxbwlMnYMEFqmaoXx5G8y1lol6HhOz9QBVs9eiF+YKfp60Tb9mV8j1M0B5j8tTy3
KCRgM53DCYX9OnXYU+1CujCOTDcDCELB0kuFOXmCQ3zmqJsW9u1YWOJ17jccOHCH
kBa+E5gTVTIszoWNPTynKtlj81/yXpqyKw7lkhO5pJC7fFuGmog08nMO1tgbu33K
bTMTi1N/DlhtS1r1ATya7ZGWjYAASxmmr1qpArvYYVaEuDpq5tLuZw8JztbvNGgQ
7TMqU9x3XnIPB1t/ZCBKY7ObKJJCcvC0wWY7TjwWvIXSeDLBuajpivhK1wFTM7Cz
28S3hQ8jYRNdw9R6nr4C7JYDvdO5JuwAGv4T0TpGuunAAmVLPj4Qb0TBxWfzmr+L
foaTReL/vKsXOvtbs8q2C5SxK+daaxQx+Exr2GKKVTQguQTAsS0C+eX9BS9p21DW
MJc4y2o65Q8Dd8u4oT8iL9peabBAu6KJZnP/fjZ6FDEMzf9hcwecPYXr4QXoDEtN
nnQ3LN20ZHXyUiAraEHCWn+8dga1mb2MYMshckM7mddKw5F26G/X8dIDL3O00Jjt
ox7nLKO/m/ImEtsLwEkRqn+cZGYvaeab66WICbFrJrapvW1jhzHvAVSZKMDKdSeF
iLH8Vdgsk4tkXDWtWh9Gomb3G0R8504p9kp+3h/R5nJAgoxBofz66hGLPze2KL1H
7rTWc5E0BfWj0C5BJh9qQlE4wPWUFTK6aHHtFTE5X/N8bGMWr+7Um/zV+LuXPmSz
EzQQEeSGlIVYO6VXsCFvO5EWvcVZTRAgURSfUXShmZm8fRG7igiCne09mYySMkdO
15fjYJhBcp0suTlOCGQxMtHLA/3UvjpG3qSxMd+Vsi9IOSsaQ9yDLmriWBGvOdVc
zdqWYvCyUUNWbX0aOybnsW6czYhKDGbEElSUH1teTgSn1rI2zTbZ4RCSRmBfAd1H
4wTSYpZtMDOF1xLo0nB2QsHPAPWtXcu+cgkuzFmUa2SGSYuqSI8SQt/lpnH7kwET
fw/lNxu6gjOfsp9hU3olUc6vx81rLugUHVzUwPuUz0bdD2jzbmAFNzLanNxfp9Un
+y25TVakJLbPrJ+LxoIFJAWOT5W+6U03GLuXI9P7WcY9JP6AM6w6RbCeoKUc9olQ
5BrGAD2LJnW1gFNO6W2FPhTAEifGZAxEJ+hPPA3RwAQryywgJFsBOwy1Cf8sEEHL
KUea2d3pL/Z5qV+aEtUVTn32iVvdth74N1aziuqsOhGbrMWLJ3/4Ahy41QjTlMF4
My5YR1K9ujHcEh+PhsYwQ8AF7jsLmy5QfDsGIRRb7AaamrQsgOq3XbYBBhSXkDMO
d1SEX2HFdM6DuE1SuolhMvdSCehxAV3koMnbAO+GSbJptLbOg3XZAdNLHbS8VA86
eFL9kAQZPVsIt8sCH6L0bvoAmbFPO+jSZbeHUXF0XUBhlG8wQRxfo652KiTezw21
bUIk/QIsptiV/1nDq6ZN/gYJEDxhQocHyUn9fonAEgiNO21dQUrbx1PWEyljaodK
WAUP9H8zbC2SWxWuc/2SPIyhKCrP8VR4fahH7bIAQ9GkuuQuvuNnEZtmTs9vuFhl
LubjgMjlxgKl07xR8/VozD4zdV2RhvZHnxnlnaCaRPrGQyIQjP1wppDrO1tsXyKG
jWlvH63m1U1olyaXFyqDeYcE97ITfsFyUvKSrfpNMnlyORgobFyQNPU22vqluk/N
9kl3po7mwwA9zs0V4qiWCJ+YLJry84X4+uO1cB0oDLeW1SiZfy/CxsIUYXDiPYED
yOyptqkvJgd/SZTskLqZNKXdJuBzonPbn1D6x6wULDn/SISR4esufP8ITK9Mjmkr
5sPR30ZNbQt4Ylf7wifAYZJDd7Kbs8+mp/0HN14hGPXCy9qDoXqNIOH4xTz8Tasd
QYcIMGqKqv4Uwe8FyPE9Zhd2h5cnlpPDHMTQXzyktkBd2mGN3ex+GgnRtODLKbg4
aotjEQ18xGQKTBponJXf4dNGt3UVyRKfILYXd43VPWhumBNedLV9JhaMaovwjVHY
B7TEg9q4YB/9pgj2MfGev1AtWLH9ok/vCnQGrqwhYAjFTOB6qGGE18TuFXmd/4G+
rFAbM5YiAfWHnon9BRqosZVQ3Rgpq+foOllAx1Ls/L/XjiWCzZt3hUFGhNuhJIHB
5Ih96DVM34kimXm+CRg5gXnvpiQ6Z3f5f6OrFH0T+VBUPsssZP5QQHiiT+SXBfGe
OlAbfmiGFPt5YtOZz0M/T3TahFOwqs8gb+PS3J+XXvCDp51kW5dkTwR55ssltD+f
71Bye0Rf5TaQeO8NGeesHmK/uzmXECxcH+rC1aNMOOoheHlgMmji1MtgtkavZvV7
MPozdlqpC4Zv+/kKIhmEypL5ujSrPLcXTMCrS0FWenot3SETnyvaRovYbttOJ/qE
ozXnpqUWlhzYSLdKDhb2DaRaXWTb122wcsHHncPTmuDAbiJWXkqRK83/qhpa497n
wLNAWirQU/KoaS7EOS/qxniQY1V4vgut0CCMdbcvFrHSwVeoKhBtD4ngKw89/a3z
EncppsvTcn+V3ZiN6f7Y/fNcE5mTT1iyKpV2Ll/s2XhycN+thVD7LPbGYP7TCvzy
K2oxMxfPTVIo92a33PWGLaihKdFA7eeD0cSpqB7X/8heyI0PQ5D2GBwD5Jn10DTl
MMeROCibxZz7q2z/GAKEfZhf6DBMiCi/6D8XvctDPfqPnzry796vyNZm4Lt71b12
Gksd60YKcEkLdZapw/I/mu7jNAHPdAFeHyT9KaSFTnKCW53UzaB7a5BM3kxo903S
ZV+qZCMgmQ7Z0jmjltjx1nJPG4eiwHI4A9TQdwS8inoFPC9brGMqmeHKdmp4N7X/
E867qS9jTbZWIqtQBi0DsH10C7vUZ9iRv0f67Np/iSsSBBcwFd7Y1MViqQSZUNon
qhFXYm+z1XPtldmPTbSlVAqcwtaxe7HW1lS3GYDLDGt+AQRDyDoNDzacXu2EpRSx
XrurfBwIk31cKYMnOLp40GQ5mZAtuzhc6kucViASMc6k5ofvHPxEG780Dd7wi6yk
ONyUCIpwwjz1/6/0Z/RL9s2R54Wn7W2ZD4+0dlGnlwcDP0It6Nw/govsmnnCdic8
zBseEXm+UvhmQaJmjiPINJaUTX5JLpBNoQzXE6CHfJ0bCz/hLRoD73ngGg6jhxHw
skxqKOXMZubAbSVyE0LK1w7KRnoC3lw5iPgm0BCdbrC0Pymc908v9jMgmhyjyu63
EnGkO/Wj4GwqerOfv0TsYciSMqmNkeSdNSo/464qeIroy+GsTc5NS2kxXcII1GDG
vZ6d9dDhcAUAxBbIAMpWFa6zG3BnGeyUhdTyhjsBMEEIqd3ouFHBtbJD9p2nQZZ6
lza05h4fbtkOOj78g9LmJeHmWVFBJwanF7+ThFi2rxRMHGRtui9F16ps+Tz8wjXU
+xBxSdf7L/TMEipbFiiRFKg7qFIhVoB8XwlA6/7PVj6Obo9IGRwiz59WsgXwHLeW
gVUhS50aSGKWgfn83vb4toWfp5Q7Bj9l41pxL5lHrCVYNIqu5YQGNxUc97MSL+b3
pB/6b2J6RQ0GQAWn1ysx5RBJSqeWjEcNrgq9/Pj6qtrl3GE1Oxv0CbAwF3p++N2g
F9in4Sp+92XiF+MPAghhV0Imaib+aoN7RRGZ2s4NwMtSri5AZaXOI/7zf1GKPl9O
XrgIeiDsf0s5j4Px/+p8og==
`protect END_PROTECTED
