`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
veipZ015ZTa53yj09ORYFLNROvSiDF6kVMeEnq6DDQqvpURWNgu840BTFyIufE/e
GlYhDWa1vgfbgfpgA7wSYOGdjxb8HtMZ7bh5Q+RvVQV2XcQduLjSUq6KHcQPASi6
TziwKgJI2OTS/f0gWaLXXP+WJu4iBbJ85yt6n194a7RvIChIM8TbLTzYEx1yUMLp
L/g+3cCp7u3qvN00zXdPU1BruDVvDvYbEjNIK1IG7fR092IdWD2LTdXq4QVDrFnO
di8hFurhnsAhbDe+YlLJNqf/Y5LzNjtrhu0oGSqX/HNZi//76cyC50QkQ/9enTgu
2uqOY+g67FuFveEiPcqysNJYXZlJaXsQJJ8hKffJ/IWf+JrbK2d4VoMmCgbwC9m9
2qPw+HhorisJF7ED8U5wsOFzbErhnGwovim/M5ThJwOoKnjlvpCTrrkJQX1Jx99D
fiZHFSK03Z1J3Ak3hK8ruV7euui1V62rY1vr9Jmvq+3IAcCJVPiVM9Bg46xjLsEU
c8i41R0JnSOH5ccgs9mjYv22G0fs3gqHgZdC8W4V4Crllk+fRpCabof9xx4q2kVu
bHUJW8xHUn0CrKdp+pt6OWPTCMY2ggy0FePZ9i8JkZJXAHCN1nhAzfrzD7XCOy+S
MZTkHdfsjBob9QlTo5ZNiCBqakF3ZyPrNtjkarhckKQKUcGEZtpUhbL8BXEXBdNZ
wnBBGBdNqspMgEY0ThubTvbnr2aG45yJemGgti0RLwFlyoBZ1IZriqTqOnXbB0+w
mlcpGnbTZ9FtXR1eHGdV6tSB3+asy4KpMipEziHS2GKVRrBn1G38MipOe9d3lnNX
CI5sI6E8PVZEMV/bAbyc4uhvvudGFDMgTTX+7fOI2XjKXMwHykCizW2aNqWb2mD5
jlEgSFMSNdmICxFtYRETN6tJ+89V/TeQMP9ezcC5M7Rg7XBZp3VXFdLxrAUALaQZ
z/bH7xf9s+RntP6gAFirQzlzklo9KTnY12zy7jzo8KmvkSnWdLdXUZXI0jfzN+xX
cs73d9AyZ3jRbmwhq04CXiVZdX4ovkWCB0KbTFNudK8ncHf2YtXVcpgiK3h0ExlA
vHwmljbke9MGrpn+SI+nliGd6PZeCzXiNZqi+2SPyQj5QxScdPeqblGsFkNWlaQh
IP3HnLNNXkOFrHEhLkXX/VsejwkQzxf2H496Y7lIO713HR182jfD1VhAcAOTQhhP
DOZqQvlQLu/LCiyCc0BhxZatrno3Y98qmf521eXZ6hjsB127YbodGpa1ZNoRJvpj
oLYqwX6hC9JKryfBhSRi3boa9r1jnYX5sd+WjAKVxaUXMRLyS30Myo1fGbIwi3ht
wd7ZkA8BtfTsdGwARiWh/IwAZa4vhvzu/JUeBCsExDPzO48P/b3pq8OENI58n+mY
4eT5iTu2/1f5q5+QtTgSmPIhPGVPkLgOiBnQAiv5yztVJqwSjPmpa+Dx1dLIqFWx
EN6HvGp2iJb7xIgeuqkB1oP8SF4PzG5Cz7qsc48ECYRQP5gbwjNda6pHOzhRE0Fe
g3bS2elxWtGpRFDWfKDLNtdIB5nilqEfYh4N/EXaVf1RgZHALDT4fQsKJrczffCV
srZnrxZQOutvehnddRUulr4yTdR455nwWEinZem7fhjbh6aHx8HZ5hsd5uk+Gl0S
ohpuUFKxLPqsUh/jo8V+IU81Q1ufniOgUe3AHU5u+5v2ioyZHHLCe/mvL4D1023n
Cbp5JhTmk7mCYLE8a0gWwI6kb3Hk4MnLXm1+Dnc8oGCQAYUxPtQJA24KBQECcadv
XnSlvpPBc5tZLPPAHsFeTJ3uA4widZzryUev1wPWuTtOy4OSg9DTpX3P2v7h6mVV
LuPe25zfAQ7UtOeqLl68t5aklLqOLDnmGSPSFUViVWY=
`protect END_PROTECTED
