`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RYTlgQhmcRoWYMM2XHDsMmj3KVWqlcP1SG9w6jeGcqeR6apBT+6Q16t3eoGbvLId
vBG+6jbw/Mat+UaJMBg8n7XeL3n9KjVgAcsgrPh98GD2hlFrSvyT6cK3fwalR3FE
mBeTOlDt5qrDJmhsnZZAKuNVk7fL2jJ95yHuX14BnA9tcP/oYaBEldJmyCDj7hFL
WFhvNTLCSTbIHNZRxr/x70eFo/ZgP9HCD1maTVNPW/NlUjtaE/QFjrXrJTyG7hwQ
KOu/VQ3wRHiCkxpuvdHwD7JmOtqHSr49NucIN4BteU0ZxXJvRZMbY/XLM6NYYBdr
TpDLBFDsjeswg5MxYcypLoFf7ei/n6Ty7xi7hKnthT0VPBfDNOG5Y4bDsgjlQQh6
JpH3xJMMAC6EVpf1KOX4+i+Zm1rRMSEV84io7u0GKSEHynBd/jvQxafaenLJyMCp
q7Z14bcqXzKNNaGcSTJflPRL24u23/+uq8m/QKomqxlTnvHdcUlO66Vj0HmVCMMt
SP9d4xtuse93MYa6MeBA5b8jPZSVDayLTsG98K3MpN+776jNruN558hSZxYPZft+
U+Uc3p3WLw4CbVuIwcTer9bLxR+dwzJvePTl9YMBptK3KWJZ0iYy13z79OMO2AY6
MIoD227f3vZnVxBuLIt2wn2qAjD4dgDhodgmkT01MQKkB0+O0st4ADq6ZZSqR6ay
B2aqy+08OoHzwQhfDQty+dxh4wq0TsSZsLEJ3nDLMFWUsBFkiDHOk9Yd6qaRXLoH
AKkWzJZiTGMaUnPddxQx7ZW6ppujghbNKrGlY2ZdIojfM5IaAybUFVvQoWvrEx/W
e51q0kAgl490O7voFBYWrSvz2gN449MCl12caqzpWtOjiZtO7hmeACek5S8Ur5wL
txkp2C44cfoUGQD+vHQUE//itPC+DOZMR2vNHUZbtIdCG6ajlurf+EhFcFn//iWh
bf10/wbk+Hsp0sufQ/wO+VRIeR+pXCiRZdqHziMlJEkVPdLvK0wOneZjjMrjgBea
sqO2y4VgMLsG7Gps4W/v3KiMGHuEbrjaKyq30QtJB7gYPDAI2glr5Lz2lAOEL7yh
dsK/tk8DRQhBBj+TTe9VFKK0tIjI2MB9kE4ZFbSJamSSwBCPfD2z6QmeugubuSBU
abh8sq4j0x+V+BdhTsFpgM0SJAm/ArJet+++pw6exkjoTUC3g1KPrab7Dep2AvKf
PBX3QeJ5MdfKqJdnlj5Q1Jow+KMG5MJBEXVMwYHFUfixoydvqwxfPqihOMDwSYy4
NiAzeCbb3sRbT5OYjppjDN+mIQoS7Rl02E3RAxMrIC+DYKjJDnI5Tg1Mk0CmsXi/
DsBDbd7NXX5v+PRK6s8QvrwZrjTzSOdZAf/x73jHwKbOQCoriuJws0XAI2J6yyOY
suRlX/yUig2e2N2rAP2qzZyb6gozaSg+o69fdAl9Ha4=
`protect END_PROTECTED
