`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KgHsAbXgyC5w4iu+5j9XiVfb9cCxRe1DDfzjjjSgu+Lm5ct+/mQMk/rON/HiTytu
n8AUJ23MNIg3EOOBKL26TBUSvq1lIpEE+lL8bVRUnNiZaVtuMtICBCOc9t1XSbdc
1tH4SJWiv2BvIJBHh8p2IkgjOA6h23enmwuMmc1zO7I98OUgpw3ZMdJBXFaXOprm
4eCFl4sPr8EDQ4E64ucKiceNwr7LV0VaLj3bzZwQzoBW7qE/Y9VP5sYUO+XMImZm
nVbD/gF/Icuqy/V3FedRd7MMkaPMOfhMq297SXGl4wEaGqJ2vQtflIQD05Z6s2kc
ne+kX9uApZnfT+sgJ29Jih6nRO03LLkAa4k6Nn/TYOv2t8pElvKYsLUNv3bUCNRX
XPa4EzNR/53s8J8xPIaxCI38+XSNV3Ve0K9MsQpktaoH7wY6pm8iUXARV11zBx1s
tpCskcMc6JxiOrmhUbhHTwHvUm7TYNiFOvaEP+zL/OevatXg7f4xNqewAW5o9IqP
uUjrNc5nCFselcG9YH/7PG5WiO4yrdu8khgDefG5h37hQ9hceKV411AKG4rqj+cA
acyz1l1qtDPXrlFhL1fBDH6aPTJOxzeSk2Pb6JXgJx4VDnJN19wchsZPOWZ8Sud6
XNr0bZSZiASWIjGatE7OrMyybdAVnX+Gthhe2VdgdHXMoG6i2M2pprwmNlke6FKy
DA9zcZGManIO2Tua38WazBwvkfQgE4oeFWQxGT2o2qCda00wmlvwAtMYRFziuWb/
Sqgv/7RJU+HZgDwx11o7uz1DTEr2OcBE771Qb1zuVUn5mUKT/qY7sChP19KPqdu/
+fdC37ywRA0l8J6O6YiMMGzGgqYYq8GM2YgZ9mIOPtx3GMhwOX7tdGa1M7qx6OAC
1TIBURZlQk8apZE0wC2mV+/SM2BNFrjW+GQAjMr7aWOKdjfqE5mhxfm1bRwY4vHh
eMFgzbP61g2bH5q3mmn0SnfG/21L+wU/AGpD7f+AqMa4f0TviVvDLmlcG5P01z9v
M9xw9JUyAIvujtD1ReQqgLkVLMLoZZ9pA1MoMlT+HuT6bh4EmW0N1xBR7QKc8GTR
9Cnh6BdAt50eN5IAV2yVhkk0IvFlfCoKadQVX1HQYyXQXiZ+EGWN3YX+6kvrPMDK
oP7bFoBNt12+XcJx7jNufyJ7I9fyINNZWBpLwfGGxytX11PeI4xdOmX7quT8GEMJ
j87b/YI1duZ4ASIDYs0yIpovTKAnvadKPP1/Rsk/sqqfz37qh1zjYi07/1QLx5M6
IgkKoFtHfh9P56g6iGBdd0cDOaUvyy3zkTnWDLViaYUbG23kd/S4ghjbTbdYDxxI
qJZxkRDVbBTBfqKvQFYBvDGju+4KH2zk3d/Rj42ulm4gGSNXkHk169PeTN/nho3F
KlzNlkcxcRgNK4DKTlUxNJYxbAt8PsqM2mm+akDKnjD9jqa3J2aEcdk01BR55a2O
nRfLC5YETWhYXnKWhg/dqaWfobJQDbhn9vBfBy+jjxR537WDSBz9aWq3TJ6S7UJ+
UqSsJjqNS1lh5sV7cc0/d+13aTdb5JlJW3iDSIt1WH/Kg67x3wAZEcQtgEPUz/mv
sNcAJLc7TRjANPWE9wE5I5mhoGq6qhNMrVAylMrrrb40jDi+fYILYjTkkVTNx03W
9ErIKgMzbamyNOs+0LbHEtv7m0848P9iwAPVRralPJBrxTOyOJvIfrWXp2w/oclm
soQSFlWQbfA3T4BPPQNe3KW1VajlUK01QFXm9KSCIZLoMnVUwLFjBm2dJQJgpdRQ
4lFNS9zKj3wJDtNEUGSoP37oskAn3nMOjbDI3FcU5yn2AqVS+BZv8x/DQWr4FWiW
I2N4zubYbh+O8oBp6VXEp5L83xvJaQWvlD2UOK0gBbIM0SbRkdv7suHPNEYsNvbZ
`protect END_PROTECTED
