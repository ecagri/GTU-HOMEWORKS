`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GTgswjk5WndZUt8c80ID3M/zOmmWh35MzypTaPLijYdLJ4QMS+HEwcpYEREgtLQZ
yNVL9atsx4Yxvtik/o9Du5t1apUw1M/3MKqecCTId9RC+7bhVj0BHLMsXVk46lcO
VRdRprrbHNhhluwlnHl5ERXekVe9PLIuilh+5Am3ng906mFQVjjq9Ywoo8aVx1fh
BokfqC4nzVxiT1fzwx6G+nx2qo4iUUbgL8rugqKg+mP/yF5ezGhFLd5ecoP4Dxxg
Bd1p/9r3Ed+/2M2dh17d4zY6kHcergkQoa07zPsCn81Xa3/TxmG28NABORyaM7Nm
gJYalESbexbOgcrw+to74YOAZ+tnc0A2mSwpJI2RiwMynlsCcOeHgzbCkM/qM4ZS
c6P7ISL2+HbV9Cof/LCozsR7Vy49aWpJKJk9CNi3u5ooWd5mzFvmgapds6/SJaDc
wM2qE98xOWbUPNILBqVDGE3Qfu4VA4CaHYte4hnifR7mVVidkTKIKxzJL8getJI0
fmwRlOriACuZLzeO7nt7VjgF4mxR6+v4mrxb74ct/JkOhT/4EVq2tiAn1px1+vzR
pJtOzlFsGVIF0c6u5vWr11tgRnsAAtfK74a4mTKsiJeO+xC+YrdWRttPeDek15Fa
IZZ3Cn70sy53bTFwZ648b8a1mC3CIpH9tVAykp0R2FRetcdBh3UI9mdAJdN3wXn/
uLKDfqyKCWyrTnwG0tpdKOgIfY2q614ZsFLBp9Avv1VWflORkxY9GRZymUnYQQZH
8G0tQjh29BINynQ6jYVjrRCTR0fp2Q/BhQbGNs1qZNI8n3yS0Ih1ea3QZHVOiPXs
d+iwu468RN4OW1z1EV9H5JSJfvLchBWwGXrBCpfBJ08tDCUU27tLheh35wwCPXWG
uyiJD6vUDVIncCv10WO37XKD0WXAhJSdbJFwRELE5aGFhaDdZZhbLwSdex/wBPoU
OTSV9xFAx3J/6ya1Cxx6S7Szjnh42Hqqd01yYTNbqSQ2CyKutdWhW9Cu+yv9fmLG
mgeRl8OuXXYPSc8ADdA9JsH8+m90DFJSyT1G9/+BZ/SYMtFdVce0Q//a3OYO0H0o
AH3XaQQSM17FybW7MysrrEaX1uyD6E2+Hdf97anxtdHWeKdOcKjdg8sM4/pRQQV6
YTx0OSkx6MpPRybt/gcJrifX8v6TqOAlkaqI0wRL5q41RvBiPbkMuI8TkxaEhi9l
lVTCfiGrzAL/lcmPrL0/a2fCiB4S9NIUhauVRUwgMBK3keo12D2TOPbKMrH1vONH
Pz9NTJOP51alzc+cI8zP2wjXwubQZgnyoClaVLeK6WjVMuKpl7uLZX5kNcIKRQwG
rv1e3FHbxAXWbOfC+yVBcbVs2jepPJ6FLIfu7EIOSvXGDIuucppXCV4/P/HJkAGN
Q3Wm95wDlWe5+4rQbcnJAPGCt+m1RoX/T82NdAn5KH/d9p7NxMDvcMKXVckI8f80
It2R6hKB6gRVs37HUg5reRgJkavlkqaEwEKnKLdFENijQMmvQXR9DJI4TS4/XADi
zC2V0nnbgfTPr7BX3BBxl5An6IynnYU78N2muVKW4DFKAOyD8bTfPyjKsquJrQ3h
gS0Wha0JbNbOQ6+1pCqRItvcA5hytmwQU6AXrrhxYqLdnAhN1qmxt2q/rCQpiKA2
EhoqorbmDvHM3QkxWHGtLjvoNzmlDkDxhDIF9hHOqz2YWapFb6ZW+8CGWmMRn1rz
OjfF5f7XAv7bLS1U4LAFtRK2U21l6hD+g2mksW/Wvu0dKNKwE4w+Srhnn4n3oLEm
uP/BfCxtbhagd0LIVr4reSdn4tpzIEUoibmlTmLW7YCq4dRggRE5qWaEbdIWd7ux
OTfzYheKGBgenwEDmZGPkza4qTqo0yBtg0ArGLKBdV6tkEGZguPsmOtCP2E6fc/8
HfI2RffoKLqgVeHe/B++l8HMq6QA4XrhY3ppZ6QeB96r/ZPVQVL5irzTJ7F+6r+H
cRBfjbXy3TnigqmOtoZWYCwnj5qCX9h/Cq7bPL7U5hOre4QCjuKpJtgHM+mp7AKT
q1wmkhFRNkQlrJstH6lii32vgy3kVFElithJRRBrhV5MwxnRVN3TmjblhDg1diwg
iGrF9KF6KLeDCEgRssnDg6J1hASK7M8xoUQq61Vbn21lbeNQTdrf/OTyAIRyHSUI
bFLy4HL1k01+YDVf/ZHy0N86eWV4GXQMPuRHII3cebyhI/JbvmlHJGnoteU6+u0W
nlTDZcvELnSJrA64EOPh3bDLi9IeHhJU7GU06OBnvGYKkjlKivtj93OUkb5XFZ5b
XaoDyfa+3GT1EsdCzGRM9xAco9usw7hGGXc48KIe2m+nj4cp4UDdh5bAfUkJsRAj
7DbxdnA8fATLY4GLItgRCa9UkdokmzRU1LBHTe2/o0MtN9sSqnaN4ESa+zHa1eGN
wGccT/uAkFVKzWEZtHP7fa1mmqf50ZXRhFWyqSkYPgHF6svADMYWKl7OWVDNLC/j
IlyszUQUiFp/MK2HISRQRHMA/BYhqJdyJmqnh30tNhA=
`protect END_PROTECTED
