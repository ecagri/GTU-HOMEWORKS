`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cp1g43RfaVQjUW0SmfD4GGqfWVtkkYaihBZgo4dW601TtirhlmeoO5FgcBWOVFWy
H06hu8lfRte7/t+xu0pdR46rcRFiTjsZOY5N+2qcdx6AVy8tqH074uFLVdkyB+A/
J8k1auRhxm4tzSuvhoUM3gwHdoQernWJtOYcs/e2/sHp97lkzbGCwgZFdrVfZclj
jFOrehdabHe55LWAZX8jG9u1JKhOMm3rafySs6hX+aN49dNURGyILxlvqxGMdsfa
EKKwczLbhpJtSjVbi8VPo/JqFGjARgXz+7BsOMZCLgnBS79k2Bcf9B+oX5c1pml+
bUVgX44INQ2U1QY+h490wurkrUnJPJvtUCmwsrTmnYhGl5K/1VmWahmgqvypkEFR
3e7H6OjEZ7RlzYHfdPT773VoNYd48Jt7pORKhESYtJlP0gjSCRJMDwZQYmxz+a29
wlUXCSn9xhuKselcu0mqOoS/cfn/dSt0Ca9swSVt7j9/q8YlexfvW5ED9Y0xMAVL
ki/Ac2JN61YKgbDj6+/nUbtgHmbwLcBmeT3wtVt9PQqv5jIEoiGHYEluacLUd6ZZ
Ap3supgaJ2y6iEoA1XsB3mRMsLMPz810T+a7n/iIKgo7c1iiUeIFM6aV+OUM5AN5
PwjJTBAkuop1uSZGTNRUhlpP4zaT1TV7sFIP+JUvu0uXHrSC9EzymIutc+wIiXKe
XfsPg72LgexDbSmkq8i8bsJ1+LJXVvfSCOITlTjHat+s04+KTPPsK+nF06of/Lqf
s7VwUZJIJUagtbFKU24N3+KtLn6CrKV+zcWHLrlm0dC4Ml8Cx2+Uf2sU8SziEF2U
iN2lwQb/pKZpZt8aiIImxwCjNzd8mMO+tdhd7FYBpYayS3LhG+s+h0UGbVUv9Jtt
b+fpivcjLHVgHg1xKr+5jp1yJEmQCZ1buokMv3GvNcEJSHjgkN3230H3oZ+aNn47
h78cWc+aQUh7S5gtspWB1O77sfwAHtSKgZmsd7LDcpKOs2Ytu+uYSy8NrZxMCNSd
RKOHSeyxW5aAXlFDjM9qpSm7SFTdeoYywufpaRT1SORbYgYPCqyz3CKRkytjI/rc
FzAsXjLScbMX31yMFfn/hvNQzo2KWR1VTPDJW/3o0zhufE0pMIjMqaOlGCtKcjyf
Lx5JqmkCDO1IH1Gdw5Wp2XGrffjSNCrvvh1BNHsbPp86qOW4sETRFow6MKQjoFjw
eFD9cB70b0e1CLmtvlArq5OEJVHPNC/P+uvLTU0tXPnYjojJ7Ny3V7yMrIeTnR8D
Nc/EIjxLFQki4cs+eIpkxhVinAxKd25gmS5WYEjtTeVmb9g/icLSf1GQlyrfarQG
igt3AIsOMyFhapD1zR2Xh6lZoprrrx3dgc3M9yZbXZOJEoOL+a29AwIxEaXqaRwB
EB94m0eLyDXIHZu7xirdxvit/u9IsgW6vc667u7fg79Q3748epW7gf0HaGCDBk/2
IsUy6fJZuJWbXLsC32GhuPV1YPE/Gfg/SDv83wUulwy0ZIcFL+Q2wb+P8J1VQha0
/F2igZDewcHRSDMNAsvFmwvKc/IkrC4BFGHW//5FR3OQXHHU6ymdfts6rGp2UzBE
IB4WaEqMPOIVKonJrsg/g574WlrfPkeFgt+9PSLDULP/0BvcByUa/imd1SwQOdh/
TLHvgLsx8bk3IkveChD6SP+Zoey1zU4KrscZbjUQKRirSkYJC+K7HtsMRynlTcwu
xppmIsOAdR5T7xbk2E5JWISGN8JVJv0El6ahnKM5E30lsG/6NV34Krv1V2Buyzsb
SJdBeyfwKI5C9jnJpZKGWxOXYPAoUt6TgvPiaii+tipWRtc+bphW3gxHREeL1h/3
txkRZoDuf1QxOy8CFjIerMcukB/qGhNaDsNME0vi15bpjTolKJES0RsawCPbtiuh
JSVc3HMbsAznyfP0bBhN9hU6N5g9bdXT5OBxwAV6EOSpVFeBrU5Zt7wYhzE79xVK
0Qc5LbVOs1ZnqxDdweHmyCmZAfOuW3bh0RgDBG9WDYP4FQ1r8v+FaOYsL/YVNKhS
v929pu0gHUCXNjyGOgxbJUmxyoOr2Gv1rgJehuPBcLNpn82+ZBJjdiWHajWB7qPe
hvZuRqoKCG0VmVPZwvaX03V07w4N6zkBvZlNo7i/gYailp7zbNkYYZDkh0ZLM0Cp
7nKvUHDqbAjSJMAA1MRTjVuHbrR5BZsDLlj9J//3qdYZIVV+/zk7+6fvkJ3OUi9v
ZB7HnrrXnwG62Yg13yo15ABD7hMos/V2ig7DtpXC+BmA/jk2TfBacSodb+8T7o7o
oNXsuEYFykpAx71w+GCrFwI2AspV/HZiS0S/TOUFw2gPqJH5236uzRNC19mBEvzT
wsIJkkrpMoIYhelzIFwzsXt9hA5btg2vG1f9EhgyDvYiGug4iCZeA/0TZBT5dyA9
rkZ2518z3NpKzrGOCoJgqJ0x4ll3yRsHzVj1yWGQ6BZ3GVjSQXWviSzlg4HY5jXw
Gji68fSFqJw4h9QWiKuLxA==
`protect END_PROTECTED
