`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uGT+vWR617Ky0K5OBQpFc6sqWYbw/h+9MZef3Rxgqx9VWDmbhEn+HoEiGQ24K2Iq
dbESDQIIv0CA2Ez5UYxauvMrQaQuBlDY2LQ/19Gnwnj1x5DmdABiG0WdVw8xr+gM
0NU2uvIe2cx4ACTs7OpUmLM8hblrsmtZuXP+BEJ6qAAdwvRpzNfcYRbWDd/XwJIF
lqustHP0zKMju9LneqWxkmmllx074PeqAuGnVpcAdmYmdcv+ELsmzzF7k66uUCZm
lc2F430BhISLoBoNY2Ywsy66tIKkacjYKDa4XFJc9AGwqgnocdWzkkpvpdju/Cbj
kTaOSsG4UZ1JNQxFHSVuiMe16tiLIUVmEgKGikt321hSQoyM+nfyGERPGxMrPGOJ
xHU3d9MMn0ov1Kq4KCUwIBYhbcPLhsc0H16Kf/EqwHU35lmi6zk3eUj/buhnzbWK
GDysbVhbzYFp5fALRv+wIWIABlverzb/RkR0W+YSqjXshZQWHSir/o7qhvB061Pp
2WDMb8Z9ngNohKtZxN2xAvyaXc/B/+ZLvdjYNEwUouN4Vu55xc0iAqDLn41B+wO3
GAVh+vGwbVgAJrMONPzUX08KD8f1PpiLevIoMuy2SJZhhg+Ft6xkkvEHZTHRzHO3
mQeutG8Jqm2FLSvEs3nnsDpQ/RwbNK9KGpAbp+ptiTg6uqw2UpIJVY24uWHGD/8Y
SVRevOkYippguiiDMTq0LW9je2k7bEzQ0AcRZalXO9gBgYNABF+lzanvPl1FRIXE
aeKZ6/EUclgMRZt/RPe5T5b8xXRh+glAbysndjWuZ4MqEH/GdwPxNPRNf3JYbUK7
yZNrSv4RoZlpbgz0n9AxTzc0PNBWO00oBBRMpFWQ8F7XMoMpH5C0iJChPWcQrh+i
URdkaHIlw1BKm9vKJnAGC6oNGphdxiyfBjnpBuynSr0LARrmcuSlpeRNpgjssTQu
rxelvOX+VN9iSOYk8Q2VrRkiydXYEQPLq9leYI6IGQ1LB1SgMPyCCvWuAOCXjC42
r9S8ZxyKtiwn4rILMOPElqp2gpr2jxWjGQmhcaxYdawsiN3D9T6zoCQ38o+pGxd7
FPuncKGijqKi/nEFLXZxK8ebXmvD8y95B2wvhbypjkBEhsVN7EuneZZzEa6+A2iD
vCehLNU39QNdCwwyyf5aOibuzGivZosO40GgVgTigaCNunzE61VVa27kjyCxGB79
MSTXBBC5e6jnVjOE5p9aKA==
`protect END_PROTECTED
