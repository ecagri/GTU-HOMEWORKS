`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/UY1BEOWVz36g72a+o0rDCqwAyVifNIG1/Jw5164F1aK07pK5S0gNkr5K9wWd2ak
QPzdd/tMI7SAGkly6KtLg5Rw5kx2V2Zi0fkruGkU8BpnFj/9n/DVVkp7jbzHnB9j
znZGPGbuIjgj+vgw+exb8KQgqScwJJ6UaXxg4FaW0Y0+0gAYEmGf6c9BKLiuC2R9
gtMTUpdRpN4REUpwnMi7gtxOWpOIFYYPmYmFquaKjB77qFFS1g+edkLvY93mITGY
EUewek2N2eZOwkUvgpOSgbYR2pkZV01wscivVWbL4HDOUIJ/by9i9RU2qty1UGGs
EvHVU0qgCtsRn/VbV+iZj1AFmZfF1BMIZvXLQQ+eu2Tlz8/oo9DFHtkoQ2VnSaJy
JKwVo+vMvlkWKaplHNIlVzC9f6hbz45F6zqkP8WBMuYrAUXdO7HthVqm946x8E1v
vy145U4OpM75w47MNbooNN8BZWBgDDG5f/40ogtsOlVsFPRPa3tEm5P7iV5HpacS
wEqZ4Ov8jJoWghXFMD80QBccL81U29+MEUWyo8dlhb3yRnrFWh567cW6eXqvydsm
ms6YuEsVtXh8sFjnksXx4maEz13rSn3LBLNTc/yDa0uznl35NfGjuUzRpjwGC+yA
HeGkpimpjG0jEZTxAnTYDCghqukd2814KiOVQQujt2AW3PtT0x8R+c9OjyMDzRHS
3gZgMVbbEMQ+yxGN+fTshFF5EcGGH99Q7ODQmm5GJIBjMGpS5mdmdeKFrcjl2ZWH
Tkw7KMqueetf7DYlYlxDlrDFi/hD91BENIfHz/z2f7dSHCDkeYmk+wyphsnB1gqD
oAQK3KL6zwKLz/UZuTmjf3OVJla9Xal5IAT9NLuWY+l/psgJFnbcoPYYvRHVXG6A
6BotxEdFDGePSnJuGf/WdKQ87AbLkGBg17CuK3JEOS/9klVrlv9o4inzXv8crgFw
UsJkylSLnEwBpfOzquL9Lya/0MN3sJy19NEhhqpACFAvteugVGr84/BoXAt9lKTg
CwF7R8orDWpGrwPGmzIdNGUYxxJmNM53Dy15dsXF6PRDrAS0jyCCo9Bp24M2W8+2
6fGA9hxvG6XdAhdvF5+DHtA4suljG1PNHtB75mxixo5t4n/bJ6TvseMlQAabFutm
8+CDyjjepm6NRCn6WKQBV+c/o6hYXl74f9P8KKFl+ueNWCR5e+0VaFWon2FOlYUS
Wk19wh2dG2I4WuK4I4tWXe5q4TmgHB9COAq/MExQrkU1WUAajG05aGB5ohW/OEI+
EJrAeLMlHp/ao/8x0desaiYvxtzoHp1xwp9qumxLuNZJHpH26r+NYnLA/qxnIFoY
TTDTNt9nzlhPcafEfKwanOurUcPkAkV1Bqn0bKs7yLiAx8emtjnPGRyJw2Vbpa9E
ofY8NL1jDHKj/rfsx3ukAY0SmkNg3VBX5RJsL22JTSibRXM8tD6c3vtW3HGeFnvQ
evfKGAkU6yQJkPYhAMmFhw0t9P7+aTv7uVsxbk0iYLD9D84ME2sWhV2OPSTaGwF1
L8R3kaelyeO1EiHzrcl5rwIOmDPpdN3dg0SymrgYSV5DkmidiG6e912p2JZfFXOA
w3RmzvQi4VTjDuGzXHQuLy/Z6tqPEH0TkVBRsmWERWQnX1FiOchM1+YHY2zBKAGF
YCbQjeRbJqy07hMHJN/r7XDXTgz0nsBO9Mgt/1nJN4unTd26E9BtbnTQqEpJSAyZ
1izkBeFAmuQVJ2WF0XdC3rfado8OnLVxLdKVvRKwGgDM4rvyXosKVsVk9h2yCi+L
8bW8G1RcOagPUlEG4iQxi81d/kfseIER/DXnFvUfzxU7BQZry6Kmuprc4ossufRq
kljm9MAI1eChfW+rVPrWw114QiaK9bY/N/j4hau+R8CM1DsvK26eKjkcRnP65ATr
GMubsNAtYi7mScSKLix0VPcLoDP4vYF3OnteBAZ3UhZMG+YZWrnt1EVccshKQFKB
gh+/116pYkL+A+4+f9v/+4vm8DqoW9MG4+hJA/qqXM6lHAiBwANoZoi/4bW9bNiC
3ZWXOb2K9BNKeQjn+LfDMOOgNfHKhu17AB5AG9o+g5rCEZ++QAFVBDE7EWLD2rA3
TGOLtoYRVT7N2mWuN7ryfcUySpJHeeGn8BELaCgb42Ij5F/fIdbMocugEI4AKEdK
wsWc2B4MY6X9AqJeFpNv4s4p63vfSmRQDJI2JPdyLIWfctrxkh2FPr2AJ5AXPoZK
TGqpybDIrlPa2T9iXWs4S3KViVMg2FQE1JwaR3uz6pjOyrY29+6Q+lygheQn8P8E
OvIEdEFT+a5MO3NIky2/Fr+CNSyDtyTdtEOOSxPhjLZVApaySJIiyoVpewlKA+xl
V2c7GrcqpPCictsR6mYpfZ0QPX3elf/Kf6WPlnVehToqs99guy5gwgTSZB9yBDaK
3oiqYMu9AAUlhbRpFudBec/v1FCrcgC+t5f8tCjYrLeaGe1KhM5g47uSpWfQXVx7
RiSIUKblsFenl5lxzY/HBIjf59q8BzXH4gDCJQW31PVL7Im96JEzeWRAbi+hVmWF
hdv4Ie6uYpUD3A3cDW0QFmMbteavYM/iD/GyNo5T8b/2iTjj8RzhbcE2iSHbqa0P
aOlpUoq3ztdR2CS/7w7bNAX7aUhrzZQ/2UHomAdZq2V/mf9mOt2OO+JZ8QvLAg1S
/yJ5S8q+C1VQFkGqVmwl+xJHkBigj4eq/A6dlv6PUGnpSOY5dVegZ5Y8EIvCVJVA
c+1B0CQGFfl0ozs+7c8hwr/bcWbj96xhNhVq6ed1JoGrJOhKvnJiPDaEOi6vnOew
I6hthOly0sr5fRskKi3fiyXPLSgXXK/qvaUkCFSI8+xyv7S89LRfQt+yXSg+N+Pu
0o2Ofcst+EXLoEgX0R82GCKlRb1vS6hxtpJWKV8Ajn9hKxfyZJ1OEEtm5MNxVov1
g0F9Oi372l0wTNH2Wq1RwXFKee7R5cdEmhbchuCc50jx5hRFMMSiBMEzgUUlfpLJ
IuJc0ekf8lYyduU9mWDP9Ao5TEyjQV1hFPRz1vIEjTVdVQPKvL/Gec2FUqDpJCZH
zzj2+nW7A7MldaJHSqfeVl2s53jDsH7J39cy+aGBoryyTyYNtxtY+l+2gevifb//
NVPjLBK5csE+CHAhQ/dr6bNKnssdivzMuYZqgu9oeYKBR4Am/xOFQgViM0w3DLUd
a8mB3/A1IL+UvuqgIsgCkAAUHuDUv81lwo4uwMrwNpfVoBcszbNTj6m3eHlPcaDO
Ng5rJJxPhJmpFL9Ln4xCzQY22/L9v4PYGkoRZKV2TXs+dGPvq27yZ6bf8DzSWZtL
XeySMZMTrf1Ud0rDznl31m9XoMxTiD7ERuZLiYyfzmlrZCbHisx5ao9TrJey1j+8
TvHF5sXu8hg9VRGjS51RFvvs/zizvsYIjaAjrP8I+cgfklrFstq9lWmEHxmm/6v+
Yn8BTE1AdtVXuO8X3wfqH4osac+9vpc8+1AfxPw/jiB0aN0R/jTOrWoVKynPJ3NL
8Ig2cC8IprXC2eLTqEjOQaZm/YOAc8rN98JYaIZfAxM3Fst9xGOQMchuPKy72x8h
8akJGAO3MFzx+C56M2LBlBwkZxfyr70PZpBVk2K0v9jcXz/BfQFa2xiafqK6TNLc
0Zbf8QNSpIhlJMAH+ZepFD2ugjQeqaVsaS9z+CQH686LId72No77/jue0cQ/W7/j
35spP9HYfs4jLQ/Aaa+U5Qahe67hsszVoTPk94SojJ5VckKRtQRUAf9P+/zU463W
tPM0HA5kaIED48kEEp5X9A/4l8XrYiCc9aAYtIMOVC7AVZfRt4XuahOln7anRLGa
nrHJm/pSqlk2lCyeYmvA9Nbk3XjQLKCdEo6TgXLFUhP0bc/60YeH/UNfQNyLeovb
VP/vPCh2N23ZQ+tgFk+/QDY4fqx/XA7PAIrnBpkHdZhBksRYy9wreMNFIAAoTuWU
m/0l2fxqeyPRclRSXg3hbQ7ke+XL+Y/LYfT3hrM02nknLYWv17ohgbHPnQlMowNl
pXo+dPusoL0I5BftXA77gcicujOq3+VmKVwjjaZ5ti7yzN7gnrxKKlZhRrOloWnu
ZSBpdK+TCaq9GD94KiPAWy4L4kU4Ve+oO1aDx9MKl9Le2Zk/N92qRCbN7LnXx40Y
983KQ+6uIqHx9c60X5GHdOBeKw+kQzW9anBgw4JFK3ioYjIEtX2oPZ58Gq0+/xsJ
93DLprLh3TTnz3zCrPJ926o3JBezi3TzR1Y7rcMSk2iXDy8Zxx9+9lVx4PXHUEFK
0JjIRloJF+sX3sIBwjJieGIouW2MUYqvD+k/cWlsD7X6bcr8cM8pdHIPWKBzQLyG
1wDlXNlaMavLU9wgElAI5TMSfKd0YlhJhzOzgx3uzAuSPDA7wEbRwgL1yCYtW3nl
aVY7YHKSvKRHu0cMinVQ/YBfDrHeQQ0fpTJa/E4zzkNvihB9eOxhqHgsPxRlhb4/
SBjpmC4IcY9nOdlX8Flv41nNq/NgBHCgt2uayMQzDYcUgUKA2zFkpramnomcpOy8
bRCkXEk70XU+NexfvVNnAKgSAqlymRKY1FNgSElRNUUk9uSdi4lfywAKxvPvGNvv
SqSp1CKPRyDe2Y63zsLCnGs/kbDM0OqPllNJ9T0HJo8uYax4FE+EPyLta8zY6pgA
ab8X8me62IWhYcJ61nJhs3TNP5HjEJ35tpwfeOCVcFFvsvc2Fe3rJPboI3VibNZ/
pHzXHe2/SQ3Lz/rh2Wx6VihQAukemkp7/Arza8rDm2bmxUBqcJH6fPGZ/n7YUmZv
MiXqLVsY94i34IBUFuWfi66Gym/oztFHiIWT2qJo3atAgVTUK6Vsbzh+VRZYDX4O
Q3rRb5oOTW2zWZsJNylhSyzcMATyhAaGwCnOvTXI/ETWqyRBlXuTp+bEQETL6TcT
eV/leVfrJ78a5ll9OKNNL8iCJ1FHBVMLy6dbJJRO+6NmKZYQw58meX2sqUeCxr14
MSF54jJhRA2msOLL92FgAd9ngefxReC73ClhAaCQDuZoxdRMPUOe7eVMencMqVmu
DAyKmjjTyyu86c1QwSGpHrUTzxl0KPUlWS6ONU6v/ugmPw1a4uYu391LObs0iAWx
03gHv+u0LSbPXHW6ed5vcsxmah+GIkcwDjqKVqAgI6iCboF1Wh6HNczzxXY6YelP
QeqqHK6thleUZfOSNm/ylGcQbxkTJCgMPA6CyC0TPREFqjeWv6l5bqA0xcD7nnEI
+AT0gVGbJpWadJzSD0dSjkwNyxsTJMaGrc57xtszRrA8FbNa9Thx10PJQNd70bgs
YAHjxGD+xQMJ7QT6OelSjksVSwUMatcamDLZA4m4Lkxnysd9AIgVacp/i+HI0I+A
CRDuUwvKI1ndMrxZ14+PdmjXB5FZuzBkku5oqQ+y6hNyTpTxd5mX/7SF/kqaPWV5
SDZxopCQZIvLE/r6MsQllYX5GnzjDdhPvQ8XJKlgYoMszHixqcP9PnnMEZ/bQ81m
z5xis+idrWQuZ4k6E5X9VSRsrYVdvy0j0ySATT57OjUUKx0lsl75xLGg/56dVL69
m8jqDk4lFKGj1ao+eb3hkvX3AWhJdXi6I83VI1pK0zYSoffLLahhqPYIEVAMFTI5
zqfxNuOWFLTaYOrU9gUE3GBN2uMQCurW5w+XfMR8ExlcDJtoZPjFLEax1Mo602jJ
3HLTolVRHRT9/MFjg7EVcBC0wrB1gUy/on4DWLwhVyFamiijjIkvXlh/61SqsbaC
A31nrgKDJ01Hb8bEta2Nz21SRja4rloOMUX1IjihgyV6HPFTvjQDxvRyjiiWTd0P
BgAC1Occ6P5VK2E6+tzrwG1+Xz3kXHjKFyXsIHJ9e9eQSojH6BjGNeX7+7EFsUfb
VpgkzNJ+mwWQZ77I4DV1qjo4cTQcdvEdQnHj2BJKzE9NYM/W5mF+iwuVUUbmh/hf
IbkKRHziVeRtAohVimiODoM9aOuvif6TtVYYjp525u/5ShJjjjxi35USCfDaJ61h
ZljKD9+OBB7GeVyON2SC+ySei4uIolYXQxEAKCh9sbaRE01eTXZX5Ob9rRZfIiH7
iAkQODxu/zrLTCqrRElhQ2KFOh5m/XFjEV8MCoR9C42vIVCcB9/CJQnQ2DsYkB1Q
NC54OZcaSOnyxufstTGp+d7us3vipYbv4jRfuBUuy0RJCdktay8OGa3qZRoToqRp
tdwEZcWkiALWp30KOJI7w5HkQulIFoh6celFyvJrnTGgCOtGWrPN66he8SJ3Ijek
w++WkckXnazN+T8aSB2X7tiFH0FUyJou3xANc0OY7aDAewe+gAfYyX7VVhvE+a1T
okYIu/9VwjlLwdH24EesYwabPSAsFe5aHLD0GKedE7jGSHz8gL3gtQ4GbqiVfOSP
grjgDjCp3Xb/eBCMb9TOvWSQPN4+Ui3gErUoV+BRBwMlxVi0aSXRIL/YlDusttre
XDaqzy3KBTMgYfJgxEFoPP0V3kuX5b9IFNw6J4PGyycOeNiLIZaw24tIWxpQ26RN
+ioOtHDen5Wjx9uGe+IiSZM1GJrKmpPvhEZmY6f5v/G2KfEv4XS+V9PYFVO1d0dh
Ok7ErjTTvgatnBgtLNpkfP1AnwNwPt+pC4lsEFP+qh+yNwEasmDHpHh5cU1sgbD2
Rs58WOYD5WTOy1Yd1OMmn5D9GIkkJIngdqvuhzgIAOA7nTHl7Zh6JQKtEpjlGvqw
yoH7StaJb5ZedRCH97CnHiOT3KbuuUupSaiNl/NULkhVUNBWPX4H9+k7uCx+Jx+/
VXVFMgZA92ym+WxKUsDUOQp3QhvpBaOHXiQTz/qRlZTS+biiwGdhjh0hFNRB+2cV
IZulx/LFGQ74cNaYNfZvumtQADR/uz5Vll0xltY5ybJUiZ6KT1oUrclG3g2PHmpP
G1taix/dh6lDtOZA2ZY/iejGIe9mfqHtEvShb/PRs9nXECZ/ZnJ8pHWIG+RCzVMp
xPgG3jCIAZvRXytkpg2r+48b5m97q6aVHIzGqucQVDXxTscwJab6U9J4UrRrHuZ+
klMp5eBPInlfxCxJ3C6zL2bzauChOM1UAgYmNixXyS7FVdUWwMTxJYf25Bwn9x2m
W6KR/9NKtea0y6NyodTqRIJB8Nhz/cdQGeY0HfNixLCGnBuPM+NXmi4EiD166A5G
GJ+ocIysCtUaSJbqs3oZMAJ+jC9WbGLjxLXCLlkuF8x5jXnlRtW6ZVlsMtBMERbq
82IjMhLyS2OT0W20PamnUg3C7XowJWn9f4JrrKrF6jXEVz67ZferaMdpxHt7JAFc
Y3VQcxu9JLB4b6caUy9sL9Jf3u/gnFPOcYEmjoPQ38tzjf9Ux3m70GyV+n6a+Deo
drKnNEGAmRGt3ZuABkqIohnkU2b4Yl4W11llDq7oR7CRoESrTdCjfc27nk3E5oH7
ySzV3PhTDENub2zxLGrzFuUhZG+gqJGHmWlFUcMb/JRAJ2gXiffi4EyTtvbxlfDK
1SLbh/7tSKx00VAebU/C7Ogs3598u7s+J1R0O/boORFP2n1q/IMfKbVqe8XfbAIM
3rrBKO4SZKlp1fzYmY8A8d2PV+lhdp7GzRUm7ZIr3fK98p3/v4TUV5h2z/BJT3Gf
s26AhBJPnhkFgZOqJ1gqPN+hdXdo2Dd+WhhnHK5vNU+EyLrtIMz83S85ekCogqlH
yCD9I/73NpTm6SuAXReq1mHtPu2EH+gZRInAP8AS8X3Pg2jrGHHyqfwKwdul9FCq
1AKlA/A6CcgJg5yhZvEEg0myGOuJHOmXBBbPhBrFMpxhv136ldIX8rSrNyH3SzwX
KdB6YJY4y9yg7hx5ja/BhLH9nkTtoElR7aMKbPoIS28bJVgPUlj4ac5J89XyXyNq
eXyPlZTCCdnDcppJhjjz4E1f4eGPIOClUrkonX/SeD3CK1dZGOnppcYnlW8l503q
8gzKXn/hCkuFVBoT8WUU+sZy2ELgRoAcWD5FBL2CHRjwlf9jwGiA4QbUOpecZKli
fBVdjSWLhpVDt4HPxu9TMGDcLDljYhdORAZaL89/1VaAVD3Z9zdWAKodAEDIy23i
/niH/KoFlpigoFhU20PDAj8MSJLVA3gUCzozxBg5Ey0jUSLDnfVjSJETJ0c4v7U8
yuQ4mxxqZXpNtiN6k3uy+Mi6QF0HV5KleRTOxnRTMI45DifJ4M0NZ/yZF3wZHaOl
l7fvocjgXSOfZMMU9y22D2CeXNZRKKYf+BhXgCpYqw0JLq92skRnJvR2P0BhS4Ed
p7ENuK/mdZIMNl77/HquPA9AodbM4h0ILsoGVAX1qpMAp7WtoSuFu3RCW8guvYnV
DFdViEx9yj33D08QAzChD0Nv/4AiqKxFZxcASsVUhFVjLl7dNvAk8DTz94kp7FZp
WbdYKUMYE7mXoJ137cqhVIhb2GvlJ6rHFaohvdMKQAGGyAdlIAcGcjtCN8vttkG+
PuF/WL+p+uMlKhLo+Ms2h4fpSUfxB/Elbs7vxz21MmbiS/z1G5wTVLvZ7IHs6DsB
+t3B54h6sOmSVpB7wDnnmTpIx4mN2SkwNNOye4DVGoR4Uif9l1duRidnCcA2AbJl
gOq39mG7D5dkzKjpDaLVjxaQXltAldl6jBcTNhazmay62mTgYysSQoHMBywTmRWr
v2pDXffddQnKYR+9ulHI6eSRj4aZiGpe+WRLeirx05MyBKJ72sKwPpS//XTsKjHm
fe626ORX9exK8oVGAWJ9ItZUz8DUyvtGrkuSjDVgtpvABhzFs9CQltlVpTbfd94l
DZOPyjtmwotAu2A4wkBOy4lbSEMulzic0iHG18xGH4BrJsBqVr0Iwei555vjaewi
z/4OeBw7ux2E3WJ2E/dpuDpQhrf2ESKvjMv9yfm9MhAbJGkXNIVceWJzkc7Gslfo
yvm49qQEqduzEpp6WmHtOC2XTi+3kLZk8onsSBT5Ep/gck+QABY3BNz8K8ZsHCtM
sPJQQU6oQbMFDDV1UeTGcF57/Szi82um7rd4DIXBiDdy6WMD3UJivAh8HFlaLnBZ
rrsY+s/KwWZe0fTYpJCphCV+TcZkjmoZQ5aXjKMjcdBOkgVZV/ThPUpHHmhMDl8p
HPiqAaVtV2hS3eUSb45SmGwUPaC/RRVW4K9I+75tT7eWBFHfZTCGmIkC5tyql3Ul
N23Ic5Etj3qloLNZGsOJB4VdJ/iZXdNHwYrTfRdImIN//77ZP1DImA3VBYp2GmyE
I2NmykzrSVeK1OdZgN2+aqIqxq+/mXwAXSuAB6fbaxAUL6BTHmC41VbIsMB3EL0S
LWzXexBpJBpGKxp2Jt8CM0N5kXRHwhNW1tb0v/8deVwZCFrjN2aHJr3WmIkAicAN
quK+ZkxDtf6SC4sJOeQZOZM30xOdcd8W6zQEelOeMLoJ+cOREGQl2uMv2L8OOgt/
03eIEcgI2EYrPiTEmYD6eJfz5E3PDX3j94ZKHlkYzlAnfjG+V3hOraQJplV6yjJ4
MP7ux638Dcl4padI6NxCW6tuNryTIqsNf5zQ0ApRNnr15IozRkS0rcOPy4fj/Ytd
eUhkmVW7Bul19Y7QmajgILKrNvk2JYqQc41CByo1+VjTHEk91OMSBFeP4CTZt5/S
ocqX7ftkBhXsRjIkxmD7XaIPx86KLufEUb9AzXT6vz65ctgT0eBs1uzdRpmYF6pc
YKqePgjwTE711WSgKkV1C2aXAAj7K4ZCqtu0KkOJinMrEB7WHqvdsRcV7K5LkWGA
b+sabu27HMs7/jELKn2uJc1vmbLfeFH28LsaIULqtZiouLUfiRbpwABWHr/nrJq8
ZyCOq2Mr3GRTqXFoBUotTDgbx2lKSiplDeJQH3tnbOuG/rvGHqlJvEhMOWnAEdTb
Ax9F39D4pyby3V1z+xmzX1Y1NS7+KlwnR1dOongYS4fzgckPgqx7zRuVBuDDVc0B
ChwQs06LjVeFK38oRO4PHKxK3JeYTrHjU0xL1u+KDmWjOc78DRJoSfIRxMP2aw+F
2vfcHMHBfOqyzXwIwsX8U+OmtTklhJkxoQJDmpED0140Ive5KU0YyjqAS1/+nUYx
JWHBryaEK/r6MHQAWOVLy2FOGyT+pZnTKgkEaHSYUDFHnsE+FCASl1nfuqgJFoyk
/7eUdmySHWHL3lo/JeztUI6ULk3/YKMMDzP6wSK9sGA5vk8vlYtp3lUFfa1rmo+4
ap25ArVW5B9v3bB1nCcAK5gC9snb182FnScxAxGnSzi5hcr2WQ+V3UndIBhxExV4
NiEDhfNEKzUfO0dGQZEXObkqrabKssxW2OzQG0H1NGRr464omBbJGf5MDCwxjF1T
Dc2iZReYrHMlBoVFHtJ//PLxfGC1WEeG4WI5mC+V4Z1XtJ1VHvd3gt9Re1lzt/ng
leEt/USfbZR/eRLsyoNfDH1OsuPDg9nywTQUcYXMpDgv4MMFmLNwHdTbnV9uQp3R
7sgSsnpkTd+g15JZKVhA88GBbPA83RT54s+ZRRf9d063ExVEcbUKq0WcqrNWGfR2
VNjh/9/ue60Fhvouoe8kgJem7cPU8hUOFvDV+gZssNwy8gZ4j3RZ+gperGQsI3va
AuChjuQ0WzYTpQlnL7xP9VYrpwNzUl5C92lzKubCN6TsJxx2GwgPtagHrQbG+Gvf
6pe9JZeTQ2JJOqk1J9/i2C4B76Kuf3ll6/rcWpFJa4MHF2pbBCXEry3Y/GpThqIo
aTPC9ricJZuStHlziB1NQpWXBXFvmxWHbRNGy4EbMAi1vZ8FwGMCze1sGjtJlndk
14lreZlIe/ERv7kKr9irir4BqyNPzdIW5v765Yh38eOv2e7lcOsxlY1yzpPvNUXU
nQwxA5uw2ttULPixVvEeKVnmlHETYq0EB+kVQizm5PSaWyS3ncRnba/s03PQTMRD
2jpMYQQ67TC3ReaiOrAXMTQ1gJ0gXSEh/HUDaEi4nOL7EYYK+bCJdSdgFyxANHxW
epImS3xtyAUbciSQ5J5KzaYUZc9Qe7XuAvwE2b/DZqehU13yVA9cqusiXJCX3bzO
XGnaYd0c6/BziQS/xIx6yKO6l/H8eJvDSvWTiEqC334C7lodPLtWYOMmn6MqgJCT
Bkh+xlmenBn0UN/4020Y76yxrXpeG/H6oWnsKwvIPzeegxjNzB77PW/gzrh0GAB1
Ynog0ht/IVv1usVBYRLEpnWk4NvDoboj25QkHrPBHu1RpvEKTl5CZCftkmqBRSqt
rh07sDANSfYD23xw0Yvkg4l9Jaf6+mmrG9hQWMuWuxZg6bda/muOZTnbGuwf1h/p
Tj+6SWwyIBM3GhfJchFmq2u/4pB73MfB/jwThsjSHGZ7NZ6Sc/PAkjzl6DKtBOMC
m5+6DEWW8uv8696rP95d3KBw6TM4tb/4fM/6W5N1onM6oTaDNTVzWBjS9aQRrD31
YV5CjcbS3usZxcLUnYIHt4zT40c+62hTi7MoTm/qPiolLbQy11AF9Nw96M5IPvft
W+ZEPlH2Uw9Y6rc4prfeIzZzKkftk1DElMqgP279EVGo3nK4rOri7tOxsSIsa37q
DAg6z8UvgsXqabeCqUcF8D+1TFzMse133JO8Jtpeg7h8mokIokuqQAzWVAi5ab44
9nawjRqEfBbNQMPcbwgx3YBqAuPjycizmFwexS2vXGGdwoeHLvUhbKwUc1tps85Y
9wqicVA69SUp4xehKFS12eeWokPPzbKezlcyXZ9g9ZxY6O5g536GVTFHso+1gOBY
t/ysKND0lrA6guZPAt3mJvkrePDI7dDB6BkXdsMlMyzhMICBWuJOk61FbsDHnXju
B2TywTu+HuWFFuGRqdY+PUF7O0q1cvFzXefS5ThPEsXdDPtHF0sRmoVeP/Yev+Sc
6GEN+YJ4L5UrJqeTajAgjj9cyyhl5Bphm021s85wKiW54zMg8BuKWrSvjkfhdqF8
ydMBwGpuNyK1sIXsjQ7sC2mtJ0t24WCUibJUKz7vduA2w7YCz50rUYFkA67Inm5Y
hzUCsZY8VR7RTpAdJxgFFZVDuhXElEdIfNkslIL0u/4eHmSG/vZU0eBjevoy+Hva
yvVd279F+1wHuwbCWBHQtZwmcTaq4v9Zgd9wDXwYiYkBdLWi/Lyb4N5oC/yGQGNL
NwHsixLkM73xJ3JFnx5PVS5Q3SluZG8WcIYAEnLMrcnLrfno5e2k8iiMYIzcUCUB
KxGptTZgO7cCLzGQUKilUquJR6VY+MMihnb+k7jAidpX1EXyCOdWk/2mLRa6g4hB
eR90DCiRubxgqknnlkIxG5MbBkTRbkIUme5DfT7e9msVi5QvAsnH53XWbWAPIG15
1QvwUu+LUNaUohz7QoniQSXOpzWKyktI1uZvN+G35ibWlR74vXnqA+iHPjKzGcTb
bsHvF3gak+nr2lG65+/tSmxZgA5hMDb+uYt6ZqggCpCCvQFfXzGrlZR5K5p/XmAR
f2r4giWrShdAHoi/OC7JtddxYtXWJ//UI6xL8i+2OMGeJANIAtW3WHrSkeGrUNA3
0xKDc2OnqpExWPxqejZNMpcGL9sYQSjw1RaKpcmOBOTqsl5OubhH1JIWGO5Eatn+
JvfFNCKwKEo+z0ZHME8aAu2r+dquLakQ9v9tEbE6CGoGKzef/QpqPSE+wBw0/kbX
WHSW041Vo0mhjboeAhseUKX+p8QbbpN4/WVO0ardu0ZcN2e2PkGoZPHHUEEKpnVj
FU3s07RNQXZuwQZ8qC51czlFTAED+/Zn9XHu4e981J/uTuWiCJUJl8jzzATEHcCd
aukH4l8V6QLDazeufMAdAu1udd66y56tY7w++y654WeKltScBBB9OHzSLkCML7eO
9oq316hH/L7QUYySUxVM/zgXG2QSNZQHbDw6OyL7yPutegBNOr0BUdHmgFmqC/8y
KmAIn4c7qqV92aTKOOsbYCbBH7M6qMSkeknFFF9OuO9wrULJFFsrRb5kUxae6E7x
Xy0+kfKJwNzePhgVeIwTt4rGCT1ugKQy3GxG4yISqkWvOM6im1k6bWZVA2czqqin
mJOG78fnDA7ekK6Cu9RnLF1bcfw4utBusZ+Qz7cjr08oDaU0/ynUPLdaeuFYYpX/
350iFYWQYLmvS9b5QMhIHMlpuRVYprxGDU9vv7G3j3lRUSlDSDb43eLDnaLu4m5t
r7GhsBi4WC05WxB/Yf8LaZN5DH+0OrwX5+XsjvkdyIXKzQ1xO2TKD5fSHGmm/e8A
tQzCpjTtC2kaPJEVvjz/a7hxs5Fb6RVcY5CuocK/lcuo/zLMI0JkI97XB2clEkT8
12Utznh1Pvi9asJOtRcwDmLnn4vFzgU3Q97eLpj2/nNNvn+hu9mo0wxI0KXOTjDN
Jl0CILWPLtNBOkkQPFUMWJYcr/iQL0rfH0BokQDDn8Q+8BoogpBldneCU4D6dmld
1w7jhBfmwQBB9mweLwbpkabQyWzsMgggFWxYly30j54Q3Lmzn8mpGaxxmhRW140x
e8RplKjwJbNfsVsaV8siYYcfHnKiwmA4IpOzFQmOmM1JCYEDIeRRwvEcUxbaGwhE
vX74T/TjauweA7D+cgoSVUDKDN27JadrhgDF0I0E2ua20yrgnS0BZKR8+J1fp5tq
I83H4l5MV+BjxYBhbRa76Q4zAtcF7y/7Ro/8YRx5VQDvLcY0eFX6S/OhTzPQJT2o
v8eu800Opd9ZSVtV3ZfKkzEg4qmw3Rvu9Ufpdsv1ae9xW6nuhrB/qVzXDs1Qm9Xq
E7kDMJn/TU383B64M2Kova0FPHawUJsMYVbToQ7U2udGxQHSKEoRd+eKI99edvlw
DTE9Ac4UuC5coORVxnYShHgNi7pjeE5rjqtisW5b8edAhWqC2oZAyei89QdChkuF
NT/5+WmtRyU6IseE7VtVbux5mNDVouOTIesLSwndvPoCTJnQs4DovoWYby4jaH6m
WwOz8q7fASxLr8R90LfLDuaqvSAvZTubRtECdQHY177gSEgNd3c9nb3NJefteVYV
4fjprt2USrhfvMgH4umeFgdBZLkpKYv4VjTr+Lnp3UKNrGaHrCm+BIiNjLgSP+k5
cieahsGaQzPg5n/cRR9Xra4thFxKJu7hTou7NMQdKXJTlLARO3WPC7/fvy3qG8Ds
/ZRxd9yBdIB1OppnI6RC7969Hy9xxlqviRQW2uP/QZVCixaJITolqc/qxgfdbUqa
T8sONAE9hq8AZLR7DDC4+TrLZ2EFjkd1PP+5VCYc/cjA3VEPia92JW2YB6E693de
HcayjJ+XrsAegfEUuY+ZjSqNBz8MMTJM1r/dGPt30DhlT9uHVAnb/fK/XqkHs+Tq
VJN0m3hYh+fXnln9tF1tSo01pU3zZRnZeSM5KXtoGpvqKMNMNb0P5m+o3Xm0Cb3T
yy1yXNBoa2bYLQ3UkGipe3OksJw6aCH0Hp4DWKvjB0Z9hmYMujy7GatHYh0X3v8n
Hmz/OBkwqeRz27bMbYM8tREedQ9vYNqqTWxCaiqp4LwZiefSdNLPsdzdAdRU6Dpt
kQDqJDuQF9gTYvhNpKA3Sq2sByMUt7fy+UZHvu+7J0/p3QGX8risFatg2fuH5gqO
BwowuCdLTUrFpc1oFTjAfgPNDeTUDeDIYvZIQUnqEfOxTDEIsw1JHWnfLCKtjmyB
VQBhi0kT1PFo+YN+GTa13fhBw2mvK+wW3Txw4CpU2niE+kbVd43OgMQ+ECuqcyqS
+gx5yl0NjW/iU06EY+sVruvb0NFAzT6humHB517u6rjHi4jqe5C2BZumLKFSbiih
FO+qLrL2pPTEFqD4rEjsI0MPyfwKOlwkF9k1dpKz4wSzht7cdIxfi5QWDnaHPb8Q
4Atq1E/IOqM9qonqEcmHbV3MHBLrHyEaQoa2ch9ieRpQaTDwz24s0hOyAangkm6I
FLV8SOGifEFxdFnm7T/zEwtn1OVCwM0fwo85xD5ShJCCEVxhpZr6CQbv4zgAJOu0
V1p5DjLvtrSGEujZCvw2SyXfIh6DryRrY6Cuff6SDWgrrldlTwShDJyfauKACIu+
r18L9mxowpYW0ipGrr/OH1lX5UBX2n/5d7Sb7/fateoFecN5DbKXa6oBylnQkvpI
mtxe6ii01Gyjl627C7UwTcmzH6Rw/Qgfhea62AsHDmtTO9yluhp1X6JaQKbACNXc
zeNX/AR1CveETuwGZ/6eW/XVa9NuglLfw3ARH0FGeoClsihnb/cisexUqA7kTOVE
U0dTydeSBurxwRGR9YxbhO5kf4htWIg9Ic7tsHOD8/Ok7JM4XbV2UNcIh3jm6pef
IyK/WmPbCRBgh8F6mBFuzwWAQCMC7K5eecJzQC5Xjoh9HdbLoQLVhR7nYq3D/n2s
aK2by4yGjlP1u2BZR3cw0my2A+xvNt++dp9i53GQ6KjyXdCGAvV7PAAnEle2Gd3H
zFfisXK32OrGGxGy/p/lXWumhPnJX67tIghj1C70JY7vYFpz9oi/yd4mnMb44dc9
G2E/rYlopS60mzKw4TgPJ1e8Mx94MfhgqvBv6nJl40UifpIzKk7sFJShJ+1QZJ6U
bBbQga1UdOlWxDtTBqefRCyyHcK9HRHG3ooKl7AR4PKI64MvN0GGz5EE7FjaYE2O
zoJ/ep7W0cgbDMP1Jb9mKYmigkM9EAnYANOhvn9eRzgVN3BxVQayNnwF4bBpuL3X
N9mhHJiUSIOotoEhZKu7D/KlytpDCiNsvnub/Cd2Oi/VBTa3TiSo+QzEE20RO9+z
E/VNOvW1hppOz+RDC/wdpN7ul38R37rUp431kSDUG21lEPvtkGRzGcRUE16rcQhp
lbYtCQSABAXqDoie8+6mkJhaeDJ+VWPH65GRq1WoclNs4HmpWRyU3dLSIF0shF2v
kHw1xop13JDdrWGdDqAJqUoV3/S+bvAcZ/ebxMdGATInWR4FxHGvxMvfyrUxn4aZ
rzYxaAb+0TVbCoo8Lm3wyC/FggXiz5KLayf6rxovKvcm6Xcwvw+4ex8YtCF1HsTp
juYPq1h15uoMk4x8fBS73XctnBs8P/jwGmxf7dFD2n0pXSBJDglw6bi3T2VGGPc8
BnkL8JsptH60Xs4qUwVFZvWOnPzzDwJuAGbXqxYSLAtE6QDguP8mmIMuh8MxiIGo
g94haN37wmSUE4N3LIM8hDZ/hHSKkckfGRo1F0BPQ2O8rHfSFPpEufiEvfIPqD41
2ZwWDJdgsPCaeZFduatoP/JUTNLZ6vrfHc1gy4BVhJh7stmsFBq61d+XU4lS4wv9
DfNU7wTFttP0wd/TGA5SpoNUl58ZkgdhppCiF1RpqI7fW8KwpLwDVzmE1M55e72W
DC6/SIirHWXgv4W6Gt3R56cvkWDxgs/YMMTU7a6bI+VewLAHNiTcmXPghZ+3Gvw0
TNhyvZjzYrVU123uptp7+6hd7D66g6f4/yrQtHwGtTONQFbM94zDouKZHjHkMVE8
QhCznV+roQbt/9KcqEjmb09z76fNw4IL8Q2dWyeBIEmrQaMuOPo58GIBJAldnn2T
lp6aV9OxQvlEKZ7mFo5SGrim2PI13oPhfwfqm0hUH9/KrhPLDBh9dy5y9P/BHaG/
DE09I1WZX8vWYWggjUHX5Tva40++X7hKufU6kf17FncReKJGp+UZORCofi0EdKlA
gUpCQfH7rnrwycNRKhuStbOpOFzNH3FAB/LS4wN4YAyqHudLd/CoGUfjZ3GmGktj
sbYenMx6Kaj0xoLtFedtOdUayLSMYLH554AsV9sZvRZ9OWR52Uo9jYdBOHgp1CSg
hlO9ANBfvdPD37YAgAnGIArhnHbkpQrlu5jLvgZuvtrBGLRd4h6T7IQtWOoZH7Kk
arWdZ6AyrANxVF6fG+k8CjO33YNptDEKBqGt+hng0CNkev8SygGfbPRVZdP/OWCT
MPlRKd70UCnwgPWt/Qa10NSNffv+RMSA6D/19UWi+BhcBrFNsaMb9tlzkQzcNiAz
WKfrKWDVrpBuw8yIQFV2hWXUnIcXUpwTzwWyfn+Hd3LgAyfBA4iyHuRLqd50bXdf
w2umkrz2Ozl8jdnjBJxTw41ETxzMMsPkg94L055qYJwo+Pkm/EGKjOoVdKw89A9y
KMOq0ONnQvv+WhVKj1YVGM5/GEDH3DKYLfjZ5XFuQSiY2KNLPe4eI8TaNDH/VdcB
v3L5k6cEx/duowr1fEmIAL0CLI1mQ21HnN1uKFwm0iegPbp+oM8PX7xwv8Razd2N
Mvn5WI/zYOdtP916DcEiQStfaaTe5OcdT2wTWE9cnt+nEkpnLB+sVKYJ9/Xv64PA
fcv91nvDN9G2v2YOjv0xiKYKON+QqMfD7H5PUHg4Jpwa8WVjhj69WEN2eQjXgOps
cB/c/g8IlhwntAK3Ik0yNT9A/AQzAJSZa/xuHQp3y+Fes7xC9zPdMNDAFQpm2+j2
umHtDq4/VSTZ5HBxud5tLqkTxmWS77QAe+k5GYx//IpWeh5YZ0y5u95+yZ00dy2o
PbRWIBPQZ18oxmuBoQnjbG5eGSDJeWBp4+82cx16RnjUWKd1VQdrudXvc8HPM7UM
Ix801kl0x9ZeVDK5fsIUPkxwBLez3yqB7VDadc1sTkQ1I73eerU1Sx2JMedtadWj
E2BzPR7238OXE3dfdNb3fPZ71fHEVdMm/m6wHNMJcU2gR2CR78OKmwBM9azcj4Ew
lNKEVenv80TwDPMP11gMvZMuqC+4/X/3VKmNNQenVHZnUajxF61FcsL5sTtDVLaF
d9mP++0f916TTdBRXZkId8702SupHVWXOksetWqDEsmYIfSwHCWhfGpaPQrK+Kn/
9AdR8NRTAjHwxX11TptLbsiryaala4TJbzPYVp8K0PVIrk7B3KXgL/fiBhChXU5i
drqa+UqVw2d/fkWEgnDw5JUbW/P3RqWjNWHnwgVC6yRry29gJKQuF9BTXR5uZ/OO
tcQfHCr/VOg4mDZfMiJrqJQC0mUNMd9XqjJ5VhPVZAiuxhJ8brwY0ewFOa2pk47r
2ZddzUhBVFOXTo9ZFAkTgFjRj6eDe+bR+Z/Ox2l+ScW/xJE3SJQDSxeq18P1aDbe
U9htLg006HxiBVtgQLAGYrSEqxf+1XdmrFkI/LJrtUex5zgYR/2VKF/XapShj0nJ
wasGV6tTdw9mr6QBMBWkLlhjLCcStWNuxMTDWrah19PVrv44d4sJJ6ITLB7s10Ld
o8SLJcXRqyIxhO13Q3mqAbZ+seHtqZDEAtpSxacTVFZWUoNgfHhHG1yA2VtpIVOC
rbnet9a9Xk2BmXHRJ9gm/zJmrSSg7UAAAFFOKgrCTA2hRgoIdVA6EP13cHqfzeBe
BxXieP75ceV4PbWLrUF5iq5xHijaeHtDGpvOqHsj0yZjgw6qJCw0vIxIMARYiS7r
keWIId4hg7MwBSczrJQGk5/B6bFi7HRIc40apF1XD5mr6nCg2Fwma17f3YZhOWSk
N7OEdYdYgII0u9JyGqVemszdenXdcy0vQqZy+5hg9ync/WowiaHDx0F2ygviAerh
B2WPGirXxzOcXkvhAzeM8DhUzcGgWH1nWZLt4xKbZjcAGNR+Hszeb2NVDaeSLchX
Yy6uH8e9qmOEmUb7XJ7PFuvbd6+p9XStShUlhuLA5OzogpxIVdhkhqBWyDyuA/66
oiThkRVIzytBTBDbCxRx/EP4L6q2j6JvEq0X+qHg2/m/Egbp5barBildmiO+4ZTV
6IfRPFQYJzHOeib2Mcvga1n3Ukf0du0UehDrIbHOhRjR7xXxBDu/nEFKdIFbH0Uh
vTEW8nfoCrTppnBOYCtgbSFgSmdS7+z7PQAbUvKpwAtSX0u5Qjm999FyFZja1/Uw
U+VM3rY/sxLQCLNH/RUgxgqxWDiiMBHL43PFc4nRbm37VOoCQX6D1WRJObMppr6j
3N9HywS3rxCVP4D6gZ97IpVeJ1A/94BMDqe2UfIG2s/Kf2tLAp+x2pSwdaEmRFVz
FdQ5uPe4YXgnqsKyL+nGL21POkL/V1L2/P0u2geFdxP0jX6EmWucP/BP9nhuEDQl
BYb32YIrazD0M7uXRI3UHhzNzRSQYQrlKG57bORy0JeuVUqddHJh053hD5MrHU/d
cSZ4n1FxPKzz4ecY1PJrT7CvaMiLmzQQKEHanyE8ingmbtR+aYBGM+0kR3g6eYjE
lUn8ORAeWqoTYLiR9iwj/nJpFKHRExMt2rLdzL6EPSttwLO8mlWbzBIrsLPsVJlf
yEqB1kTOJA+dWmxIV0Di4pbNlTdBJYNdPvljcWfnazL0eyLS28cOX8fclNLOi0b+
2RWLkOqV6leoOlosKfxBfIo/HZ0MwBYFt9sKeacH91J/kVdV1sY0PBdlLJJarbq5
sUPwEC73lNmlc8hXWCSNbi1H30lUgpadJ7BjuTv/mNQPnHEBmHI+gr0O5Jbycc+M
+vzqNnQp4JpyxVWXjgbxyNtwsjfu3ZGXkgdz21y/nu7t86qnZTmo18syNiwwNAxc
XtYkAdj8uS6OGO61X1Auf6/BdgswFmrVCQswflcq5fWtyyWOCdZ0i5p5jNunuh1h
UUEi8laGZVjGi7w6/MwalUB8idzlA1Y3To+1GLj8Y2//ADvix+0N6kkLxfFD7JmV
6LXbBmI2XryGcwzbA02P/b8czO2wz+WtugAf4zO10W1Z1fLWaJ7m2pmaVqBBSiTc
l8rvt5qeG1Z3qN+sYf6i8lsY8U5YE4nFwZfhjAxqb+zLnMktWuTvPW2ZPh6h+hvj
Bn0YxtzkPFfCoSIYvC9P1T/8OcPRycKglV7VFtuq3jzlyvsU6M7mnRGAgzGI0Yxc
JMQUvu7F92mC9td+rA0lxlcXe9qEX1xTrzQmUSIhZZM9Z2NXfKAW5pQunvOijo8t
47puxXMXezwaIure+XR7hsOrV7IOCn/M7mEYgu9PngbVseD+1NtQUX3GXgJVB7NK
cQqpsDbLR9rvla+cUyy9Cis3DNIqvqeFiamZTufXuFe2ERpjcwd6rw5wJ/ZRNqJe
6/YnqdyeoFyE/a7QKBIZyZFmGzJM5VWpP64mABcjGOMVZgOrmbWrUSmAcIqqaXv5
0ox0+eiORpuHe+shz73QoqPEzkV+Nd389v6R1+fuVRgTfTSrkf0YGpekkrRIPucq
fgRndPwz+unGl1MbdXe3eu50NI24jlHwBZVUkskrrcT734eiEGNT47V7F6GCEYQH
WqC+CLParuMOsFOpgmGzgBLp4wFzdYtU8+MnY9aRnQId8/ba9kZiBu37gFSIb0Bm
PUFNM4/m7tWuTreaY/Ocl1ApDWXMmlUZx4RZtvgL148GfL56KN3V5aLNzxjXGOjL
+OV9kVusu66U5jcdXOb4uId4MWGIzW+SACaMt8l+w4OOjTQPK92PAVtnaC+ao2vU
NgmFsbih7rzcyM+orvqNzVHgBWglYMWfY4Nl/nQjEhz1QME87yL8rpz+SToOVH9R
2fccnhsEDUsBRIKIINtVn77LgFQ+fcHbLS97n2BoNP/IoF/Ys5d21bv1UQm2x4Fi
dlP+KH6zQhQ8AAVHQJCkhilxUF5WJoSje8kQtkr5nuc0ikQRxvaYp5O9TKETnZWc
0es0eo7oTljaxNNagJNDCkgxU3p1/kvzwJKmfloeZuBLTyE29wib6cw0vu3FElW9
d/PrqR2QUZrCC+hLauESNLRXHZUFduL8I9f9ju2HJ5rczRX+YlTduawa9QA0XA7o
R/IR2LShhksZx9f0qEjU2Np5c71uZ4D7SvuQ52Wus8uyQ98dmFbUYBKcndOptg6f
Gb8wcb2NhSggovN7EExtgWgVDl/YLvAqoVykQz3wKjzu0Rd57Q6etKE6XEkN1aAM
qADkYicoLcswgxjMnn/KOpGbZeOPjUyR5VJfPKHhYBODQYMBoum9/vFPDVPK+QoX
u9nznzAGCCLngwZekWtfP4JVeZXQF1T5AwUi63IMhhdyoOyqUjbGzr0L2ZXRVDM2
gr7Dt61bo/QLiopmz6IcFKin9j/cF7OuFN2Y4nERYFLO7HnobZ+H3A3x5TydzsEl
3DrwffQETfBPBgv8UX2QoFgullOPM/2DoWf1CkwDQ7UZqkMvU50FDBcrI4ASfUpx
jsJ8FKCfvdHJl+mhH8U/DcVVNV5iCua+s6PwezixsKWVikCBZ4v8LvqaLKfxuthU
/39MSW/ZDFiH/w53CCmTk9K9Wr6N0JfM6Br7wz4PhS9wZkGHRadQrygt5w9BxZ25
a0h/FNijOLpbdV3vIcbbor4ytlF6+uGrvo/jqFmacLHiwCj8tcQAUrt1kv5jMcX2
Ouq20Nq09D0mvF/0GAd5LQzrIpavZps/WFBwW67O6EnLdTaDXjJiYZQgC1Jx0YCj
TbxkdG5ZfRIOfZV4XT0KU3RBzQNhgrv0VEwdv6d/v7mvvSBpotJihAM8yJQ5mnh2
QmH09odVIDhHbXh9yP9IqM/3LpJBfV3Uvz96bJ+eH5vJPaZktElPXkkdO+CiZICN
bUEm4vdrQaIPszf7uDEcCTosJmazKdMvrIe0haN7BvmvGYWLQyUVMXLjpZdAVYhc
VBImQvvo25floW+K/5iTpZx1I4cwi6EwLvY4zraqBoVUkJ/RGJE4ON628uonKD67
oE+FS6hvIUvLLOdRaGE/BpWykVkw9E7hrfrWbN7MhOixgCFQ7YkzxPt8GpvU7TiL
`protect END_PROTECTED
