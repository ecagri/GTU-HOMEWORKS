`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cJ0+povgZYzU18EUaPjocY2W+hW8MwF7sDbXIm9w3HA7w7Gnx7SYjHaRRwhlEn61
AxGH2fsQ2MC9X7WISkUKZgNEsa/sLYbXtfNj02KZDqe+bXvyC4o4IDY20HAC/KAu
/XsYXi1nYlPpZr/R2dtEU6FyX9yYNs0KYFcpoy6vDj8S75dR5ozm/rMLWI8E6QhE
vjK5S6toiozoOnn59nL5VDHjpH/4b24Yz9BQDDdjumup7zDnVlhlRdls4cgFFPgi
f5p8JzQ74LSAItcAseQjCmaCUtkRlDix/lkZy53Mk4abZsb5rOy0NYndwjsnQIXU
UKZ50h0RnYYenlhgp3W2sjSEni9fCENnyCW43+YpU6ddSypyqcWXw3a31q8uIXmB
g6kAZuJdUAXWr8b+0aa/w9iA8QAEzaDQcz1MFS9kA7g09UZvZDFjkVK85E5ulqNx
1GISZtcqcOHs1dB810gG6BZLWx/uWjTdQB1S3498hBeH26bvIqoJMwI7s06eFGKl
1+WYuHRyDCHNw8jCsAmFG+Um5sIiqFZP49873vkQqkZK6x0yakC9XYDvxxLgZBgt
YYpX7EQJcTwc2u7vJSw71o/JjzEfNQ8bnsj6A/eOhVqDluh0yTLz74M3onzjrpfI
C0KrnP7Kk3Rlpb3VxMQ1UmUolGU+YXOEe7VxdQ0YfkdJwoCObmHS5Z+O2UxdeLYa
61SxVk7tqu/4b5eHOf1x5wxU9AdkR87J6FJ6vbJsgL0Ws1COPv3XzekwYJ5TiQIC
3YuYx0fFdk8Hi+oTx9sM3Jgpud5kgDSvX9yp8tnjoKlODidmjkQWsnmOIfwYwhWk
+ttthY3uajpgqurCmWHpTG2yfUnxevigUp29Ky6HnlupNdgn5GTANJTA93xLysMo
P6+RwffjrdA/6Zbg32OYGcuw1kG7PTAyQXWyCmbK0YxVNHqIrbCfhjOcvDtYGBgd
P2laaoGmvQlDhF1/6X3LXS52tEIfmLy2uemXpbcAD6Fhe59JnF+ektCGA7SATm/P
JDOX/cP640RJHB5ymspxNL2wn9b/IUWnZml2WmSzojBBqkRuCBpZRoTel7c1lS/z
oNwAaFQy3KwP8me3lzGwqKO7IlhTHtHJl7A/Ao0caBM6V7RHWZKg4yIGf7fHBoZj
MIxjE5b312SKFHl1hWD99ZfXrNe3rks5KxELG8SR5r6StoQrGxc6j+ePmWvS9ZR4
LHTVHiYFBw467JVq87vUEAwPiLp31W80iiRg7bnQD9yfghg3Lq+GuQ7NfKCFH/BB
CuMg2n2CiBmy4SiXL8F5ASiLQcEGpsoWjyfvXHs+2/7vMEKZYh/myrw8YT5USuSU
SZlb3aFXbUsDxr/W7FQ7rQQ46KXrOaN/3DMpMutdwKGKQoNS1xe3xCs4vT8BWI/C
mN6f6Y180cm9U27aBLMg+JNWdpj+sanKDFkbrWiEu/eQQUikn4FvU8buspPSSvIn
9AryJWop275KHJabjqAA4HvHbg1TgbwqY/TS+obIyKxtea2bPM/I0Pprk7ii0WGQ
iqnZWV5TH34QpD0QYqKT0cB4+QVk+fsgVW2drK8jEZ2JMyP24SHzxnAZmQCHRzjK
fWtfobQKdqMl4mMGgZZG0ZLa9oib6JpS+Ese3a6wClWZ8vLpOJjyl6i7HCMhYohL
Bqk2DFj2sMbKJT2n3JZvIoI7IWkf/dzupUCJ0DSF0YhYwkXLIfi2Pk7hnAfx4nzA
kWszOPiUyKv0SS+87YklY6anms4dDS3GR/OUedGRTdbDLSLKVQ9ugLAC31KpUttF
QhxmOJ8+fs085TFa6guHNuG2qimpM7x+LrwnPkZi3w1cxiinKqKIH5F/qcuW/mgX
TDkHAMxsxM32RcuYqjbh2mhuO2+aamby8YVXOOcDBUR85EzVnki2eb90ZUym8y/B
CDrFm2a2dlhOR7TKy0C81hWB4zqUqleKnsuqLJivvwZ4pSVjwtTbUF4vHysjQ7U3
LZ+H3adfPhxbGcTGqY7CA5EmFmGTyxpzOrkVbZv1ZIKG3FxyuGmQ4T0a+9wM211W
KPr2VFSVSPFfMjzgp4c9qvo0MNHM60T/u2T/tMXuM6sr0sLgLlOHH/z1DQbJE5Ot
LXQOoiKP3QLJZlo5XX8B1DEwfTluPoCu/xOkz0PhiVZaKjDio5P91Bhb0dLYOaw/
9K+B7Chn+S2LMOe5qf3uDUosFSyd3pAfZ+YzMNHKczwoFXrHB1bFnQu4uD5ybTh4
WgQg6U5HwP/LkrD1dMVNS4hGddBveKFHJTMOAvkI5yMAZQXTcZkx5iBg4M9WZ+ej
t0sdnYTR01ocB1qIC5w2YG0CPgGgVv30jTycKOkpBAx/1TRvXx3HSOCcDDfPuMo+
IUDhbl5YRc1Q5gH4dskaXdAYxipvcdNcCb/pvePhGlbQTaKtM92PFRlGHhwK9ukx
TylzWxRbYKYq4Oskf0myWrJMmbPSSqpgtaY8hvSz9vOCo065e0sl+8Tvn1T0KDci
SvcTa94Y00nk1r8obmQx2C1S3L+Vyd25N5l2+BSlJ0Z3h/3sKjoQJmAOcAyhce+d
1Wi6P/xiPgkoayMwNfLlKnkEkULrZDw0vm9YUWphD/D3zSfFS3n8oN9U6W9pPib9
gDf6/oKlUbCxNQ4KuwjpxEiR+P7BeDeRbQzlo9VaSewCRy2WtnVYjdmlmFDJTggt
Q46F87H6S347K1HGlC/J1rFr3vepBxp+f8o1XLdw2J/C5cYsBj1ebwj8nQxCoFk/
LVHEUNMDYrqCyVpcKM8KG7eMca6Alj/JMrf1IrbWwQ14jslTSbHHMhOu/f7OCM4l
q7nlVoQeKVE/EYfq/AfLMsu1FgjC+r3Qxx57dd29RD8PtPe8uzr1CHmL0P+fTtA5
5qGGMBRW4vbhkJ5i2sCiB8WZWMuthQlAwuIZeCvqiDZr0VeRaoTmS6Bclf4W6sm4
csDL1qKdZEySCCUghkOXX+deL/74wsgW9YQS5LUU+BpuMepKd0JIcU07zjto/VX+
CmRW7QzaxZbgc5J9JY4auqWE8npQWUEomMBaMq+vMGUtSN3vB4iozhwulqtFaUYx
R5o1OeZFvx+W+TppgaIucXW2AjTBZhy7vEuURzwibECZXZRZpVP80JOnizXe/REe
rwWBHkxn/s68Q+YO2nYffjoUHaJdPM/AcLJd2XQIeRXNspYYLm6EBe+Oluz5CF8w
HyD9Iryr0ojyhcQgTb4ib1F5tnc9GC8EPxSmCC6YIpCxPMwlwtDIB6Un9iO8fkSO
0KDSEeKL5mJSbMStOfxBFgG7j/PUry1hppjmIc0WreZz1fTGvAmuLUZUz7uN6+lp
58qKWn/5QyG7ox9nrgSWcyQ2aY0vyRQY4pg71fWoWNC7ZjI4A1mt8eqDcJ+eMq4Z
+0yMYTIbdKRSm+V6SgScwG7Bow+UsdD6whLIIKoJ9/Zel+n3wwawij5WT1et5+vp
Dn54MiXXmFwBsgv0xlf39gQoNq0VmWdOSLRnJJh3cVMrXGlvA6FJokFgAQzAbesH
Cnuhw9ZiAFhCIiVTY2belAxZQCOgdzCAk4vEKgZyt17HIMnIxYyp9YBa/zE4xGpm
Mhc7LvzdQz2BD2UxrydkrPlKwsUlbA4BH3305fTLg3wS+GXSwB2UfC60QF3ZfyO3
+fVPxMsG1pWOdSZG4Jr0Ta99isO5lY2yjUhKykFwZkMbN7aYl2BR3k/0rjM9e3tZ
GLPIq+piqR6+SKQPvZTtRAqr+GpKnInV0mL9R9Aw7EKwe3HFTok3k1fG5EXvTMOA
rZy7XmFKm9FDEWa8bhYSoxSslxYYkKHJYKCaxQ5aURW5zmAPF0F0r0mqfKVLO58B
94cBgNIlr5xBa1CJsBuvCyxjWdFwsbSlu1aQCJmg1ci7lC1Ih70ybGzm7vXx6l9G
e9UoEy/gZC6aUKsHAZGNNvuMi8FtIWxZqhgBgjf/InFzSzE9/FU1FoRJJQdCN5Fd
npJ3qu0fAK9xqenkmPKvkzf9UwrcnKvXCtu2fO7EkG9LT+QbE8oQ3CaGEPmtKO86
Lu587NdXuAyoxLZlA7jKULZcz62dQuTW7oh3ZSYc2y7h73q7BEChNJraBz8H7q6+
Hx9FiSKE0UC9vd1piOIChxbY7CFkKeL4gCRcdB0EBw0CTgAPlGFnS6AKwZwASPN6
2bWN+oIsV3CJkoq5eU03adZlvCqPXvNS4dkMOfU3mLSMKWvXfr0yhUzYYPCCJC+H
9QbIqLs/l+AfT96gQEwQNWoE//1JxesWJTLu7kto6ut+FEF3MABLKcwZjaCsm37q
QQr3AjrML2A9zjB1obUJelhgyO45K/ilQKQgZWVmvFtUj43HRMG/5aroQHpyZSAC
QV121bZc27ypqiHJX4DzmKry2aE7U5beSMAq2sjHmWXQsSuINn7pvtCRlDTNXmo2
JoUFb0S2mUeK6DpBTp9tC5F9V4E34NymlAS2o1apPnXkmuOkm+CI08DfM3aBS6hb
K6JHoOuhavyqTgaX68jV+pSkCdt+9x4mkqK2kJMzj6nY9Zl1/1aj0smkHBBlCxIx
IeuetVvADKdDdAxP4ZnCDvRyzYzyHepmULu7Pvw6HeCK0/ZBl4n5ybTB4Mj1P5ov
84ivtfTVF/f5urG7HJqiEVim+Tg5zu0XtBvlasHw3waDPXo1EME1BlUMH5LI7u0n
GhptaGbs5kf2fT/64ZMOIOm4EQjAyUH3dUrDz/7Uy2F7Me7Ss6z1t6nZVmsa8Jtk
aj4BMAKzKTkLhNGSJpAt/3sZ6+Q8k90y1ERFwB5YTQjE3fR8k2XlU2CPLkLCLElH
jshPqJrihbR8BblClAlScL80FYANXNn8Xxe79qpoCRUVEYQytBHhJgAaIzxKeWv7
p5jTgpWzz8UrUeU67elRVdL5tQ9CNnlOIRP/wB897Mp9cUj35m4RIbs0IPrm4HYr
XCMJ/jxr6trzLmmQmLUAEJ9dDnw5b3iMP0o7vtCWyeEoCGIy375NluiAVP36Zw+m
XoYPmHeWkXbET/+NYyUlc/NjHDSwEF/qazInQGlkuzK2T+rlKKxVOMmlifufydnv
z5J1Kv+3/ZuNIFsB7y+AFoQA6LytlSbU4p9TwNFlT/7H0TQQbj4U4t7Fi/2VWKCC
E+khnHk++5eCQjGd23nfGnCc8bljgtggVijt2cNKauZudazsk0NzDdtTayfs/7YL
Y4ffPMuwd0LtxtfgWbPv2HegDpD+RWEihaSCrZ4J1+ZLXFlIgNgXkgEXoDtuJ5vx
kQ7x2J0e2jOQnuoYcDSCmnb8YGmOjvQTiLgUnbG2ppOQPiDH5QqEOZ06xa1BJosV
0JwcSDDGWL9eBld+6v86j+6uQ1x2LWpXufJVfhGMrWSmdj50eRvMhYFCxZnu351R
hbWJQJ+ufxSpQlePOef9u69byZpeXHzlT+h7aWp4ffk6gcRGg4PbdZudll/5tRkQ
5X3FSKkK1VW9gTMYEhUbYOe1Q5hvijY/9/UBI4fZxZldigcD/L0zA1Y39XqlVY9X
eXX8NEhfWuTdcw2X99BsHUPEYD3gBlsvhE9nXNG1/OrkuXVIQ3toJQXmIKfCiDm7
qTUEVUIH4913oXenc2suK20SixAv5E2002DkOSxMrCW3qUuAtTYiMwHtNsISoEEi
SfiDcE7sQH9yHyhSX0NHObTXjdz75r7yvC1GNtEaNQhSOodyxsiVfE86a6XPA0zU
ecHQ6WqnDtm2KQfSMOWXr6OAP5zimOn7BDzUEXDSrNtwC9bT3SP4rXlQWohrshX5
eryGfhrS3D2LuvJkZAMuhtZS9Nwa637v4WjL79g0k5YwMcQsA2wj7SvDJN/jVU4e
HuSufA/0Ptc8jrNryLmLzVpfaJkIbvEe4ZKr8Wr5yPBOkMQAs+qlnhT8rQJgtoff
ZaaEgrAqSLMCRJnS0wXWtZZNRO/B0aOPxmDS4aylFEES7yN17uMxHciwnB8ar7se
AD/FvrCPND5b8XHxwCCOyEVfOxpNPDW3zb1QdYsiyjkSEV2ema/f0KlvQAiSz9Kl
Wx9Y7PC+kTHbQgHbu3HVfI2Q/cycHe1nI9XKTyCQZOsW4dfWFqCBRW8D311KFF3D
oxi7VccNbqPR5Voee1qM7SFPwyj2UfCsgqachqaB3eD0b0I7w1ur5VSOT48z+Gq4
w/Ez3EiXn13vvBJALQMfK8lY2UgGStVNQGwMU84ToHuC4MQvmIrJSs8JomHCyPsR
OyQIKqE+r5wZADj7uZsX16jOv522vC5/iQcStYU9GtU1yTC19pBY0F7VPzojbmQw
65LbSgWfGGrdgJpfPfx9cRFGn+n62Ca9k8u7f0ljlXmVahUGgwJL2XkuU7ugdtj8
ZeydiOD3SXiDrLl6bafDi938aH1C+EhlAUr09vsxab2fUsAGKDyoCbrh7eUJgRuA
UI/WWVSEB9ODpJOZ22RElW3BeM8yEyg7VA+shjcbLa24ynQlyZ2P0JokA3nXSPFR
342NWu7z+c8BqHUkfQeeJhmg4kb7wVVVKY09U+N8j5T4wAkym3gfeleZQBblw4qt
/43J5Lal0N12/DrbyxkoNgY5Jo2qwEY0Ejtu6UVMHTwJv3DJTO+5dfhZRY5H2E4i
xljUkiP0u7IFN8N35tiW0HtWfI6Splxn63WerF7lCuQ9oD6oBah3LGWEZI4/ptfA
L05OY3aODubx+bRnhBuTXjySoAecr/fDAnq+kzgG+hNcjVTgxhIi0Eo2GltQYv/Z
LGxhTq7hHKROaM71Ne4ciF80xEeL9Qi2bGsvKqZdp0kZ8eZr3yEGRFcwhHbj/aW/
MvFfWmgbfvgHCJLcDy1OanH6Jh5OOxM2/3Hc65wODL347EtnkCSnLcMxvAes+Qi/
INIH4pUoSo5ZK3eixfLahT52x0AAUHizyyJJuEmEmnIPCvmcTv107hpXREJaPzgp
YajpsgLmQZezxyiapir4dLyYBSf0XfNeucv7SK529Ql/LIF/gj5BNWWGPU4sFQME
bL0PGVhKmaijmXqZhFiTTILYZt6ZTj9IxRv+ScIpFJlN1r1xLh95VGMwaWLW5JwS
AOmM347JiFinVANQHGayunIbBkocZ9EZHfjR95y7EJrlDrARSL0Q7E7tCMqEZlFg
MnUqwyNCT4hesJVCFZ96oprSvIJ0uxQsNCOf4siF48sNyWxiKT3OVkba8edrHd1O
ezm3FhUy2CYycR+HsXRfT/6hpo3g/6iBK0M1WJvQ/zUEoLp9euuH84YV+8mAbl/j
pmkwkw4qpUTolyw981AcC9dRsI8rZ2KQfyB4v6wqX3Xe01yDJdStP73hPEQzF+qI
3F16RTzKw1K4vI19R6XdfYXtDPGX/mHhvwQnZH6j9aH8rmOuUdsraQOipXYvLW0C
APEgEOU48XjN7K8No/BQPADw2cmh3NjfiTbuah8psp+AY68WCTsRs9Szm/Agw/CE
sGPxELWBJVZRFIBWdg8D3Sy18CRm/gVfgtpx9hXAjtQROIfPC2HTA3dAmpTwn+cK
aBseTwoOjz+5wDqh0mRr1chf67E5r5GyCEjmhTRn5fdOXaH1/6tROdGMxm/YGvzX
FrgTuQnQZFfmF6L5OmMmZMI8j5ADYOb/uCiZvhzDTpsDve8cGsq3TqunUDIIygOw
YDZbi55DP9RMP/I5IV50wQA89KrwiO4OOej7nJEI+MVyApWySzZpgo0MHw0nQkgg
gbGPcN2l6QRela7l+d7FQpeDHiN1VYve9KyMH2Oy0qW605b+cMtkJdVIsxaaTVM7
mYdAsVfqpmUnUMrpBrb+vOVUS/FikFfaoDSGHsvG1VYhKxZ92zX39JfNMWzjlo1C
zzbIsgnQZaia0v8ptNaGXnPfLfxvN3OWhvdqjWGsXcVeitOtja9uKIpUeeQpEDyS
87CXoPECQnSdOcMU9qKsgBuAys2DKtQgqvSjLZZf4Ide4vYzIGdQ7ZV0J2UMXC8V
NF4P39OAmvQEwORv/YiXbgwZeC0raDLcp+R35Zy8WRMVrQ2mrJvMyL5hO879jTlx
jljl8VB6fdFtdFxB/tCmGXxvOrEnRm8v5/283+xWDz+EQS5ViGobWlpXRI/A8QOL
k6A4a05xT90M+/ln1EdCHwh5Em7yy7513pewLB58R5a7d7UHYzv8lEnd4i+ECUru
v/vvrFtJ24hnpYyqp7yh6+ns9YuFjxYcHEuN0R0ESBceahVslzMiXAiCTaZMGVR3
F5Ff3IKGgykaUhI9lHhSG/oUTluNpVVknUt8nBI2W0xPMCk6VqUW2liZXnnyJ721
CieY9nhH0IjBn4dKQ+e0+1PC95K95awhfm3NRFNJ56WCPisv47Nc2v76b1D7MqiF
olDtF9wzCbz1e4ECEgvDFoYHq0SgeqiSlwaoA4hoF1wHhS9Qf5YsI7KhSOvphQSa
NlZJY2wcZ28xuW3sftNaxtKA0JlPx5u93nCm5FdyMKL/KFpktTXaiFNKkz7iH9Hk
BfGq41ftvdOlF3V1AeVNfzRtb75+t2SoCupR7cFBZ8IDx3L+wphsXpK5TlQW/NBv
/E85iTDoNaB2yb4QloWYyAuFszS1toQjxg5inNYdx+rBpd95OeAtHg5s4GU+m2qU
iU1SSwoB70PvjbRP/pxy1usxNd0YbOcjMfBHUJspyW48Bc/nmeOgp7jcyixaPa98
sDj4D/pBf95sg88VOekKNSchimDDRGUFbWNbH9ShZLzwpFYJFwP/ItQeA07SfQKQ
xoWwiiNtlFxydLWI03eSfLoHphgMUBfUeNL9ttYn45a5trVxwSJkfAIBIkfWlPwR
+N+Fh7C1yPvzjxIO5uTqQq+oRJjrxP6lxLkRyQL3Ot02+926Yobd5osTeyUnYS6a
B73p/avr4urK+vvBP0EtPpamytJ1KhlYTbi9m/V0oX2UqNN3SC/iLhrIeToLAQbP
2db36H2El7fwXoy0oW3R3sfbG/Kqc9XAbVF8vBVGj/qnL4haqWNoe/6Yn2VR2eYD
k7q/K1ixQh0nTVavuo+Q3SwvcufHgyffm4V8tsCqdOcLp65F6qBugct54rrqixtv
b5qJ9y7VXjVAlfL+NkGB6RXkwVgxJO1W7UyDv4+xJqVv4gwZ97oQ3jfPfeE1cKhX
nbX63n212/E2fYff72nmy9Y5ctlAzJi6a21xPsVcRSyEQ7EH7o5r9u//kEb3/VG+
UEw8IW64PzdyU0WFrmWguLBjODAh8VvzWcYfAuzPb29YbmC+m7u5l8ZKpofAbQYj
pM/cFDfTqAhPWsLXmX+1uCQcVEliusmQmhpONyYjn2PvmCee+VSjz+CDyT/7/ePp
RXZVUqg1WtmEAz9ovLFpFMP3ori10JrfQXhbUJLoSNwMFJz9ZAc8glDt7LabcQiP
ugP5TGPZSmrQ913rKNHqWoJwdnW4uaO6Iu4aOCos2lB4XhlGEg0xF83DrTyfEWMB
IuD9B1N36dIdn+EK0Pg7Gmeu+17//3x9OhqhggmtINDiE4nyzALg4RzXTLFI1++X
exjeyyUjF2cx7ZBwzEsylrrld+eKQzMceXgHZyWSKrjDAPLOX1eGo+3ky/YdMVfy
a1nweOlehoQjD4ZmqMWmm5hu5lP4iPr764D9BKn4ZMtddY5msDhzNuv+JPZc6hi8
Yqc8CAn7iey6ecyQlbmCp6BZlEv+x1SjPEsZSSqLTKIq36AxYnpU2aLpi4mm0tIh
bxhG6u+XzqoETmAq9n++aYPzDdaxifdOtI7LPczEJBP2xWMRQflHqoXExi6aWZOj
fi5OsEsWIHQn9r36aAjpf5rv/H2kx1InQVcJ14MPGyAHYgGkFULBxKJ6ps0xrJLk
36fQRii6Do7eZs76LWoeMbby/b50VflQuZUdClVHb782A0jiQKdkWNbh8hoqNhcC
CpstIgw0M+XMVN1nOKhQfZAy0+hxzDkmHgEJ5nzheImVYr4gY87um/3/f9hgUJN/
bIcCkMoWY81KXwLngTYWuNPL8oIMZO2EfrgyegPnv3anWc8hYoCYCaSPpru/yxS3
PYHGZZ0wCGXwpbtzbo5nD4MpF+hUaYD4TsbwLbSxVYknozrfDDGq1UXjhO0YU9xf
SBLunHTadTWECnsbWMGKQvcj21XQ4xYnPmWpe5vXYPGuGRfRoX73EuyQRh3vroRT
R6BpRDqXa77opOGXGpr5K95RXur8gf92uO+ZZpxf2yUWMv8JvZOb9S7PyqlBgBQF
YSFmLp8oEXfjrFdTuWlFTUe7QoFdwg5DRL5lQYVU1czsrLYbWIbwyL2dXCVsUoAO
xFxso6NbkLCSV2gjZq9YM+P9npO/ir7NsrHMqzKr/1aHPU6qU29aI64brMXYV6uh
eq5s/TYjN3UDN/801SfkSYzbUgTr6XByCz7Y9mYT2Bim554X+Nk2FEgqs77hbrUf
Hg3HWURpPmiJUAL8fAVG05PsIUPzI7T80JO26CgNJKT+kkmubCCvbs00FxZQt+5E
qJBDJRdzAaE7Dr7FJ1ziG63h6Ba6VwIUOO9Z2RYa5nBUDc8tX2vvdYLZg7RQcda8
7ggO2Kx5CaCT+sXZ8beXi44lgQ0PO3Zt5XfNS7STt+Ip6MMMUn9KM4zmSFjhymmh
wBo1nZR579VW3r2ZUihf7E+gVrcVS/SDz0PGTKSiUojsgiByPK+cNuzAheqr57lF
hq0u7G338a4VSlc0+qVM9dWt7lBiEF1oSKatWnWdmj/j/AwfRdeyBCRijGPsLyo3
uMmqO8ZEU3mdxgOhEBS3hBXf6rLHldeObOMeTyHiK9kyaHGi/QG7+9Z+LHN5UZuf
7BWeFqwa05SJjF6Yt5LZUw==
`protect END_PROTECTED
