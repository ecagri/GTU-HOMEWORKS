`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6M8iYTh9IMxVOI/eVidNaOK8PE7uyviRraF2DylggUsZRicuWI9scwPnerrXOLnP
mUawrZ3nRr+Dj1PrbeczfJ+oWXMotT26eDhjwWvvdhUi77z80Zjcsy2WwlejjjMH
8/urR1dq9gVx75ZbmhYDc6cxy4L2D8O1YpgzEvezRvzI8ZzjUv8o+tChH9O46vhx
X4wnCExjWS6t79OhSORHf72Dbe/QC3ok9rmazW+9Kj3DCxzNLqJ94NelwpwZdB3q
Q0ryoYVusNwn6R5anjTsMVABQU1QdVcRAK3+Md+UftpNzhrXBtYT2J25hkvsYcNq
JBmo4MjuIYlbfXKMdENH79lb/kVVZNUja8g7TC8lPJ/GsSJfMHuVuU9qVQG0n7h1
XaabYb1GcmIk+HzlYMDX2yaXuB4NuhpmGfqLcawvzsVgSqVp5DK1Mo16Zt7d3JEE
3lq8QW7V25EHqtXOs9906HEfYip75XKzIx5N0d8vhPriyVoX3I+xJfCqlf9CioAq
CdKg0xoH+ropQXJHvLfYI/1G2mHg2gxgs+fWx/oPYfyLUWLn8/HDCYUMDA1+j1eZ
BCk8AhXg2GPtwQdavfO8OIEKXy3P4yvAQEX1vJeLUMOly3TCN+2PsAWPTanLnHLg
lO2K046ZWDXlbiwEjAdXd8ns0kR/0FjgGYXwzU01BxeFqwF+fblS3bb4+WoOoPF7
5m0uWHwZI0DQ+9JEooWS7yB7oTsR2X2XJHap30EIioMHZXpBdK09vWb/s0R3sePa
ROTQtsJYFpxScLr4618OtsjmN1qyQ/tfZAwPsAJ88U9GHhnzBddFGCVrnEHgGDiE
q7FwBqQQ3FLi20rWOmoY1e20FN+6m91ojgjYTFsCfYU0cui97D9TWSULhkDxHU8N
h1zZlPZxvX1Tv1l3s3AFuYK48C7y+RrAMHb2xcV/pQ3/k8kyiugJk7Kf3GpoTQKJ
F9v8ti3Gw8Eo5P2OA7nM3FGzWWkCJh1Ct5Ft3ax6w8/fgZp9aiS6423NoFhK5Kb6
pLFAZhiNNdU71DTsJBVIZxTZ3lMF1Yx2e/K+Nw3dhnBV+mdlk9hrZhkKQwlF6Wcy
pF1AvvrYOQ0+/Tv5DrW4+EHk8tObYuCzRqhrYjrv0aqWVN405YdL3+TaoOCAXQ8F
i0mEzySTsD4MsRo0gss8ibjDVxD/bw3s48mvVhn6Vooiina5zinayvXNhqeDEAUJ
Nn3hcZXTPCEBgOxFH6Yt6zSgNmgNEpfnqhFwmmzWXGgnPINp1gEcJSKEH85J7UmE
CJ793tu0hUsS3jY8+I1I5oI4wa/2vmkXqBrf9VoA89dmUJ9H9D4ik7veo29Tug25
uxj/LHGR3jiHpI+k3sMUXJ7x6rjflG13G8O0FbtIVBuYIwAhxri3iL9tK3csGd21
r9X3wjqIF5uNxj77XAYnOUhFnPqD1BkkTld6MWeYJpKKHRdNXhzfHaHHO7fvm9TP
v5YQFbCs8gARtDzDCNg7laR0WAaiWubfcVA/wnC5MkK0kIgidHd7cKh0z21vjXYE
70gmTcJfJRQOWYYyMVr3CkIE5hT0oqB2w9ik1EEqGET4iRBiL/ygalGajrTnXSD/
quU8o1IBc2dletl4AkIvZdV/Ff9zXK+CaC1WK+SdOGlucBM9Xr+Zm6Jk5OxnAYVW
vKREAMc/vvRNuFZR89l3vR87CfJnGxmlAyxMZtXR5VynxX2zD2NI0iZ9W175rxEB
R2v4ZnHrrR83YyRRBPAlBYu5PjKsADZcVVllhXn82gbgUxugOVpEnMsqOEI09bPF
So8+msxrQilfcwNRH/wsQHC15bXDRx7+512qnvLCMqtX1NHN5bevlNszk2KrgC4g
pRMP/fFj9kXu5zglu/DeqhQarDizmSXxfr8YZND7bb9iC17LqFHs2P+nqvXoEzOy
uYRiHYPMWj09FqeXYuslPuZmVytVaTE2ik6MaJUUi5u2DZ/4PavyOJ20bKiIucSZ
8BFqiAcZi8lJjABTSped6WAi9CPpMUmy9h3dOYPHnzahtbgA+tKUbOInCFITDdYO
veCPSpLl1r1Z8zVzL52uYt4nNytn+mQeQtkDQ+ID5aUDFqKTfPFMV/mf4RBCl/zO
HpNjy4At0lxjgk2yM7dz/eleXm87g4ugmfEqy8CTwcwiCSw5LpahTCgHjt4EHIKX
Ze/lZGGrGhLX5AocFx5AynItcc8TKq26LvdNC1ziZyMpYJj49GgNpkcp/H/q81Rg
giKH6tdWT7Q1QbCnhnLMFxc5M9CmZdnnzWsEvvqs9S9J5AI13j4EV6yagSBWBmem
Ku9fQo63yc992nYgRpt0YgfASBvXDulv9dwqC8deKIdbu89OUM7f706Zhs9JHBtG
fvMZgze81wRH/FC0Pk28eioFGYGpbQyZbeSIKtNP3k4tU4aJtjewqeoITsi8K4ew
IpXjy9ZwdIni4CCLCIvv6+LbhxhEVj1zhGCNC+1eU1bK6CTjf6hfvQ8GPpLYPsxH
F7tDIM4l6GsGjpkLmnE+5ODZ24nVPc6E2rWnKngEztd6G/GWcUcwxSmywSsiVH+o
CDzTYS+jO8rckFZJaMwDf+Z+TUqPMovgS3CTbRe/F+e3kbGRUIXVkZpujMzQZGWy
j3rf/SA9nl+5nB8Av+2pgo5c8jvTdWzupkLMm3klQ4dgbbTxEU4DoYJ/CMbJbykn
gy+yKE0xCdYFORH16YwCkvMZfFKuoZSc4Jw/hLbbVvr6FVntAbuMAvb6q/AGJdvP
BYNzKq/3qs7p3h/NK+eaoIpcfM8TkF8aR4HVlJz1njbSYMxZhK28TFjcojRerFyd
jlrfRzGQI/VP/sfDT1mzZXnsxUtojr9a+3tb+jo87Gk=
`protect END_PROTECTED
