`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CKaBiNIuVSDOr0C0vpVEiFTkCD5B1DcKUIzAp3RjwIEMo4HJV3CHNQQBzLzvRIQf
6jvgjYNHQtp1jSphSnO1KAuqw4uTnx/48CQAtHYwgHwW8gEtwMiyVcDKUuBfzjAv
hqo9Xan9aWaCwepjc/b7OAADhoWL71iBNtkYa9I7SIgOaQIW+3osthJsdVL0KMwR
cm9l5SLIT2ZQxQuLqdQMNlcL3DzhTRnMBivIloQONYs3G9fC1HaR/iKFY+xfqqQy
fsRTJ4KRTIzkgsSRsjlF0U9oH41sVT6gaNWMNm0aGkSUB1YzsytGteJwEJb//jYu
GW3rVMuc85iMXaduZ/JHY8cpPTT4tRQ38JuqGxMk+and7xNCE+LZZt5rxJv/c5rW
k/RdwEMxQt8z9RzyWQzYkq7N9XnvwSGLbrF5HHVKiiPCVWcdV5EuR2VlKKGpbZ++
9rUeVwhyJ2k8sZI1+dtedpLW2219ep/cqX7DNPfSXiim5JtbpGpjKlDGamqMuvVT
6wm1uCfQae1IWl97DCBatjzX+HmBp9c5qutVm3oBndiTUyHOQkpJ9iQ+Vkgvosiu
JEci5WIfw08NDJSMoDeqvC6kpXZRmvdLtS/SeUFIGVKLUYN+5cbZfFdycyWfPvUG
AG8VhSpbkEhDhpicQ3V0A4DTxAmQYaHyvWkC968xFM3CtYlSGYE9JGY9rVlYbZeO
RqPox2A+M4RYXcxPfXlFlrxqMYoICV//sz49U5LSGTih7lrCz4RXlmppzcHoy/zm
mGMFfaPpfURmi9otJ7N0JVwShaY0+V3A7XhWv9lMeT2T9qbRGfesOe1D+xxIDPhV
hemvCHqlzA6Bw8bpfLFmB+7ItdlARPFQWncNShCgalDUR5RYwGSjPT5kLt+qKuvQ
fpaY7yhF//ISXkcOzRdl+0d/3LLmziNGeYXeItyTgFnHdLqX/FqYMGQuZBQgknt/
P82bI9DQDLcRAO9unA7s6gNvZPrTeTojWxAlMtTPntBZRYs/1g6+kTZSZYWXtEvU
tuC2HJjxEH/wIMwSRz7SB6p/GKNX4SThn/dmpZfyDsFdSYs7y8CSRPVT6BxMAIYm
ApRb2nwNgMbqfQ0ESXCt7PbXeX6rIkkh4UoaRWlb4CrQKU531AHqH5LgkAAE95iG
OxOaK1illuftCKh93aS4IGz80dEgQ65XxPFyMsoBeQFdozEtDRiyVXmE9tRsQaVv
Ws4+FhO1ePOh8stOZ4zz4+Lay0jRkcwF4SVVU6ZrC7AVKz0Wy5bSsyHSzPivnpsn
I9sjJc5xJVQ8kI4mCNJgUel9y4AUKtsE1gYWotRkT/a7dxjs3lQjrNoVkQ+r0mIn
JT5yx2Kl3OBH53IoCVsWtD1sUB6/NEnUH/udRjG4hqNEHTInHSL2zefzmKGdcjot
Ptb3CY6RDgDDpPWCy94hMsGuMz7Hkb4k9FOJ0VZ2Bt9sFLIonkm454CdG6uRzXJe
cOBoDrwx/tTb4DM/LANKkNrft+7U1zg4Wgl+6DAQMesW0xsoX4Uebev7m0Tv/1yX
uP360ODYbfbWfVPnQmWeZQBckSFEUT0KIlIF8fh/ZlNlBIsXTPD5NNSOXutvUeQe
CkB5yjizRSviKFgijgI+LplyeVpMZv6VVjXIDXzTwX53EKshZUqhgP6eDjEU4d9N
HLZEyRZ49LaLMQufdt4QyWhBQzJeIc2FrckWE5vXWfoIakIwH5UAooQ4HC7W66Hr
4spdGkNtKPzfAiRUXKcsrnPnX0cCQ8CgEKe4oN9N4H0jy4L2+wB1j/N+NKx5n/bS
tJD3yjYCygtYFgNNUIJ2PLaq//zCYtCVq9qROG2oGnjhs0lnfTgM6ee2T/RRAXBT
5doawWPurFIaSY/52bIZH/9tMkqdkOBUDHxrgbJ/NIVlb8UaChkfmNBKgCMMN+Jw
4E7duG8JvfR9YVAghYvuIkIxpX9PdxItCfYt+6s5wf3kk08h7ePS/pJ22KwGbKA1
pSeDLO662ZlJ0cmRRJc/zvD5cuGbKOdyEC+ry1gLjAaHO9fJYYhVq+OhXHcL+ZUP
IqTqZ0VkyZXx74aggw99UIMv/96BTsXLD5LuI5+N+lYO/yUwzRaLhsNYNYF8ILIi
khDV0cqKhpApL4Y0ew5FlrH/QqHzfQGLPoKjWlGXvmvsNbaZCEN3TzL0Vw/5NRSc
Ab5sG9e+R2aLSDpxMGps1hCWZshhPv5zreoXGdEbu3vTzr+MxlgedcETdvnRKnZA
sOtiesY6Pt034b5GGAytSvN+lHi4opzZ/t0u8jTe1LvIA8NjWb5faTEpnw6Fn5ac
aY5Lmc8B5J5Tx0rTzv2Q5/E1nAp7BpaGXBioIZJwDPTZCnhH2YOtmlvQikb59V1I
67LCzkOwrIkrQhgWBhjeoIxX7EyecXekHu3vZ7m8MSXEXmcUOWTozx49Hh7v+aZT
2ipZJygn02OJsUoJd4BTFd8lyK2lw4AMe7uWDG0xLCHm7B+/r3+hZnfwysAD98SZ
OVK0qowS0RA/Jizk3o08yfk38/3e7sa5ryDNKfywOQgNJcrsJL53shul2i0/2MZI
65qtQKKl8O201hD/2+aXC1H3zY547Op6+eJS1Ixl2NTgmenRLjXuQpOg+PiUjloL
60Lx+0mIjJEhVOCm/AQBnthLGs8uWPGVioe9kXPOVYOiQB42G3E19iGXkR+KxFpJ
D9tQkv3WT7YYavnZ2eSaN9uPfXBS6BAF9PPV3p/e1Eqe9lHjKSJIzc/V1xnzoAFy
gePFjGmJzuEuDS4LJSKXjZLxLgfcq8tw2xk4iUJbC+G0ROWpFvoTBCPv1rKDMcZt
gwMBHmfW+X2RKpMlo0yivU54zTYIfRiPIHau5YiayiJCZgf+uP0x84U7iustRRwl
3pBZU9eqlLHo8SMxxgQuTLdxp2tE+MTg9jiXNIUNog7vE9jqFwfbA022PqD+WNF0
NN0FM3cc9MC/NliiFy+et1bIVZZCBv1xVRct8dUsANUc2tfb+P77bQrfE3KrQwfg
SrWFTV2MBMEYfblSGOG4haTMo7hdkDsx7+skEw/2F18FVWStdXxJsWulLTOWncjp
BC3UWaD7XAVTD8pgTSi12oN4qnmvLr5gQm/jZhuskRDLoL7x2LGF1e9P0t4tmKYb
FYMKqclck1QCe1q5fwsZpANdA9froznK/05HtPAKV9u6WI42O1fjg6fC3sN7fQm/
nO0mXb2MEpMtxcfwsCkhLeOZCN23Wpcojw8I7SmEbzhH8XUhIHlq3rqMqUzDjaks
+4S+TnzbtA3iGY/wocPfMta6Mvc4Hv1P7wNMmuyoYSI=
`protect END_PROTECTED
