`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JQEIWd2FikgXQ37mNft/Perr4/ZV/QNNYJqIdnBd6qJu3FibHTDMSKZDy6/FG8Iu
4V7q7JhKpq3tlUt1Cc/m7N8oTYTktcW+YkxYrx4IBO/A+IDxZAKxBBHXsk21P99U
XHMFvbo/X22ZLmRndnzmPjZChh3L9BBlEboQkY4BWNOx4RJnB8io14jLUFDAvPOI
ixMdRQm5b+BuOXIc9d8ehlrAE5hZicfBn/Y580kAcKkm7wdu/B4sxFABu4jvnUor
LX+9RpXt03VXUwdgMsYp+4mN6HiWQqENU9C412EEzQmDLZ2N5vHh0qgiEXhybdMr
pEyJ+EhCzXQm0l67an1luXUjVAfToEeA+2QrWJ41wWfZOKxeJL6QlZKiWXUHO4xI
WXCdtfXGVnDWtOBIisfGJcOCPMODgE72nbQ6njNeKa873HoHGVvoxa/ioOFFGKpj
bRXv5gxgFVs+CKHP6PrDmR9ojnDGUzDW0DzQrYQ7cDQWyn4unFv7YGcAef8sMJ+2
0RQGFp48ssVxl4NUdr8YbLPMEjwM8WrHeS7z2uxLYSTKHEBo8lZ5covzJaAcQ1Zs
IKX452JXEfcinGw1hhTBDv8pqkVBHiQVKKhGtB5y20VPHkp9LoL6xC01aZ2TfhFN
y5GnHSR85sYemdSe4t6f/xG3bNYCNKP4L9E3Jh2EA4k+QhmnRmXsmXaFXMwqgDd0
BYK2yYyPrWB3K3CVeWTMr7zftF8BaRTI+7ACBGGNEZIMEv2tXxBTHnquJDdt3v5W
iqbHCnbwPhGUDkxbxn63DeB2ksG43HjG8gT4CSkqbkJeK/boinv6af1+OkxJzEyZ
JrSR+881I+AbWcgJ/J8ho9LN1pBLoIOpXeRFbLWa+iE11KYlX53OclZucRZ6N8XR
VnBpU9iilyFCETt4FUvFmle+Vb50UitJTUteTy1M5yH23lF+GBrP0jVc3P+JJfdA
bHkHni60VmS0KvIFDhQKvzHc9oO68m81Uz0bP4CxnYGr17a+dYjbPsTUZoQGKx9p
FlssPSkh8CdepL7CWM+99JqK8OL5yo3oJZyPDjdJt5FvgdBT5p8KzCc6OMY5NKGO
trQKIguADKTqz88KQN/gVvJA0ayTrgI+SRyfyjoR7RbXECuOPgBxdZ5DebECyaD/
qkpXtFA8Iy1N6ODRZyW8QpxO30ssE0gWfaApliX/Ro9VKds3hnomXsfEchAht7c2
nfOcoPIHlRT1/YB6G7+JUFzDtYPRTtE+ZJIjocvhPpUPOge/ZyQ2Q8BpI1PvAXgp
QXPm/D8MQD5/POO74SzqE0XrVf6Tmp33OLCjxjOr4Tl/L+3pFXtgOix0pCNYCPbz
cB5Zil0nIkBgM5bTLBupiPQtJN3WqxMT6gXkCTjy+bOMohY+Q8ZKaaEPCdAdV3KY
5UfGApuwUg4/F/HuqJ8onTrCw0NmYzjEi0FcyQaIECriSAuQx0lFsTP6N94X5VNt
NH02co70BFXTxBhmnAXZDjsLXNO3Dh+qfsZxtB1kcra5U4XzYaNm0+9cI3ZstFIj
hYI+yXj1U+hFXobm7gShzR6jpmyqw20MkwfGRbfTvIGg23SaLZP7Bh2SmmQ/UxMn
AZ+Rvlwk8+peimlTEOB8bXTY+S3MD4w12GPQAdy1gAvqGLAJcrldyUn2kRuSUBYp
Wkgxi06IXekAZxz12ISVINhro0hlR82ZrMuadwspSlDjjn7Lwp5Mnck96EK6+87q
2GUQVna7lPNzUmpN3lKwkGcVJJdSP01IG9yG9kSX/e9/21TgLWnQ9u3WlOv/VC4H
XZXvIM+DKgS9fL2tr0xd07FGmt5iTfofBjfIhdLXPbOuVrGD3u2a81uBrb7/RcLe
6pVW9hBTZ+kWY9/M93J/Fstp9nl+B0h4EcRiSBKQWhS09JlDngrnc5pb9EFP7FyJ
L3c+apkr8bojnKw1Z4dcWufSlqHgICz94VIQ00p3hTMMEu5brLzKb7+0q+UFz/u5
`protect END_PROTECTED
