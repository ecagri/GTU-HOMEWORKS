`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E0lLEYdqLglC0BaMP1xchjgX7/rs373fjAbxrm3l0tboGft8OQ4J3WFMHN3cr2vT
aDJEMkKhdPzRXHYlSMtFHD5gERDgExTNhNEXL7V9+82ZHW9mzRzoCj/L+9CkyZmH
DLutNruwf+2l4tKksi1C1VEdoTysOH4Y/Yc2MXKPCX+D7uhNvY05iv0vRAHpAut8
GCxLeWDjq+ic73ie/zkxESFHnsCHl6BFW+sfvYrNkfAUb54DSdW0aaZ/hLzTJWyh
9uUA2CZrgWWo1Z0Aq3zYekKYbuXZq5WHwrveeVXMTLEUQwbEe8edcOCua+LpEcb4
9iXf4S3JWicTJn+8Sx5LSri0QsRuZTV14iMBdWoA9m1NRtDdoX4wNBi63kiIajPY
k76FuNIMQKFMXv2EPLfHu7JAFozQ6yP1D34d2E9JEhK9C0TXSJupEMEZ3Flki/7F
fjm3KtEUKYKuJh7HFkoNE7KXvDX3GdIMaYEl/qp5MrpbsHbBDipY0ochw/pXtJJn
SKzjhJSbkGOqB2EfRlZOoQ8JSIj7JTGCmBCb4tW6FjVH/DHoAUh9t8P9kxsv8VB9
102BkBlGX+Y1dTctXOxSiEjIMktVshzrfh6P94DrKodAeTi23AjVvLZ7RiWLfWAK
IZ9IULE7BTKQUtqvLHsGZVKIxj3yr0XwzmXqt+O/DvcrKH2q6rknDGN6Vx4L4t43
UswuDzU+EOsPPT6D5eQMC6G8sIaUdVz0whlIC3o3ysplZ4BHT7vV0LmbHdofF74G
wfbnV/OpFxZgHBnEpuBEa7zLBvvZJwMb61FrWHO1rtvSmCyXfbzn7axkhVU2dtyR
gGkQHiG9wGxIjy6pld/SUMhba9FjwA9X2j3n/juR7PCHd7F6MJVYMtsNjqnN6x1H
9BYZCO2GJ5HgJ5kcNov3QiQ7yqoCLt7Pd9+NsyQuJ+aoYDxdv2T7QY/D7YyRJcZh
fqLlfaiXLbHb5w1noywxVU4zBCJeZVBz9bcg1C7+ATT2j3qoUJqhS0JHTAxOgnZL
Up8fJQ4cY8X3hcpFJCNk2Jwjp7i6iuoIcdkdzUf0twqwpKr3KZjz9bdrXZNtAx0c
3kK9fTPXBvZz3+Y9D23rAa0kfG6GCgl9SlTwUFY9kpXBpVtl9ojTKxr2yLrkWkSU
7wVm3zMCGiee+dWetdnJiCAGds1gdPv+vZcPAvNFbbBdcFlh8RNIN1GwQD07w2Gc
cgOtMsrENknMEjHxBBXBb9vvV82PRDmz4FQasMvxi9Ty+RLlDxNnIk4weLtzMFan
Ge0bbIlCryzODQ6kv6/Vj+zvXXjeJL21w+HYc07fBjnqdcvZ08u9gcDUWvKIBNST
yMYNLpeNszHDmJlufgvqcMTo+sHEvPDm9Yz6Z/I/k2D1zO+fW+s8kBusxHZFjVui
NUh8ReKcz11BO/AEaHaO6rIGhAVCJoooN/Bheb1sOpJSxAuYBn9pO7OpUks7vCXh
jhP+2ta7RhxZgogyBH96LREggUACcQrI5stOF1QQ/7JF1o34O6H7co0j8w8sxxDB
hCYAPUgb10S7cpc8ldmQta0eS70WRN72WFDhQD/YMGKM65mqRZL+Vz/VHZ++EJSs
+uqTeSKFlSc8rRLZ8bTiaCMbV6S778bx3yvsQEwoab/KclUWBEupM9aSqIgbCOMq
s6I2O0UWsO1SVge5khApHC7zg93+pTNgKrSUln0NzFbrc9aIVDnBL/uUtdPQOkiv
+dyoRVFvQ9TOynP745Rr6ouR4PHe5MO/iJmImn/6K8CzjWOwSGNuYNH8Gzi1zWGs
RDJ0/01IWNYqCu5eVVTmV9zScEE0qMWkRbsbaJ2WJnYgA6jWbhZBOzK45o+oIfNb
4deKZievj2/4Vqv+MGVeTRb95ZPLzn2/lc3Sw2W1JWg0uf8EdA5TBXBWLVg6zbk+
E7UnBHrih13GfYeL4J+kO07fKz4viMdpADMgJ6+I7tnLpIgQN51ABsA6ooeSeaen
skaGasnV7lSTpliqfuowZho+HzqVJQxOdXw38FKLH5CWuCuULr4j28xvGjSubP92
d8Kjvain1z8hmSSbk4wdreb6nUbCu5cWgwzkRDzQHoVA9jJa9LuDTD5StAXXhmcG
IU+w45Gh0f00+NMbIGxCh2rlFwDbm7tNh89JcBbqRa3snsU1qA9UIhWdwPEJ2zft
0DW1fkOt4WZ7Ieuv4DuiMgLGePWkeZg6AcsMBYcHWJvIpHQf1DUVyxANcr0ALTzz
s6QGLqdSfwn+uPpd7/LYNGddnb1j0+8TNgE4Bm0dhHKwVpDwtUOCchrSo7Gx859+
QiDxu9YRYEdNtjrFdl2T4BYAXXaDBjshum7cMsdgNAxNmIhNc4SgmFalGmBcQiWC
Vi9ImyTDwJhHModyP3syhuXWwnIfmsyLc/oJ5kmWfsBm1HEUK5mZWXfeXoFV6uit
mLl6id5ABXuqINMincpnX/XYT8xhZx37r4oal+4laN1GFCEJYxdsB34Oq8474ukS
kv1sNtXYfS9Ae4rep/RbKCck/ka6dygQZk2sc7tGlRcqPNE6XltZRSfUlP1pnN9p
tN+1KcylN6HQgi2Nord777ad9nvDlylu94CmPFu0urxxI/sw1t3hjzXye0k16cJP
eN6xJ+G+1uS/2BBouccWIurn/wlLkW6Wm4CaZW74OlASnThK8EK1JsPFhBAB2FdG
ATESTRhjzOhCLGSKiFeiE77OStK1QidGWC96u5r9PLjcpqR/pXLE/o+oI6ApeR9w
QwDDSBMqH4UChPwJPwepkvRNFZ007ad3+ye43v4jnTZpnHrVWfvB1ofIZs628Eca
4jK37ULu5LG7K+Cw94PCf3+6kfiurrJNXQFRHofImc7CcW/t5jtVH+kfPK6YonMy
pmI2gvUix/cQmnHitOusl5pVbbzRLBD6XLP5EAcJj4/AvUCCQFQjgORdt3mYNp7Q
QllkBDYVmHzXKv4poqeiSy6j/u6Kx1Juc2xiunMtX8YNva4Q/N+6P6kqsv6c/l2M
o7InjTPHvE6bdz2dXzFs1wWOn2Cr57nAEK44nCbRTDDt4BUhWU0GEvCUoTe6/OhX
oy6Cr+WKeoUSyDEhH98ODGRq4b4Y6UieBt6/JedbjrGKbC/6vs1I7KeiQD3+NIWt
FXYdFoGvL8VhZKPM6OKOHavjAF+kD9jqISDdHhPGsJm877UYF5FbAM/d5hsbCBuq
UAsYsffhNrYWLo7quE2nFGQBHQ016w+HBnSE6ixjacLQBCOnrOEyv7e3A12XTGo5
KGFELGMAItu9P6b+yIzyz9gwfLWdMsdgxrGZ9s81gLiU2JP0E2EXwpRCELVjWryU
zgCbP9I/Xy/IIBaa6Sdx0wXXFY2RMBI2CkejlyLbXAzOG3c+4hjV8THdtuRW034w
O7phNKNVcQbhgF6TKQ/icfHz1tw9MRgbbpZ/xLlG/TqI/Z6bpxmJTvf1zL6wRAqB
Wi1NjYzkGM6hHGqaN6fxLBKHW0ZNOTMNTNcq3qYpdd4U+0cTeIkLONNCij5CQv8t
aOUNEEitKXTUzW5ll+Qnd9TqduMN5JSx+J3pn8AXHWsqL2j0IMs2oOjcUT7tEIJi
wubrEfhl9KIfnHv93S1yYdRP4CPHYmUMEqCntHape+BoLPqCKBEUOvYLnvry3Qfs
2+dHr0gj477TAeh6NwaQPmJd194wR8k+JELghQExXyEDpmCGw1x0wMPPWWsRfF89
+PNYbMIBgwEGdQYlNAmU47rDhT0+cyfrsevdqf7qQPf9hbBFd4oRqy1DAYZALt2g
RAbUbbCi50S4EexmHcW5UF9lkPJAQEUfSSzeNPUZYwEQXhU3HhB3DxCnyIzPda2f
DncPeiq/GT8Jyuc20yAYsVVGIABBACcrYbX8HWtzSRAfgGOT47uOFZsoNFVpcurW
xvTJjTnAwSm4AaMhnzobAU8SXBStFxL1EhumV4Z92YIckWBh7sywUvfJtJ0dFs9b
FOwSKFHOGSw7liRidkkupL9sJ0h+uTu/CfMpiTB9B6c+riA0LrIUOHv6vyognNcR
Q3hZla/r7zKchJD/347ryFj1yNuRzBJRdgxhG6NW39rGSMqx+kqxNPIqwWxC/5/Z
3BZId+5LOjYPxrYAtTkJsyXYIkcv+rkBC4ccDPlTVR1uRGh6KtVDnIbtsk12GLhn
U/ENr+z5zlQajEuMN7Rpr28rFwXl6kiYHTr4sZq2wb1RgsZllDFkTeap7ScV82x7
P7bBIhIHY73TA4OUUfOHsr4uAj8Dt+GC44PC1lWurTQr8hrND7rPiQkyHRRU+t+d
xbiDY5P1CXpsfNTeFk08BIA6nr97k94vaPjPLA+E3WDxcOr/93yJvuzKKqvgUUuC
p2Te8x2gghMlUjX9bZ7w8fFQk9oIRj4rnOd/5+z2zqD0K43Aon6nmv954fUzCjpt
Oh1qUKJ7RcmstyP+W1VPzqDRMLzLJLAOQWRNkWnqnNWW9PeBSRzUVvoBj9orRJVO
ar+ovp7bU5PAIvLmi88TYFvS43qHYH938UKj9641DRks0hA1MfUecAD1NTkJJFwz
li7G/74M/y5TOfvmlf1LH7i/pk9pgQ+54C/SALHjj4SrKEBJLf3DYdL4ywJ9AOvT
z8wnhHqbhfxtIku57VUmKOYMkg0n/dX9Ue4T8NsCPVJfCkBFBd+ML6hV9rxvDcZf
VQYjJqKPN0OVLwi39qhsaQzxJvOIbPQf69+eOxEX9djuxPwG+NQ4zc+clEpBZ3rd
xw3wWR2J16lgF05V6deqc702K7NMW5/wLx99BEvRdQj+m7TmntER4IoOccQVUiPl
zbhBETJgFeohtpTEzwghrf62ByQDACGo+j/SsoYalF0Ki3eVEefbEUH+aGU27een
GVYOOY4RSGt+aKtHgjkhEyMEvAtkpb6CMQ0sFV/giUiJGCAV74KxTqBHDltocD4G
34yaFlermLWqGq+A6fXPqVecKtjXr2X3KCEe4icLYfLT5easmz3BWco+oQ3w074e
LFTwaCBGEdkEdSb51Mxqzfc7TE3mDC9NV5G5WTSf4pd/vRH16jLOjJUQuxaT7FpC
eYnOkOtUL87o5VzCibx6GtPixfj0WkklmwX7Cwb14FcptbT29zoSDD6pMOa4Icej
SeDDwi1PtgGOtsneelGg24K2RkZLa91qE00qsXwfFx9iC3/Hq+77XSRGQp8yxTB7
1wx8OCSHJ77amytF07W/fu5/VAXVrwa+g5hcyNNOXt0susyPD5t6dF2tTGWAeEat
llsabY3nIoGKgL7F847k+RLgHeJlRCiCwz+w9CsXyHs1A70cPKjXZ/iY5XMrD4gN
FvseHcJX5I1Ovjak8gFEInNunk2YaUJR9k6Ef5W39GqBgUC/Tq5iHQ7pyhq6rE9o
ePHtv+Zd8UAG/s5ZWHfoLSB2ehOK2h3+MOwxdkveXAXwowoBL3QdI/BjNGR3u+6w
nrZNTAC1Gdhb9sW+v+qTHOROWkle0pWcblUtZZxANUW20KyGdX4ZDx8IIomN7P4Y
8zknd5MDGSaSDJPMjKT9+LyQLBi1+LF5z3cxaok2Jpjf80gFyc/TuzKZVUThI8fD
UjGoxc75BtPWVK0fLYPhhWz9oS/ZO33/CIKLUfb/KHo5fzwZRy9aiJqEe5OKHtyx
f+2d5FE009YG7hMZ3WsCeIJgukZwlNoJ6Pc6zU17LbyqDL1YTobCBeE6T2de4T4R
d5SSK5Tv40ReFnODO+MsDKokvn3bB1xEr3xUBCQMcSh6LwrZvRw8CtXZ6SqLkM8F
Ozns4C6cuRL/Ri5LwL14mxV1vpc5thQRfoqngciVFAsmm4f8mNXzgl8T/0VE7Vcv
pWvNeV2E7jqPjPF3fX2nCeCV3mW2O0ZZH4HHt3WBeXUVqClsvgrXTfaNoxxZtuJ2
qGuZalfjBj0osZeb2QAt5T9Gkl63YPqcpr3/ak7ZdPx2aDbOCwFoahfe0ayLB43L
kg2+xVCWtZ50BNwQx5p/5xRJ2y9Zqtg+sXZW5RXqodB3jyYvzHfjv3mACvp06QNu
2vDflNM7m0GpVWS4gYlV61ghoNy86/kh+LdI2jXt9Z0NqSE97S3I4KjwklJ1taiQ
kM0CfhFa5CRFgCpMM/1eQaAAG3gbLmDwwK3nrVVwE1m5DkZac8LBx78W6SIPFc48
Dh1tR3SeZOPpo4BWUNiWKjmJ8TJm37oGf9m7rB332WBOI4muxyXoKNPjrnTA/A7e
kGIPHG+Rk6ugvyRdkywi9skYlvzYyCjKjzuO92iqlUw=
`protect END_PROTECTED
