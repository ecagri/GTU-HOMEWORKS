`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uKF9t/D7scNBPy0cJSFw1b09xSRJYnGwBTgguXAGwCfwKQOpcrWDxqsWkyYC17ZK
NjZDVZajcVpmqjUiE5k0NuV8vujXwmpCfsxKGSTaX/epi3d2KCZestCgMLn80jdl
TbAgy19nf4qVdBTrCFAflnN/vPgItRT3WO1SQZ8jc2fy4XbArI6aGIcVF0AjjK+v
2IeYia2N+G2DmahmJN5g4yU7t3CVyh7+V1/Oa36yrxOY8xGEf5SH4cNDV9yOxzcH
VwJcenKfjFk52ibqv8MT2zDbL10r/DQ8RJrIeqS9RVz0P/yt7KQzAzd6JXA8IwTY
UfbknbZJiRi9wdLl2vsbXjVv0k/j3JQXTHQSwfxEd1jYyHBalOw/NznjsRDcjUbw
EVxW0GNXo6WMcr9hrqDVgNRgkf9/z6zgjC05Zujk87D7EL5ekMQFR5wm5K8bqGVa
E73TmE9xpWGq70T1+qs2ugbrKEi1/F6eTkVzfaJZTtx6/IL1gPl38NNfq73J9Jpa
BQ5KA+KVD5yI3xYW6+MvbBEonIrKJAfnVWmMq8KoexG2H2zSI1sdfcDhbcEeQ9ep
reFKCcBGg07nHfnoGwpsCesFAtGtSQEJUjY7gr1ptIwaA+tv5jrSjOrp+1vW+ivi
ijlu5OPPCfSqS6kb653yyezl00MWaCh6O55sZk+dsHSPaOrlCi75LAmXq48GhQ4G
UUdCXVBqNq5pu9WvQGm/J3YLfFajeAT4mPn9ZDqF5vZylLR8K+ZOOyBcCHDK40qF
mFCGUje5yWCdPbDoVT/UWi75L/g3PTnEZWBbkMMsOcVPxdIX3m3Ys9JtchaBkeFi
dJ+7Mbsr++GIEYlDyzy7PKrIOvpQl5T5xmCm0GikPrUFWBWyeSaRPI8BPF18mz0C
i+MqgUAQujd9N9qzv28ZRbTVDxIts23Q1SP9psW2LNihAkZGsFvWHgEp4FCaZG38
`protect END_PROTECTED
