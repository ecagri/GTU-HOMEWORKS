`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
78COyPZQC+xqLRTuaTEyl9QvKFI9rK612oq/VCT8StM8zhu/ygGgTnAEUO8UTQNp
DRD2qgMno4wXmskaBQqvuhkG8GQgbd7v0X/xpy3lUcVPgjQOz4k/oNyM7cISSq53
oM960JjJvqB6Sere4ymf0PHN94dWKR/WzHf8DeyeEW5X9MkGSqxCdVH+EqtvaJIw
etqQCDbSj/EzYqKN5dWDkw77K/vX8D0+BLJ827x8kc4J9PnM99TnA2uWvBrhNzkS
Voi1DSygk8E4rA8Iz6eRtHjRdR5dKyhN5Nppr5PpKdOp2DSPi45IHx82n2sci9SD
1j7cuW+/Iui0I+a+65zp/tk+1tDkoLF2pSziwmk0PdOGZzP3ueyx/JN70o3MEkSZ
baoTHCfNRFvhcJv5rYyzO5oKuAIRfvYrq7gAmRlKWqYIciI17sjYSYwv2px297Cm
PdXHsu4oRJOSoaLPI4LpltFOXj5j90CagfE7rBV46XyeHEnE8qI1Ype6P4zft9x4
4qI2V85ZzTawZ54OOL7D61BXHjxECT41bkM3BCpvMJUtibS9pHSqt6DVHlko5C6g
Md8fnhOFn2su3IaNOfJjz8/2QTRKjWcBLL6f0kplHFpiRiyavawORF4aDlejmcn4
EPe5hphrg5yQX9DR4W/J9AlT/N2Sgpyg+JLud8xD989o4xV2V6FYtaB5a0qqeU05
V03BgVYc7mgM63YUQP4VzxYatAw6iRSsMvdiuXb3Wmv3iBaHffgkqkDeJDIEEHcA
DCj3h6gMXdu+AER4hDUJ1y6NCMifh8AUjHbqEkpcGMjOtvUAJE3qvkTbmlAP21H5
Fby4h39NAtHi6JywUYDCZexll4qD1dZ9pQ5cXVVeg6bwxlWbfSfrV4nHQAaL0jEG
wPvJKuFRPeD6xvpko43qhXuEDtbsqoj9LgiZxOFaPGddNHTi7MU0yFMGNkzIAGhF
iG3KlwbbrfPYgDTT5wa1xdpM4CjpQgLPGhSS+ZhWp/kzekx6L9iXrguDRoRaR0Vt
`protect END_PROTECTED
