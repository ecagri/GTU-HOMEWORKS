`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eQqrHNVk3dkx7p+61XbH+/IlKfDQ2ALVcFV4q/1RtttXNTCYCBo7AnPFsJQesgCj
MJ0+1GviHpF8YquZMPtbBhBGKOVhMV6yOmjOXXEEilQwRqq6t/ovNTl/6Rhp2dQ3
vmtX8Yagk+63uJf4Jm66F8S7RGxR4oQ8Ya4oyrJtHy9IOl1nlspNbLePBCUnhU1R
UJn4KvZ3upJUCq6Icz+eeGb29JON7jTu1E/hOSPkGBeRoQIvBAWtLSFWbtTHIMDA
CSkkjI9V+bUaLcv8cpq7uxntd0HDzk6oP76CVGv+JiCvFwxUMSx2HlX/pk5ICwvq
Y3WKnjulYe2jK+YeKeQvZjqUvBv3OniIeCftOd1LZjhPBlheAJ2fLMthQfseYN8q
r2jPGx55St8mvGhV56jKXf/3op74hl/z0EJKv9x1qYcecpUuMmzv+HEFOG8ytil9
RTer0smSpKQsI8i3sUa6X3SVxK/mg7M0fM7CmYJXRv1jgHaNeSYZ/Oy7XSv0biLs
PNsOInz7pRZXVL6q8c1/ZOP6opWyW9HBas2vodVQrHbyP2961fd0ETt67tNv7A/M
FITZwsCOKqi1r4fFCHYNnJJnwd6pBsIw48BJjKGUr4o0DZz0eT0eSZA8w7+aItZG
shF+2IY252Tv3+mNV9Syg2bJaIGbZyJWUGLuy+C7HpyhldT8OPfyTKnCpBRdRCKH
VRHNBWXm+I1keFdz2/o/mVeu1L1AsiKMd3EztyMe493dzBay2Y8H54N6NT0CBdQu
lXQgY8B1LN7sDBsOnGwLAQXsavGj1K2MVmhrgnS9btljEZ4GDunr6JvpmjfALz1o
jTtj5C9GbX++mqRelK5JwQqH+VMkQ5yJ4RpU5HqYmCfSr21YMatV0jWG9Oyh3DSG
YE4ENFuPDDbQzigl3jk73R2UDUh4lQCnFLKta/kSEr7Sq56W8okcP8XLwC/1DOgJ
ogxuf7Xxs+tXfySRi9HEqLsZqQl1di5m93Vnwi7Z8kKCO/CEsXJztekRFIao9GWG
pY+9kSqOApzKtaWpzP+VtH4/wu6WAq5BGEFs2KJAea/cL/6APAFIF9X689V/LccZ
iV6LkaBc+A8Ub9lZusEzQn2DaP/wzGufzrGbhcc7XcL0vmiaRAEki+/nJS884Vaw
+YON6Xf9teyA7jtqzPUabo1CJQa4MniRqYz4aCZVFZrQrlLsdsfTJfVGdHzz3txF
LP6QaTzEuCP6AuUpjxAyyXUXtXH2BSlFiAeFQTbIFVMLsA3S8n/BmcPOBWIYwYdG
WtMxGB00gPO0IfggAOMnkXo7FVh2RnpwClgzYhqUuMSxNveS7X06ovPepXMtTNIU
ETLFP/MW1p84F4sYhouIY7mtp5nan6iMGVIa/0WoCsObmI7oiWmRw7BQmFufbaS+
Z05KU1b7kCOG0nit3NNMwoyPYEJ+JUp3pk6oKORqGhNSITDikRILxxyA9g/g4keV
EneMZDd7RRx3mmbOFK8BURClN0ui3VRorEgQZ1t2MnPR8Gok4+cuY0gy+E32f8RT
NADYUNxZQKTfYKCsDk98x9N6mqidbgNKnvk92VzJuhXKablqMYFTcX/hQmJf/tQQ
WbRgOE7dgE/YlRgRQS4FO5gz7cG9QeHvYh8NIFDcvYk7dECS8cvsL+5Zrc1VPRt0
/OZtgpZrhsbfs38/cTJG1ZP9BBA5dh0DO1hBwLpHPVw4S2W+Pm+iV4B9ZzF6c8pY
RxTn2LlL1UMaaBXXGWc1w/C7Sju/u2CS0EKDhPKP9uFsXaDiR69cpPJvYpD9hAuX
/L93icAikin7ozWTKekk7I0EODVIsk4ugcjAmwKTRa1DuVGZ50PnlS2FoNn06MA8
FNBLCMv6cy2REDKHLfla4Uw0foChyh7UlyRkhxz8xgitXc1tRoHIPSLzpn3Cyef9
vNymSrgAPS+MpbYTFxVHXQotdxYoCpzE6ur8wwRqXfwDuJOluE/ArgiLLIW21P/V
gyD5fgpML3v1EauZQ3fTWSctMBGllyIuxOd2gRCNgJ9sToqqu4+6V5ROr5RUMbmh
wj9uE0Y5c3NFjvA52xU10xFYJyIfI5RfOZvvTG7uRd0b+kRAKn9Pk5ks/13lu/qk
cvrMQ/yKSuhdJ/WNpPESZ70FpqZco4nrqmtCXzTwmXH4xbA4k/sti5iWShUdRQUa
hQLsdqJp9hiyfP/BwVyMEK1Miq7n5I3Hh/tbp2VJ7UPX8o8cVD93IJyZko3U9Al3
skwXjmU4EFpPF+G06coiZ0i/PN9/l1olpgDbr46MewrPnqZYAtRZBtw9aO6PzCa3
wIqnyEGRkuxm3ZZaJewkmDBC/Lt3rzYOGfBeRVIIvzeNFwE0ciFxMFEWOAnT5zXJ
YF9INKu7elZCUHLgiFSeJtqH4oI2s0lssreRBerBTvy6ON0h48lyRbRQpLrmRqba
e7n3JN1FryM/+uDLlJNyQMaENCmhwre/GTqCLpAT1wmOO4viAYhA78uP1WzlXpgX
u1kGfp1fTsZ1d6Z29Nd1IKg9BpnbuJ3iqXhbGn3Q3E1nNIgRqH0RI9muf5eJFPpG
oDEw/K5OdhYcqnVG7l25thHLloylKlyKRz2CcXLkFbq5XDD/b8WgjfSZgifGZYbA
I0DtHRTKEAHum1w1uHufT7OJgE9yQRNGWu9oAehMeKqAAGjttCKi+IdE6+pZIpbG
ZdB/yq6fRb5ELlDRoWVjdjZ12jlJKs+TM3ai8DKd+BznlTxgrwqUJplEyrX61E7M
gkC0xRhKoto3mpnsHOH0iuIw28WyTSXe1x3oNBJ1WkFU93vUc11+ZcsRHMMWenga
Ik1AcmlVW325yFicfqMOX0kp+En0fbK/sl8LZgNOMtmZQc5v14l6YL/Y4W3eiewi
gmsQ+ZxHzxETMLJRMmWlbjEm6H57SI20X2NGcdqIJrTK1MyFu8i1/sfW9J0J45I+
RxrZ5IHhuIjcEHMNbcGCAQF3br0D/fDsz+4tRo/+Va/ykHPSBfwSl4YDFC0etJLy
CYY1Qeb+PtDQ9saTQ39e02o0rogUHTS6PFrFTixjfDytpwLJo11DCVf6YyVKeQ3B
8aM91CjKvHbpuxgSy9BZ5oqKP8tT2B1P6RT60uyg11PXbEyh3kOj2+s9yNTLJLcX
vI1M2top812upCpnxcia8205Ra7OACdiuXTCned0ybCtIIFvBz2Kt38C7473opLi
3VyR8U+MZx9AAsNHeoKASHBg0fR8yI3HiVmlmg9BCJY4UVOir0H5Ji9IPz7ijWjc
sSqkwFCPRP0d3SzrD3hlQJYC4lICMWNbK2YNOamtZfwE5awv9Q3NQlkf5kQZXf8u
EUVUn+BxSP/rw6M09E2OPWOIT6VlHapio8vDNjJrlIGtAKXDhNx6WMCviWqggqyl
MAXlODC4Sv8lDjaNy5vAHzHyr8qSKpoCkZfc4JYfVzHGZDLHAaETqL0q6RqP8EZh
EPsx9Soa0qqlARoz4AvD/OFPUyytrC1pec7dpEcDGvP+h2Uxx8zYUj2SA9AjEG2M
vkYz1Tev9dXBgIn07sAShxFJDBqHKov00g1uYMVa7n51SdQBp74gY8h6Le2TwsGe
er2HSMbRpflqx0rPNDxcATdAAVUOhikbrBbozpVA+Biww5YxeM2hDs5RV1xPHLlG
XuEEfdEKQW38k1xp2rv41mpGLwwHu92APjyARCtK5WqLJ93c1gMkdHcI3/9rA0Sz
Whb9gnvWpgzzJTZEP48wlgscfv5/FZFlbxso5RcUaiEAQEczANAHe4u5na2AFbyB
PY+J/BTqhpGS/DQnXHl8f8XKR+B2ZV3gX0+L/l0v2CteU7MJzuJ4vwG6jvvyaArm
27GNkvr0VxWTvbtmgq3sBK8LIwbnSYAFKC7E6l1mOiEPB7hqVJczA/BFEuQSMe1J
Sf0WR6L71+pqtfG4GrxXiz0ax4AMLro+vanNqPOD16kUCpFo2lXCs6swbKR7XKun
1/Gf3aUBGB8ZWAPvQ0nJbE/pBa1nBnFH8GK7NaK6qaUVozp5RobRnTEzZtwVDTCT
M2LNMTZ44VXzqq6Vcc5+IYsSH7J3tnfDP7LzhQJ/adn5pWsQigRWXHeT3qTT6cZZ
gcLGr+xWhjctVYdp6vZCOOFKMauSiZTlJja3K8Y/3kE7iw8drevUHOwqZGYbxaJg
F98Hr4z4C3LuJn1dXCPlJHrY6rc8gFtDUfVGp/7ArUCadAHvxWAn5NF3j0GeKlE/
54ynBASk4bEn5QDwoJnHFpkk3P86GSDy/GHey/Z568RLaWmzK3Ph2dmdaV6Z+n6y
mRei5driRpntr/rinyXydQMhA2AFEyDyAAtjMgIGfu5Q82OG3QtVYa5AVF9hOKwp
8cMY5SgxK4XWAgR6c5bFj1FgHtqZI41GuBNz30CvBoDkXKWkkLpVxV7WL/FzGhaq
wbSxX0ANxcn0Xslna7NsrhBYF++NXm+kyc0wcPQNHuM/iqtwjx/MDxhkZyG5HTSf
`protect END_PROTECTED
