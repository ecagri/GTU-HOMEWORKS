`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ny+pjWMlTy6dKYaLBhi3vnC1HF/zZep8IRBxA37CJ21VcgBkbXyo1Dqr26nNAJQd
OEjb04KRYFZ5B5AY5fxVficv30TLTn32Fm4zEUPrIT8oM2UCfIcu1x/ww1VvdqrA
89+4ipe+xMadzrpd+vtEGBK6eaRSyX/Irckv5xb5+epudM9MT9owdvKVJvLhSw8s
jggHY/NeIgRyECGDmhgr2wr0iB8P0zIfbaXVxJO1ESgTN0vOwIzY9QvAy5RxRJTS
yl7133lOV9z6sop2QC/Bsaa6kqWPS0+a6m2pgCKvYp7XVKMyShyafCLooE2Qt47v
Q73/LHijkp6d7+CTinsx0oY8n44b/LYKLE51WDv4ak+DHiE5OferkMoCQOC8f2+h
hnKS2i1MEOJQlK6r0NP8QDyTwaw4Xpix02zPVOHm1/53TKjdf3ZqQieeCSlti1MD
/9hiijXp/fDno4hT+3qGeQ==
`protect END_PROTECTED
