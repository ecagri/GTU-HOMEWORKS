`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
limgEVWDoMnzPVaSNPOrL+sO9dTsXUPGIA9wbDkz6/cW5I8+gI3RUQgCdolsoUbM
GygGhviveMtVm/gCuArAqSJSwZGGjTeuOCcr74jCpEEuXXkHlcmgM/ijIpALd0oz
F6FWkVCcn5zzcdQjp8FAMoxFRmmZvd4Rft4DNt+8ijeAyOPo+nhufuW5cjYdxAjS
7bTrv+hyTRPGcjPBufqlZLf8XRoNE3iOhtX4AsbRL0iD68hrWcgrjnaWUg6YcOsV
fPZe2SbK3pfAjmNGWYZnRIim1mKiAD1bEsqlJPpyBFWTaFZv8KkL9RjbRPUJCGjg
8CWcqkysP/XC0aVKRRjzj54hF+tyHMe8cyGCN4KTzsIMeBQlGhDYUBCUZjndfO7U
XCKmWaydv90lUeBzjWi1E8hnsl8MVg0uypaLh2WvS2+CtkiA1wYzzQGlsAT1tdiB
9cKJNpRQxj500oa7AmSlbEl5mTgAfB6boRJVlc2vAkKJVEKVK84m2IXNtkUoxRai
KZL2AdoBGSHtraCz0dRTD05fauRnTED3WEmt17rqF1M=
`protect END_PROTECTED
