`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i8enDOUB6C33gfJwT4BMozv4+vXlb3M/w1CSRvMbL0LxRVa60TXA2gK8viYdsyoR
funjcFbZka2RvAw4Kj+4QqZv6e0DcqWoW7OleTNl3+hgTBYPRh5ag2wx9qv8YYtJ
pIa6l5EeZlaZ3FZFshPm6viKy66RZpmpjpndUh5uxE2T0OTjH0AIl2wWeTiALzPv
nT059OtN52+qpKmh+Es/ur71g/trLtefDRhmtBi+0aZXht3DjqHiuJFQDnjqQXFB
QzcX1mOXZhyA60ZpFolx00Op4ksvpsb52Tw/U7T/rUedouaNAnnoiEA1vc7lZLqT
UZMf+R0P8S52GzVVs9M38VBczym0wQ71Aj4zYh6lw68NeE7WwQD4WwuZZfho1r4l
pW8xzrSVbQf1Ss8aHlbiFEIWqpM/ZGmDN10GT3KW/t2jkqkRCtvnpmAVLfuNoTbK
pbo1TLIWAQB+jgF2LWxXbuqPKAXZCsfLp0s01DqArCxxSclIR8rPtB9omp5JY+GR
qgxM9YeIHoH+dNs4c+UViOF3oYGlnuMJMKweJAWW0mkjBdPYxwwa7DK9rGQF3h6f
BnXrL4UNhcC+a60enoT7HkcqeADatpSKe65XY9ENcd/D4CkQWSPoDywug8UU4E7Q
a8CLUXb/0JKDOFEFLrEkUGKMPl53nGr+hzDOawPlnrOxd4qPimMX8P5CDno58U/n
/nm2AuO91uV8S7Jtilmgb9bvSo91IXf9VfBTgT04zANJ8TPP1gwh880w2i+vZEPl
4qoNVnSrtqlFYcYwUkfWQ32/Ejr+cGOu0aMr5ZI0aVvlpZwXat1ENU5WA13uZyRW
MYUATeogUIBcHHy0Vlg+19R34AQ9Th93QOxZli7lD9cvjI+oUdSNmY9Q2zkP3sYq
4ZBcUpvMpm2N9VJr6nFd8GLTnhQ8v7pzXKHq6wWi5Q4fiM0h0y9lfsgQhBJ7zCID
eoTUPkJ9QcXhMY+NKmSj0pzC7EAVtzR149pdN19yo1uPgHUUGsLnNA7LCpnhXF6W
wdflcmu+fl/wULqSxDg2Tiq1tqp5lx4y/lMjYuXVjmSJwJn6tTx2V0qhT2rbe5i8
NLlQuNF/RSehu1DxM++PtcMpld0Gwl3P8it1HgRAnGIs0GCSW0EdSF6pRXhDIk0D
YbEOaVQDKQxWHtPlQa1ZBEesCBYFgfMd3t9vIBm9KwBR2uTegUKfe+ossyvS/pgr
+zRXf19xCwDE86JAU46uEn3RQ7CLWWYNESA/by+JhzG9fhTq+0NJwOm4QjEsMp4A
ct8SiftxWmm1L75mNsJwarLll4EBB2tTCJJbII/s4hrphS1e3K9Ff/IflGgTsDbu
5rO2SjaSO1+IzMqiyKgTPHSADAcg5GJ+PKQ2fFz6RBAljcA5JuDe4IReBO+/jlWM
KOoPPeNu8SgurA3LGpER9xuSu05LpEzCacWt6vUzglIwa1VuRaG6MeUo+cYJOoZX
kAYYa6IbImnGJWef2vwYjkXNlV7hex29TH06HT0jF8CHJllG+BQoLCD3Dgchd89/
Chxm4U7qs97u7QOYZRfLq1NjCiqGPlIIo0Vf64i4yfrKCr+qUXzKknzXv5JdPXeL
SWatbAinIuc1XaBbsXriOV5wm2rx7oTFlu5rOxsrULdOJ3XVhiATVlaQlh70uSlI
2zzZOaANf0/+J51V3AXEsOWa18XnYwoxjZICNvOhDbadFJwBnPzscBaQS5rqjngD
KZZGYJlO8+bcax208V8KQ5gGgHsb4YizuxDvfAg7xwffh2nhgFudn/mA92jbYE8m
LGS4cIY/n4+lxFs29W+T21S2g1Hy2xkBO1fT4HICOcJ+Hp7qxgCNoWVumNpQsJLg
7EurxF3pv0aJbFunUbVq+TbaAg6ewTF3Q+DSvo7z48XBhr6TJNC12q7qadrm5WmR
iWlKE/LjcYVGiv7iybynWXF2MN7/ohWCz4MIVAw/o/n2t7F9kpCIoKuE6KMsoOCG
976JkYMd3vnz0g0PvFShW4xZ0KX/IlEiDknDtzmz3saKd0w1G4b7aeagohwZb3kV
4MkeDKHwq6Thv36uHNW9sZpPdeFV8FFMaBp8Bm9y/hyn9MXI1g5CFkp9fGSDUv1u
4310VuiHPFUQVC0Nl2btAAZQtCdch+AbxLx5yFaQCXlfFBFvfN/Fsm7GZ2KA3m/0
WYopA36tG+57OMLS8txfh5M9XYGmChro20GHA1Wkco7U9o1RtJVKZecRVXSW7ODu
Ut0bajPdge+0v3uCv4kzajVagtWjtcyu+cT2Dk5is0+ad0YwEuep9/XEg/7dOB/G
HjVXo2mLq1SJSwfsMl/ZWhs7xTpxwqrDeR4OgWkVYke5tmJYLO9C8/NnH5bloVRF
kXErNcstQJkHF5WTHTcnT7RRSkOxDM/Ip59imP5ZK3QqEKAQ/p7Og48VnUQ4dZx0
OVh1yX38jWKVIjbMpIwuoQx1/ux8C8wwgpde3CeQ507yJxygXHxSA2MHTI2Ujp/4
4PssIh+rWTwrvFRfvmp1FxCdIjUM4xYhw8SFX7jeIEt+wMyxlafl3rpfIVfoaNak
MiRcUlfVOxyScbanFd0gmpLn6dGrmDhQmumCX/ztl3ac0sDoo8SJXh2yX2RAWE7r
htBss8THPWHT7xST3o9qBBOMn8eBZPORMu/E6FmIBwsh6toqGp0cMkPlEUWnvmzD
UJyX8BmRRe4EdtRT0CLuMnaLXQTDZxYHIThWvE2U4eHhyZ1KVLPuu6h9PXy5YtFy
ztdKJA5/PUd10Vsl90NVgJ8RlG7pvN6Aob+cim1jKJQgw7mGWfXzxTpqeTJ/iqfP
ubBWsMCXRtydPF2UE1xrVtEgN0kEEhdRAlq+Qa5clEVcFUIRkj8psWXUknpfTG/C
DiWopPtSrQiBH4E+P54FA8CG42gx8j11HFyR6kqKRnQVQuPAjQFeCKUNTJXAn/L2
6Z7BIRQTQYUCKBVp1KEVSDqK5PObcjj39Yr4+ZUCVzsV7FnngFS2oLylBF4Ldvql
W89naDcp3hyO5JQBCr2BfVjRaPHi61I36ri/k4PCigxIeWB74vcjfF7WtUFd1mkp
q6eYJ8paE2b0wLVyXYGKxpVBG01Qy5azFz3m86wGKnfeK+P7MdDjae+FQZAfkbP4
a+Y5A/xh1AKOLwPRWNVtx/DKK/8cOijKdKkF92WAuK6cXafRInruq8uYyFSPubc2
GujPR0AtvIi0GrqHI1cMaok/RNHJK+cXTOnGPCg9mR8rAHYraeoyBhkJ+Gzj7BWR
nDqmVFoegdQkCFMr5+vzMOLUkdRz23zABW5dozjbiqptuDJyfPCLEwz/me+CHVKa
oztkFWFomuISMRKJYOe4qHtyp2t+9N9C42Y7CrxHYshlcrpRHAzjaGv2AtPJMgEd
HQYM1tpIB0QuEnQhVHbJ1G/jkCnKyjS5v2cGJkRaVrbnTVDXW1sjbcXD+B7ni8bB
o8tgE79rZOi+cfqw3wxBXjW68ApcbhpqLdLySdW7KftRS7M7K2OHMAkzHbdvBsSx
8Wecuf1DCTWgrkbmmz7dmLt4bOTO1RcuNXJFOk1dVqgH9IHajH20CIxXzOS7y/Zp
z3RY09IBjd4M+WGF2NPcccKK1b+PkHmNX3si0hUY/dZWSbXBCjiMEdNnCWt9oq62
/5MqhbjIImYlYjWf/GIT2wQRlHudNkmygYrBldqFndSDfCKqlXNChqsIYf7SsDzB
aApq/KF6D11LcpImG6RRqCHxEeSZZ9ev9gpukopzp07OzStE25NSJhM7gYAHXPU+
T6ytmJd1AHyPw1prB8Cu5UrhTkZWDb2IhaBnqtYsTK50P1cE/URl5bEKWAVWOa7m
SdMrXwJIi7vQb0Thrv4yxjmaj4aCcomP4BaRrytyg2192UbDsgl25toEI0ZXqXSI
QJzizu800pZcVP6hzQUPaUFbRhwMBY6whZItgIz8niwCgsjOecN3Nsh5hxfxJOYl
JMtSnEYoot0q9qTPluv1wUMDlp+4je73NseG7/8wDIuN6uZbVfBc8JEDFzypG8od
YQOwq/xDAWA8X7v2UItioTHGHaAQIFDadEjTOwEDLWwUfPTFl9t4zU8rGRZ9xjOb
HueeksYnzmCKF1wiRs5sBci3K++rduPHJBGoEo20jMzDQFMvidt9En3UQHvU3WIC
MsReUCfm9sChHep0Tfna85OPTotmmpP70W6faUhqq8lLDkuq3QbKQy3F+0RC9LZq
54ww3ABoqsgo8vSIG30L4c2UGpc0Fj3iWYLItqWJipPd33uPnLLsb1s3ReEf+NPZ
UN0FMOaSVflvF65/eWU7IVldpO3fx91YacquXeoW0BSFwjLaEAFBj9aBZqAxIpHo
Qh1sr3/0Zgf5b6r1Lh86dt0uh2cTkJrSNT+NqPErXXKylfHth1DHNGXOuGmnqdzo
GtiHf2dr1u7/JOzGVyNeT9/lvyKd73wallO7BNnObctp0cg6V58DNkJ+e1GR/xS2
ZLCJ6HrDVW9hYk8DYu0XJoeX9YwD9RTIPwcjoXjCQBHg2fF8fqnQduFFP0now3+Z
P/jF8j2fk/76Wcq1ZZVOaOjuVJgGa2zcMc0pMUXI65+9lxFu80jnrf4F/xSgZDnI
iaSq74ID/iW/SyEk+P//U2cU9mhVhvU45Y1K4RvAAai9spivRdNSWGuLCg+DCoEM
HWyHtFLJSPfdeACKvH2CSwoVHT8aZSzUqcZV5+j3nmwqhaqaTCPwFbcEO4V7uZc7
pHEltD2VIPHgiIV7Prr1pU/wt149+LXcPLbCTPzALf6jlCu6HudktzIlQp/N0PxZ
HwMUG6/bDsd37jmkxPV36oGLxeDJRl6SepDtdzN1k++k4s3G3ABl2milDHZXio1w
fDz+zvr3kM8xjc/E9uUhpYJvNVoZOrx8PvMzd6aZMl147CQLpCGORarJ8tmEAnBi
002vf1oJaIIatU5ey2TWToc0JLV7St8LLHXkeqsJlhPab933pOqtDa3gfII1iMQ1
`protect END_PROTECTED
