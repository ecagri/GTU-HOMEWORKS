`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+zpq8K3FV8Sn7ExQ29hWVQarJXa6amHgWxaAcynzC/OZ1+XgD/mHrLHBWMHch/8m
qTE+tF/+jIUjMA3iDxOkHNc/aLZvcAYqdYSMdI/nhj7voF0k4jxOWwi0Udr/XRJ2
ONdIkKdt8Tvx3/b03oxPbiXxeaNzL0axuOpBtJG3pzN0rLxNJ5enMPalElrhXUZU
HL7pDAREvxzdjrOh8lHdFNkZVHCA8OSPHcCT5+Bj6jNWiiaci43G+uMmHliFGMO6
pNDLv7r9278q9eNJjerf1942rXn8WIN+47jSnMP40k4hZ0RpBZWpjRk4O2Hr/qgT
vYOiON9mLDJH+Xvucwif82rklJBdcGJJ8yy/wwshDrgWgpwKA+abxwLtfyBrM0Oh
NuXDLv/PML2teTp7sEGxa86jyS3ORNxYYcjUSvpOJftYEYZpr5jPgPf0i03C6bJu
p6XIsit3DxTO8W86BjNAJcAtHjxsHNDMrPQ8TP82J9J+vmaJz4Sb+990iubkZfor
uxSyVWYDAsgJjnH0GLIIG1o3AhIMK+RQo/44tmXtRGnvIet5lkvtlIWYoap881F3
rclrNV7qupaCLUkF0fIYAYcJvMU0q4IvqlKRr9s7xzfgjh9gQwHEWmRv6jwsTF10
o8B7snrkqP9g4w60U3gcvx3qIFKEeZZkvGGvNHlCe994gKS7Zr7fI6UUILM2h6jb
JJz4MlqgZ90HziYhIFqlv7Yo8frXpy71eay8KhfRB5KzbOq712CPNTAHjSDYDP2l
gIaQTg7Z8W0g1+ghrfwgRe2ScfMH8D4Y5ccUuCCeuzc7ADJUewe5Bai2u0IiaSGB
KaEV7WiJW/8IDIR6A8FlUA==
`protect END_PROTECTED
