`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HhGI9Bb0fC3yJa1kCCSCQJb/GyMkz2Q69VmVqE52iS7D6x4JTPeZTwxQKinH5tiQ
VziHqa+GdIUQ8cyWZ30yE6f3kTt6IlDXtajLmVUsyylTGYmaFafrVQMs9ad8XIiP
hMDxIcCQ668djHOCnEh5rBMglvrzDdhnDYKt2TpUfRjv1n0SisfDc3e9HZa5VyC0
XvhkFVF0yJoMgYdJgVv6R9xuyhtzXj/Urdiyy8zOArCg3a256icjOwcvkiYXbcfN
UM9uYrWxy8CZN0Cb9p4sG1BFjK5wNkzDWWzrJJOmB4UQVD7Df/fYAEvQv6EY35KR
j/0Qsvskh4DmZJqheXDNZBrypCfJau3uED8eg5Jx2h09u9ZAHX4z2vvn/tquNOSM
wXwB8Jgmc8oKrGElRTX1AJoeZr1uT5aegjwylKif5ybzn7839tAMEvEpsNolG5WI
0YijEVweLLu/kicGSTJxkDAiPKubV+KEuNiPixJ1Ij21dkh6YS4lAytXTg8YLIg7
K0C/VbuAi+udOkpWGGuw6tRPwrPiKtzHSnidPCckIQvQbf/c4QlDKqiX3fnD3jqV
ATicArG1smeairZfl/vz79nJqcI+AcQko1BzgU2uPH/qd3GC+fhcdb6iu3M2QsjF
s1o67j2Kk68RCaD8kHciQ0CNdKpleQUkljZm+Z2tHsl04RVNcgSTTUHTQWs34Lgh
s1nWqbtsKxz7UJSat+Vb+RgIUEjLecjsHdqiZCjIQFchL6/9CkfR8PPN0fUAppWn
FsYt8PcO9U6ZieEIOJvzxJuGZAjNE2Lephf7YgJvWKWc96WaAHuL4hQWhtNkkVPn
7cfnGGflImOmEgYq7Tj0IxDII1vbDfgvicKUO3r4kiIJsc1ac70pVEyEoXhd+pnL
LPdJsqj0qsCnim2PE7RTDXpwzrBOkFtY7GIiKVy9YNEkDj2XA21ujeq/APY4nibF
/IZWM57bHhrj2dk0XzD7VTvO7aNN6uZSIU4tgsmdLU5lQrJSgWS1P6DhG9GgmLqk
guOz9rnvIIxNkkdTiNdV1axxY0yof/2I6zQJt8hW6JPUWvXnGLOraK3/F1rqhilz
D2E1XpkvtMA16bGBkPc7TST3OJMbGvPSQ6PhxTHc8Xdcvt/vOeGD244rxOWbkOfR
fcJd501I88hfTppwPmcXGd7+NoyYgdPYgj+fv8kyH48tyg05gjEJfu6/64m2Qo/R
yB9evCkHlNOccrLJ8ASUYoGMwUW03yKfjVnStrXu0m0FX1+sSaIT+jcf+SiMrvDH
X7Uqim4y/dvhaq+gZUEJqdJfml8swpsFEkDsqy01cd6VRFYRivwdMUfScR1N3wJW
R90BPVF9GEG2TbEo0cj4Kezla+lhMiYVyNWqlbsEh4VB4G14MZs9b/pfJqoIda5c
P0QEA305x2ceOi3Td6YaKjdNfC2cLuM79MaBA3PU6x1rwvq3iLKcct/3j+45QtUe
k2NMqX4yBo11/6Nt1PYpEbJ2c7Pqekqr+QUfVHWMAup/a6U/4kyQOafVEX1YRsAD
yIsv6nFpRN9PX66jmBPpNRtYtN6LzJ6YWuW4LxP+f2Q3gFHAHJs1hwW0te0vQdhD
zpStzWL1pBt6lqabwVz6wHXatJ414z4XRuqWVnMw8J3fcZkRYj+nLZe7PYyBF21s
1eu7Kwwo2an/PiP3S4zEkC0ao9z0m5Mq2hN0nazMcHMNeUQpIxEFBdGr0NoJ5reH
eqqEamoWxFeQ4bv25CtK/jc7/MolFKD8GfpwdIS5jX84gR/vSDKiWHK4K3EiKGED
c3gg06mokXYiiLtombywod9+SAXnvZukBohRau908lNPt9w18NP5yw+ecUayqFw2
ltFL7Hx9BkzrFPZZgHMd7DM5dVeXbVq0J7B0Ns4yRevXIIf3rm7aFVQDUL+OBMMz
r90pm8Tv32xRqZ/3O2T0dUKuEo9nWHcubcNWr/dPUyWCvXc6GXjyVahoh1O98Ujt
CP4/68Fc/uv30Cv/17yjY+z564bHJmseiNjw8FdASOiC5CyMLPKZ2qc9hkh5KmpE
fQS/RkiT2TpKM9K41c+WS9/vkEQw3hQQqdFAf7KuSI+FlDFHrAOnmIsp5Fpd8upK
S6/uAapqVbuvupBS7vNTnxTVGbWza8XTQIwaU+mGdWhjwvfAKI0cn1mjnC07k50G
4n/XCcqmUonnjLkm7CHA7wTC0W5eoYCCEU0UIpgOkUOGTAHWkvleVEDSj+LCy3Vd
eCANSzJWfdLLS27ohlqXBz/Uocf2cNrcTn9kjxR+ZkPiUBVyizW0piC5T+1nncyn
UQAWwNKJvEFH54P4ppZ+svyzGY8Ii5b7CTgHF54DjghP5TFCB0AilF+X7KhRdtgq
6Zl3th8VKbAwS+9ib2Ua+AifkrpYfI1tnri+B0gLsRuZhvYHW6W3Ueq7QBxeJjNG
tS8Gyn4saJHWeHKeykLy0/9NdDJNryoGZ4I9Z/sYq44VfgRu+5rtQimbkIURjAjE
ef8igxJEbwCFM9VFPcFrqICmoO5VrN5zXEPpLUpXYVdAgzdHqau237xdEeBzvFlF
7axlcQAt+ax3zwQcZJHs3Lgr24ltlVPXX2hDMY62EYv79k5954jN4fKPvLqx5Ntw
kDCuGyfTZnkMnLeN/+RNE2gaeJDxRt0REm1FByOjp3q0DPAGQONgqOEXWhkJKXt5
vZ8/SW2sAcchVsS2prxEr3teJjNwK+rChoLmRjuT3c5xJ6mQC+oRfhvmzcEi0N4+
PclyHyzTtDjp+Xx9rgYlHHXccQ8HLNKOwS9mdDXRSj0Z1ikHbNE/ttjiErzvc8Rs
fYIdrZxy5XYLWsesvOUe2IEocYfKCfKBEjcj7YTl9MQ44v264zlia2/3bxh2wwL3
Eym1JZCeYxQNKlpHrtbGWZSu9417tFU1fZtqZRocp6/HOwnkxR5mK2lCTHcgCs6M
isUjyoMS0CLceQc+rIBxrF7BuqhGZE5D/yt/5Y5Gv5884vER6SaIorCGcfto0yNN
Ockh0hO8Bu7mHhk/uDy28Zjo0qNudcfhzRseqEPOGN7cEYvLIrB2LeaE8XntOQ39
gWmWwRCSPoPUdZJnCIchhokTksWmUflfaT7gkf4T4qzUWAC1Gw24bCt9Ehv9Nhmt
Ef6lBovzoNaDbfsAZR65RkZ4xKhLDPYQbs2EQhvqhcZqvImhMXpJK0bTQLL1JCZE
7WNLMmyzDJaVOEa9mja52iTeXkBYwcknFPR1ZdWzC34DGz3KK8JKzS4cSX0bmuWY
9EpczvegL/KkZTuI/VPEZ1rK5CZosa9qgE5TbdrHaueXAYd+nT+E1emnPOW8Kv5n
K/c9SJC5wAVR1HwnQLCmIsJCqBvhQ373LHkA6J4scgmza5nD669YB2eJamjW/xF5
EGfTMV/UlryqbtN3coB1a7a8ONf6HCypWe7xpgKii2TX7Ut4qMQpal7RUypW1Dgs
MZ6G7aU8tk8+itSq3YLrweqv3pwJ3yjY36/u2Uy2N2D8tclrtn+RMBY9vXPJ6PZv
3XszGhZV1fbIDHCTw0WuafJUGN/2R2vI31wpc9TKHyJd7FdUoNZ56ryKcSmg3XnX
JwB0q5wDFrwowRR7mR0imoA7o9uruW/3MNT32cxZbfFSAojGapPtE6AoGmQSln7M
A9P+tG6iCStb2S+YZ80MEs328aXz0RXJ+s3aNrQxF/W8Ce0tSZ6snoQhk+Q0VKEh
KgkKQpWVyiWX6OnVg6FqZnKWWJ7VSavJCNJXfhLgOBL5vbJN5nsTXWPivB4kbSb0
run9dki4i3t8iJ6TVh9AIEwNhTbbBds/e5BBO35/bvCJsF5Ufdg7FZYEo15y+mRe
jG7MShEPcJxuacx00V43MQ7aCFePDCYdcwZAZYyNV4vAf/0hFnVulQswfVArGy2g
FkfWEViEovE7hhXu5ow5SbYr1hr/LVYbyk+vKFa3VR6nvl9GFYgebPNKOafKbyYk
Hjhg1bDqWrcD/PHdITWUzGxzpGiWFDaGyAeaKduDM/oNCUnfeBSMZ+W5FpWyKFqU
j6k/NufatBYqTS+53D9Pt0S8gPQZ1O8E5ZciMEETySGUPTS9aSUf+fpfcBnxhEeW
F6zaF9UX5Iu+bYBaJbcnjp3lLwaZJKHkYYSkzTWHP+NQMJZD0TjsYH0C69YHPGrL
c27vZuZCyhpYmUDOmZXxEFbbTjaUltA3Xg+u0P4SbJrkm5QOM4PVWmjPjMO84XUc
rPycV3e89zvaQu7X/0dAfUrfDzs2p8UPIcwvFMxCF9AgTebD/fAJSZQNYtIZwSJG
ptAbqvr1Q8hgb650VSNZzT946vacu27i+fxijwUwRJkd/d1H2OF5JjGQNDscC2sC
jA8vpZhy09/z98Ekd8kXS/+qPSvCuzvI7GoufikLhEUGgmtSRnBV/hbuzcPHm2pX
huXdgcD66DKwlwNZ5UiR6IsxrwWCbvnInIGkNX7uR20pPLZoR/plNJtHmhGa/qAi
qsxrOiIsF2DQaCrWXQtik4JL52U8swXHSPV9LC65XBauySPcvSt9dkfXPaMXXrqV
A5ArQU8jizzb+MVJWr49dF9HuAfkVKcGZ7bOLzcb++4ohp8pjt3WSZYyDETsxwwf
rGpyYgd7a8vfS8t0sczO5uFTJx9UTXptcI/v6AOb/LHBhHsFqe7ywRW9txZHB0/1
UzoD3X7sSpsK04dEgi4JJe9Bgml+9o78znIjG+3+7Kh2R+arhafaFsQ5rXTODM7+
1nwaOfNsuAPeKC+IPPIN7JTpa75fZ9CA60Ubr5WJAL/8YCDgaibt9KdkP5v0bHbf
ZUey1CM0DK9ma0NInft5RjAyv/QnTfV2PTwFFdibR03OIAFyI+ytApBIP4muwb/X
kyZfUZ4tcXmwavPvTcAD8ebzW4h1W6wdBp6RN5H3SSapUSeZdJQvkN+FhQYbemS+
fOD4ZRnmduLej29dBQ9dlBE0nQRaAmbAM37Db/VZqAevFPPbVWRbtaI7Z4kO1F+J
VBlmhOijvmkrXeXd26YLwAnqQCHPl8q10pi46Ike43azn662sBDhHPpYHHy6U66S
IZsPn+sp5d5mWMbqnNocok1joURLpqy4EOwnYJfZmqf+ptZrb8wzvHOKCELnLlGa
XxeoDxcmNnE6Q7c1wglRK/5sxWgiNKuGK60ueSJMCwFKdrx5mkLc6VGYfJe1voV7
Jhq02Xkbfuc78UjQm2uod4uj/e2ToBVUFuW2cJnhTL/nU6d1X0NXvhPJ38M/zvwf
ZRvFV42ULOnWWsekYdITYaNe0c74WqJ4b7QeMdFv2iH4XfVR6R8d0oHlx+wpNQNE
ZckSAr8lQqLmcOxTD0ZYEBRRWxVGcj0uC1l7H2HMxxRarJWqDLJ+Z9z7xptIHMQO
huaBkQ7tg0pW3gmbtelixY5ctxX8ubU2CJGpH4NwhWON6r7+G5SCgLQT+rWO6h5g
vN/5MTOor41UoDlQtD1fE3N3lrNQEMgj9qgtlfCdmKQpXn8a8kYYlioHEtFTczew
lrEuKLfPP+TPY8bT/KHmvbSGcICY9U7SGexJorwI0mT4XXCt93dLOMwR0cLg3ky6
UT9FBhK6BeRXv+STuGG5xDLGSQxzrQHfFjNub35CcBDPx4Rqwo88lZAY3c6QwCq2
Vjh9Cn8tzcEXU9JRyipH1yeXNJKVC+ZuCLdLNrorbjJ4t1VndJtl/I9kgfZKvxa5
oKLPdWhKgCvJGoc8Xdh86OwoCq0Q29zK6smCFbhCmFXe33PRn9x1uvyVLpojJnou
weDPe39/c2QVuoDduD68hcyqbZUCuwSKZ3Z6mUHmnVOTfcdgqxl66FBvDEJOX6Cu
IwJFg1pQkNGlprYaJ7mfgG/s4xllqfIWR2hWfzmafGPr3YR+Njcqsn8GsD+KLPma
TW8wgjaP0DlZPKtbmTdobbStdjaxsv3C3+tMMgxIeDGGi3ed5cxfQcm/V84OjzF4
p6AKAzliNOF8n8lE53H5nMgr5qlccx74lPluQoMZvsTUR/LmZz1U9Vf5bw3YnajQ
7YWH1RptAFI/+/E5f4JB6hchQg1pqTgQ2F3K70EVB5/hGJ352u9ChFRoeOv1+FLF
NQBbWVQb7QfDiHgbcMcPCLdL8sOVRebt6Ie+oqrpEVl/f+UyEkxbE0/ryqTca4Up
uLFMeJJHe5Z6UVr45x6C2SLZG0Amlq/1Rdp3p1rpOZ/7NeHtNrSQvDbtNKP69T7p
Zy9SGH5p5pavoc2DvpohLISdNl0qyJ/eE8OwTMlOwWpHnoOnk6e0kUgFCwZ1vaAu
wiiHrKYCqpRXzTe3qHQn9+DtKZa9+kcXMXKCDL2vvhnvGKhDz7hi+wZhIChEqcGF
2zRHHIJbtmdcDsmFMGacq5CX3U9kiNkSOUFEzg7ivyC3A2rCUstjggNKf7+WIZzo
4kFJbmDCB8aJZPi8vqnoJFmKkwkiRYOyNZTUTL7Tn8AuMvfg49AqZBKMARdaQ3Wg
Oj7183KmcQ6XDpqsr9sKjl5MLhDUk9WE8KLCVN50UsPnVbrKPcXKlBF4gM1nwg8v
U9kROEZ2SQewqovUhWVH+m0w9zXkbf0qmfw2+QV6rxby0jW5V4ie2+qNzKfvBzy8
80M/Jv0QzslIwTAIjVMvjFw1YgEmoUd7Eqmo29Y99XYuxDnjeU7AeR/NRWO9e5fa
sEmiN9d/prThGkFmY8oaQIP3yn/PkGZpY8aX1WPecinCb1JLuqmeztIHYSdMJFW0
CjMvj/X+xYBC9w19k4oygbdRhdrGkdvL9vnTW5auChdrk+R4caDChrxe4oMNmUGO
GcwBpEHVG0Npdb8EnofdGcJZB8Iw/xfAyK3PjmQ8iIBF9jqHlsNON2ZmwYBzyCTi
os4IzTENsykKqpkYP2g1trmQe3L2saoQzkBf/duIEkPoiVVliq3TEvk7Z9Z9k89/
CiXoXv/dFOW59PNc1paHEQ/BuHMYrO1J+x/xfLiph4L1vkRHfJ/t2ROnameI3DDN
3wEOWiwfDw8s03Twht8U7NgyJuQ4KC8lYLJoA2SWGfcLRwGe5bZAmkiNk4CLl6jr
tllt7A3/aHI8RcZFfeCCJsEWQSSSHrzf68CwDYzZtpNv6T89vmxdfkAxUnM9Ew4A
cavB/XWl9DzyhwAQGo4D1AI3Wk0qnbgpgUBnZsA56tG1lJvoG2T8oAWpY3AlPMnG
/9K6Uhf09fP1cBR7VS+ix6bzApHhOOrQpWRZFBke3HICwzrm45FP1yd/HWsd0Zhr
hNaHvaAaAXy1kJJIsHs44GRulkjFBD2FVhzQQvSAHmXNgg560cUlAuqMy1Lp7L1h
cIu2G2Bzywt2iQTNB2T28LDbSBVpzmLfppJGkno9hu34aUMiHUolh+ZVo1clUD67
baJNYDXUhJroE2b6imTqdwMvsgwjqiZht27VcKQvm1lzqW3a0KoxyhIkJ/OqfYCr
YFDW/8a/j9HNZEerHxJQdEknNliqV8W6BHung3Q/fhR2nCMcftfbXNO3i9n6MyEy
KAK6bqSCsy0gN1dkU9K3oDXz+RkC8GytZzE4bUnx9eWiBV+FR3XKkQj+gmEZBM5C
T3rJayIX8SJ6lLdvB39VBdK9KLij8ARP4RXjtygGrf0RbqPz/e/scv1UAQAxsyL5
G98ieStTA2AGgBZGLu+x3Yn+TpSJ8HEAgLciu2UzkW3fc41OPOF9X31Ktv0XUq1f
Qhm5TKWrmyvJQk0CdMDsYlyGUB5iV7K2y5PFiAgMgMZ2Xb3BejPcEa0ioOQjwaAy
IIrrRi5FDxJmv8frThwdjIRM5+b8vW+Zi1qXCynnehtEiQNtvMerDMcnrKlkn4+v
/iREQZAPfY2lKMEEKicfH/ZJlFTAl8naW6upf9l8yG048a01HepCG5WmNisZv3Ln
YFvuOHrSc3bO8Mcp5yRSlVZpKxEl+35Cu9wUhoSurDoT2+hzzcynlVAnpIrskoYU
qRpA2x2BKxNi+pXI7tpkucg6eEoKI9rv5ji1t6HXgJMKUu66VXnVoJA/rq+lmL9X
r6Ue7NPo5d0+5a2HD9bvkravyvptdf3O3UgmJYNDR1zFnN4grlMq5QPZddubd80k
VlIL+N5oWoLgPcViJJRytqmeJvJz/KEGEGl9pK9CJga6Ev1gCm5SIahCagDpwzVl
6x1oI951vTYXdLsVUKOU31C3d/lyvecVU8Zc6EWZCMvk5UPOIvcM2y250cedwSsc
x0fHbzJuJeGR5LBV5bEzkl5C8XgVBxeDV/XELdpWjHAnoEvOxxgfhoT59FsGRGva
vFqTbjjF3JcP+zv5HSpRJLGFl+g0oL3iTm+9EGlzF2QKaPBN3ddHMW60dFfewINJ
YJYmHlvVXaYAmEz/Lo2qO7WLZiriz5Sd3X0ZsUFqr5lGkXIxlgcg/N7r4L8remnV
SN7EIDnCIg4qEMvmfEc+/4HAYTUcBZ8dpbNuDTVLVLdmNGnn9G/zflZRuB5SAqYo
nPhJ6TtCghHVEOA0OpJvF7GEatUvlB/pbJWbzrcsML0+v1pbZK45mO/70VAmPmRF
WrOfgyXTT4C/9NY+tisGT+cncFebM7zx4VVQ5DFMHupEpFuDELH8LzU8UntDzrX+
FsNs9hvqjXnZwrHdGhxqa1Pfewt873+dgG6uZZONrxkYXdZg60SWY6Yd0woDkcPs
0DelOHHjwonNuBd52kpZH5KVbUUFHnSsbRrkPzRmPVw/CA2qPUFBqcSwMce4ouPC
qzUI8SqA1Gpdae/BsIGS2th3n+7IAl1GBURNs7m3uMkyq5QbrbF5mSWwt3Hysu9k
h/YUHOBOslgcxnqO0gYXQ0Lx4bkuPvLBdB97omn8vfInNGiTcKDmoS6iamLYz/rg
ZUXz/mn3V0PcKkiSmo3dR2A5ifWqqZW1sH3FDXgDAD8p5AcsuwIpVe9BwRLZmWpr
akTNom0JVwpcpmoGjyPeOs4fJ5Vp+cYePHS/Kx8a+JdIt3Hs+oIlYNxgcIB6VbYa
fAshV3lmtPr0mzwhM1jTkfIePPu0jSoKhuw2LiyTXdXaZ87Vf/D+m9jD08hKwTOv
MBSlNvlHt4XG4UzpOXNe/B58s8ay+iDCSfAwVPH3+8GdsKpc5ftnF5vC8ENsHX4C
dKKnwohDWtV/F6oC0clbZwW9jvl8gpLWgr641US8DqjiI8SsFSZwdroXg/oLY4uR
S5AcpTfrMN2Rvxsv7tMocgn0IYTouhC1C0M8dzO69h+w/zweUlxOI2rwUFNuHGKJ
5TNnklFlwfebCbsPNr3IkJvpJT9ZD/zememWaDRSOw9mOEfj3oyMotyv+Oh/mTCM
m+d75CGaqSy4FtRFZOFl8RgMVKa5QaDwTtiIRHSnuowT08dYNycNJgcUIVSv8F8V
i8ZfogxrRGPH36FkoTa0uaYXJTBC+7UhCeOu6JdTh2MMsmWf9Y2Oibeuso2tspKU
xGzcSamiuno0drolUL5BBqxG+QRzUA74+3vH4zjHMHNYDoAdyryX31svPtXyq0XV
YMM2G9O9aW1/MOfZAbsEqM2cIrP0qpECoa5TLqvuKgl8iOb5b4aJiV+zx0Yw8Sh/
yMBFgutrdgYDQAM+5WsH/izV/6pD4b6WOjFUcOyjEzyWzaIpNsKpmACM/3N4MRHQ
KwxCHvb1urWr12hThE2GvPoK8jYOyrPCT26R+oRmEXEhLi4hCYaLV/lHxKWtzWr8
8aD7uTLmEaiMScWo9EJjxU/kLnsZvmN2Zkxzdd2gLZ8WDnaYm4TSWIw5vgk+tCSK
Nk0Wxhl7p5yvN6hg9YF1U9SEGK4hV07LJKli1GBcQSF9eQ3YnPg1WX0bZwJsGNDq
HuQQLDxRgogc0pXOC3+gPQV4qgBN/E/e8WgbaMBUYgW3GjXDLjL69ptVS+wLaXoB
oCU282aRIaaCX/EmZtFYBM16qqMoT6ymOb9rF7hpuLkN3MbxYknAVQF4/PMMWvjZ
gIS4V6wciZIDuWrFrM6f7Jdr6C0UAPrnb1aK0atGx/fwnTK4n3ogQC9RrGQM2fqc
tkBhzGH8DjzZhzQV4/6HVjEqgRs6tveFEqJUvmg+wL9I6TWfTDk3uD6psaiHY137
g6Cjo5pRO7k+blJYgNP0bvXXvHdSib6FKjw+5bnE8e1tSSSumqygF+nGM+6XFQ3X
H4NGJwNqIpa59NlHRIJYZmbkzr/4pU7OeaoB+cDdWq1kS+AArmRpK3OFEHcMA7Tp
uU11nTu+cMOJRnigQu9YPF308gbcvvqxgQXrDvdwuU2R1cTkRH1YwBRhHAGbVGpL
ZBSrP3SwylYmrTWlpPQ0KOrScDJd1XXMy1KwrS7QTbbaU6z2qw0bZmBX1GD7fY44
XvlXUmeneBrMzfnAj2R08hwuJi/hOookPCRVTcihK26VegqLgH0IP1pahhXv4Jau
Setx3RpPkTTj2pgD99aPPIY9QXxKQLF7LpnAnHxE92BQ2G3A5WavMBqwtiRAhtRp
6DlXEj2g/z37etpgr6cpKDeRd+6qHCorBaiwx54xUNj+vD/hXJuVehEvXeJmTsJX
eMJfNg4zj/rUHseg/S5HjPanRTPUZvvsJG8uvNQHyg+F9ccfswVgdLKkffIOnK3y
O4JiinXqBhN5M/xGDecfiGCOMF89D/yrQ4qiFMcPOUA2WUSWhtyFSLM6beDCTqxv
2yv/RrTOoZcjzEPGX9LZ80TI42WUcoV+Riywp/TYUflmSC9cduFijsTmh0zK0wjE
JyMAEWELn/B8K+hCUhRZuAu+0Zy5mQvJSKZiMiG68IGQYHu7DwHlIxfcCcBm/p4w
qcFJivql243J2hTRwpGab/OruTRSzPyqwVj1xg58sx4CjnFJfS1KlkPanRy5k4fE
D6vrcKe+NbzjPehQq2APdNQGxKAm2+t299d1tWw1A34blTbxl6BGJWgo/nWMPAUk
JRJJCQ/Pv86PvSfR9OlLDNHxPtMV3Uz1bgNwWFYu57IQPeKhI8AVtF+YxbQ59kIT
uezPTuEEAGMWpotjVaiABkOw1Vq6h7TzR3/pIvvjS1dfT5xgjyVr1yPRd8gjqcjU
JZPxET4ESU9vDnObgGHSsmg+qN7YxNYFtjlVFEG1yR6Bfuv3ao8tRrsylXu48xQY
eqz4/iGSd1UNJznR+JDahOvIrw+yRZfyuFClkeuk4CepD/4dIcluX50Nza9qlRb/
7bI/bHpX2MaUQlX+oMe8mqeUQNf2B4OZsnKTgL8j2tRhCsihrfLR0CiJk9cDQ9W8
UQRczqY0CeENBdZMrZr0Ii9otyHzVEdNkrw53U6OayZ6AJ2BR90DgQf7ANnJKMge
wPZA2jm67w09HhHxD+s1YQ1mn0B1cNYPbGx44t1MS9BwwdyJvv9ixG0oMeKqJ3W2
g/WUSddxO3hL2aJbCQN8NOva/jGaVeYKYw/2iTFqEmQ/D+X67UMvaAYiSEVqBmgh
PSfKp43FXZeLZbC3eOt5vMLl10I1sdMIj4p+sA9eJw7d2lbVCKHLwp7q1NYSy+/2
2pMsgTP8FZOa1N9AIiVpZvuf9dgYYjwKQtK1gDHgc1/9VKxKUiYeWJKLBmQgZ0Ow
jOsQYqfTMmbw9IGCPTLj19lKowtlrcpyJRymFS+2fkShfqymBbYmQP2S98B7HnwT
s+P3uh+CZj7vlKdMLXks2zTW5Jeh18O87ONuHHd23Rlc6tBJRoyxMcW57FrbvCvh
fR/f546zM5XSPTjbJg4Q/tq7S3AQ4JHQi0njBmbs7RQhfDe4N8Jb3dZP35wv9Tbs
XPxAtFyMzTZwpUymtZtVDvYJYh24ejWhmAF2gEKWbspAVx5r8h6xI9yXUDueWPPj
Y1pEWh/0ZdKEBcnSf17JdXTNfgMR9AEKx/Tx6jkwxaUdhYqq+46NOyY1X1IQ8R2U
i5b0Zra2NWiBw1DWY95LXrkMpFkVL/Qw1mOQFGOiV8KcWgqC4FgiJX3jzy3C/0e8
f7U8iu1IcUhyBUKWG3bD3II6cLl9OkDJi16617gjEYBcdSWL4nlwZhPpbtqG3tto
KqDBxM4jV+vOM6J5COn0gi4rbiuH0y1ZbBUYYIcXgIz8yZS01YWQFMgzUDUb4+hx
SAT0sIaMXMgeRNszmqEnd4JrhBGasTJPWNKDC1OiHI5qJ5HY9tz4b20VK4un/rHR
syTjhhu2itF2T2ylZmheAoJOT5FpAJlClFO60Umrc0LUMsxg8qSXgnN/w9yfPTFE
3O1HvERTh6Tn4G/05u/raYXcuYlTdTDylCC8syhbo8F5Id/Hgv/9/aMfDbxhUbJX
HH7gVGL0rV4C06PwkgGekqq9Ld/utSfs2/qfk20i7qkNlg8oZ5YS6zfMjbS5w6mH
3SKemUwFgnfmkU+vs+57oSBhrf3j8DsyWIReQup6O2lnVryDg8eBCfWRfz20YHp2
UBEE/FPUBEuMUzdJA0nyhlA0B6i2R7E2asyyksXd5K3oyKvpmLfZdB+JfyZl9m/6
elw5hcNnUSoRRRohHIC0jIINsSsXSvcCPSISXydtE3XQC2zVEjj1wXkI3vNUA1EW
w9K3wGm64XSx9t1ay2gM4FGvirfCeb6Ek5Gdnmr1zssDHZXT42rNgPi+n89t91WS
ytGMn61PBvIO6JASnMeyG1HGDDxdAgvVaAAdCJzMDpi1+3JS1llF9qjGIsbR/mru
yXZGXznG1yo5P2tCbWR1E3ue0eYRzBkRSB+Os3qgaVFMkaX7P+nG7s/1Au3bBu/S
k9ISalw++jC3V/FZGxICHXwkk79aYRKOnZ3ThSAGnE7u1aM9IYzyxR+/Q24xvpvZ
iD1dVYwCk6OtlNALuBvGPUWLjTECt+/Fvu5lYfBhpm79YJKjZZaTajMDuR0oJQxD
+3pkeQHEngj8ay4fnTgN1DcvZHQcJ9j8wVtygFR2+QLGguSaOIIvObDHJL8JuMsK
rZ8seLaP4ZFXMn9DgF5TGjceIleGp+/XUOQByNTK3eUdbPM6aGT5G1PHRf4/hiuz
vGDwUfjzFDgOP9SYwFKDItoJgNTZga8PYpiPpRW347AnBH6+6GRASOPiJBi+UMth
4WnLTa1NFbaRV4G5wNguHfXYbitb/GAHBpmeYAru6KORTy9PPQzNOggxCFMqVbQl
Vm+gs5nPSKem96To4edtEEYAy5Ufg50Gmo9cYitMyXOTQBl+F+8B48p7WQrZDj3I
m9EVIrE12ANhLWjyQjtd7G+BkSi+dTrwOaK2n5DjgyMhXqG6Hd2+JxLOcJnpJHuu
ncR7YFScRRymKzs6J2jEdwstJ7zEP2WRcdfDpay2aj9LV3b38sGCWkxIB91Kwyo0
H+ugidq0iuOn+/8NJ57VlqfVwwg+y2KJtpf+D7LaEjeiNwoQlFYy6MAYg8Og3/Ak
wWBbxJXuAOkE5TOQBZut8vez/tihyF7nr+9T4euI6XiCFRyuIGOF7QTsVx0JMvxE
ceM01G82x8Qlnc5BBsltivlO54NVlXJ7e+5OxqzcXkYptRpQlDNDdjvFFCpt5UsZ
PBLCuaOQxMiMvVSPOHOroN/3TL1SNmq67hEZYUSopbMBF1EvkO4fC1JxECFkXvYb
Z6ZhnPSQZTmSxlsQXKi1T7zRzOvvEdup/3ARQAzq0hRoW6FTqUGYTCG+cgFnwsRS
KV1+Q5oS/LbcKR5uoI5OhbNGxXGfLtsprkmbpdfrfgzwY43IHk4ObEBZvsfeD4cG
8qp3JjdJ5YTIM2kggJ/enDRhxxK6PTk4FNtSNK6quW99rsJDZKvEGTtzgUZ3/+ua
PE7l0G7FDaLs5l3LpDLRHzemNk7AXCjwiO2exMnuHlHR+BzvqYG+poQgKpXKijGP
pQupM/c7WU9Wtfk5WCn7gMYBznjTJUZ+RB/4IaDsrfY9sQWrMOZmgC8i1/xTaMVa
2KukHrtq4S+xt14ur/ML6zM340ZVYEjSL6hXXBbcmG6z5gAP628pUFWaRemmbBYO
AfrjQwfwGFn38AOezRjFGBqp5U9DlQUWxAw7g12Nz/0kxI654efcaBudrYBQ13Cx
Ps7B/ycyW3hgBw6WjBVNlAunkvvippDtGC5xoGLWdlAlp97oH0/7m+wv3HYqZzH9
42oFvCM4sZbZO/J39Osgkv508hW8N15fHhfSWIyZolLu0fA+Lrj/cb8aA/uCzOuj
M35yCrB1jmfjYqN7iX6LX6r8V02a6ADdSPDgzxJMM01pdZBJbx1YwtTu9spqZ78A
zRR61mEoaRH3z6EDRleOQq/SficH8DtIWC9taMm5LC115wNLT4LtJkxUOdwU70gB
qR8qI2vzxiKz5L8B6s4115SVXRzeTUL7f1yBtqlt8fjm4xzt1DLYLqlB0E8gVG6e
zwEzgvYMdBHRbW+2nKr7duI9Er7RJ3ci5/CWeBQDmeS1oysWaM3/d4hqprr6DR2p
qzWZaPRD9ACL68Fc4lIEn3EOlU2bi6JPf9UzGV5gyHXJhhva1o836upCp/9MUfXs
uVOFbOSGXWDlPl6Ye33m4M0UXmE6Xyv82mJlVOuT6RjSu50I5ZClvn4g3v6WgXba
CGy/ObSqdHmBuBf2gm8MbWu6qslXMdTVhIPp33s0Pg2LZ7T1TtiiRQ5OU2PlNG2L
ABiOSf/htaKYPw8ajaHuXYIACKpCVjo81ieQLzkTsB6tZzSFmoVdnqwygBXE1O3U
H5b4K4bHXakna9U3toFjN+NLu16G0e573KbmB0/7wePYwcci+9O0WllkDz1ZUMsW
TZnIzK73NyumRhfOIpnBHjzVZHPAVDKqmqPUxS89Isy81HA63/rpO2dwFyAjiVuB
VSm/pLjugs+4EPA475M4O4qJkmQUofwr1MBIMZws7c2mNnjBUyRUcQLyJEPPTDFD
C1KWkcU/YfqGTk7nRfEAn6iPKqG5h85eUEtq37VtraQpj+IGFSLNvbHsYeGyJ7gz
R2ZO8ZU/9sqzNGkQ8ky7beRY0sAFJNmSOzYaFpWefo6tEbgOxKj9SvOHWAst6VIw
jV8owkhHIMarZgENhmC9dAYRsWeH2UpuaY+DZhglw1A8UMjRRlcy3EZgVJBKMRUI
3A2OwnOd+TdMztOUAv+M6Pqrl2kbCfs4+Q8tfUzYZyuUs6LekHEDoNXooFgU/1wn
u+GWshwtjuugVLRwSlGOj4HOWG4rxdbD2hfJSyD6LxFLjnXXhjS73gRdAh5aaKpW
lveBJZU4TBWfHQO7CthmR1kfnJhnPqhZ/sGFkavWkfAN+6DnTFVCuCyDBRxwK3Bs
ck58vxlJ0obFGtGE1uBXdEzVgJwxP74E3KEB60wBcK06KyZhIy2ciJYqQY96a/v/
8M/Fwpk9nuBMqnrbu/qoCVFCkeTM1ZxdZ+nY3bRL3qDDnMqWRfQK6UNBwcvZ2cBv
VMGPa7+ID5+WMNyYvLq93AO+aOxGLL9Hdiy/Ec/D+mEVOrQv+/omIaDEW9cw8fCL
45P+YeqWo2wDOQ2SJR94F6QepE3C+YWC02lqZOZ1IYHeH2QqW0D7WFn9aVP11IVg
kGMV7rIUt2/eVLzMHRxvrH/257ufjdwXcEGjZV5CDcXyqFYk4wDmfUEAyEcV1Gmx
I8uAG2vzACWZSGn+0OSrqKvuUEOBNJQ3Lo1nL9MLG8kLODXRZZSPMHfRSdfPvBcN
aJ43qpXn77DnP8KHWw35z8ljEy4l4y0l+Jbqngfg3b/NOCUWKALsKH4XEwPLJMtr
wqnOC63uNOIWyhwGGz6sozV49BMgFrCGsysMj3IguMgODe382tUhz0eYk1b7AzvS
aWYcHnqoUwIpU66dpbp+HJRJ3YUe9opEmhP4QwNn0zN3Y2f2+O6N9LAiBuIN8I2T
y5mJZecKJS/nM/Pdj03VS/TA2rH9qkERBXy67E2ZgzVAQ6N6zGF5mGV87Hltu1sS
SR8ZCgZoYP6Rb1UPacGynvDLFxTZ4oEk4R211hlsFzSdmpqLVDap+ArbEdhZXh+j
qqLAZCiMpXqTxtmhk9kNLQt/SEVgklHwxpnupkmHWeh/vUSetHMxSLRWI7k2E6Kw
yIzM90jmvjQrNtcpv/8HPfTvzfqcqwzaCrNG93oKJZ18zAhuSJ2ogaWtlxfFFn6R
8SWiiZBSzDgknFYgOs6pJGz91p0JmRtFP4rwlzE2dMutI8dicSsphjqbkwH0wKp+
9vcFkHZcpOUnJkNW5PDBirgR4gOLaQHDmRfdDTluafwtRhhasWw48mEfkK0j3jV5
kj0ulXOcGNehZ0cmN/krUqiHC07RiNamcE91u4aAL/8MA2CfF+Ox397FKyhM9ZGf
p4Mhs9HD6ZBP3epusoTDKYTV4q5oR1tua5c45WjpzdKalZJizY15XA6OAGMXEHHT
HmE7K0DdwtICIOqdL+K9ivyY4a7qlyGDQTTWTxKq7lrNBX5Bt234cuOER2ajgDMW
/vWGMzy4POYe3CIbJAYGnpWFGXBgvCb/5yLYqid/6/uQ+mz+LaaOBw4qk8AMvtnP
Qiw5l0VIzOEqQN0uuH6QFb6RFBEuxBSXyAwaTyZAS+2lz0qKmC+ZAEN1M4VlHeZV
n0OSuOOQVAxcGHRZ8DxdZqq1g6A9JKVA2/wnJfamFmiOIHYY6UG8kg0Raopl1PNk
otf9bEQOSfwRjftqD3PelmhtsaO6+D0+BlcjKtbTDpDRxIBVpnHZLRUCAiriJX8E
h3bilHw5KHRKybGWN6hh0F5wTjHfRPVkAYfI2QNITqRPVeqjMw6vTQrCanIymf3N
Al/kqDN5jROrlwnwHcfnV9VqmF+WFup6lV/LgFK82d3q/EA31QGzc3+vA9VP+5GV
lV9+UgvEeUdbdilHYEI6atarZsKzXTvMI+p2Ilg//uaS9oq3uek8tW0lgPldmWYx
Z3UsdyUbbSQ4GxpemmiPNwW/ZPVhe/JpZyvQ0jXkQGG3eubwJZkk3C6AlVuAdHTd
9lVZvUKXHsagpe1YJBM/ik6fMD3WvC8Mc88BO5t6CrbhutW4S1MWrkn96pT5OHJA
UGYnFMxeQ1vu2067hOImUFWsjo979nNi508UwJWgnS1ghZjxey695lRnA2/LJlgZ
EVGm4lvFuqMSEbKTjcPoDKGmP0PyEsDsr5XfkVijey9yH8aY01kLBszxrVO2dVnV
HRB2DPrY0v8RBe4WAKmw2LRZ6oPDKqrKdd9h9UHOjH//fcDoFSfFYnHkN0O1/FYc
s4vfv4AK96Hb2/y8OQLxTHpieD0DCMV3nmwjbELwOsXZIdWnvMQi3YQzmRnchg6B
1b8o//alvMValt87Pn/mBmqL45yA0eIuFy3BeAEStqfVfVJwOClZ7lbHJd1/QW0y
IARpoqNCEYHLkLV9UqjrD9dZl3NCFjQOvkesGT6Dk9Ju3jLuTdCksRnOMfJyfa9G
WGRVSdWruDsknigdkLBWUNVe3EOjdeP5Btj3/hemYh3uRy5DHj1KV2W6sNHggjXZ
UGROEREizLh0xnFZ/HUYKK9EcKewxQvu3qnFkeEJN/UTH6j8MXK0kO21UdAFnGvx
AEVbhqPNlc9CBPO5wHt2nERMwrQku4vWZ1Gn9ZeKQDaCTKjOaeD9vF8yp70x2IJd
5G623ev1Pb/R77BUtKMI23IIM1wV4e5zk5pDmVQ3yoaG3/+8fpUp2yIPUV0m59xh
O6r53adiIb6T61qRqCw6Scr5PexZ+kdnimt2dGS8GDE5OM9Eh5s4zWH0PqhpWpqJ
alyivVoIYLBtRsiFBQfBqvYhK0AKJqSdHxy4oNIkIDa3EQ1kAreJEXf8nnqa2F7H
wRk5wKZejQdge3OaKgXQHvf7v64ssYpGmC1jYjWaveMMgfPjOPmhYlppd6BcbckX
4Cg56CsnUZKc/c6++TIuQg2FHShAQq7zm4v7aaY3esZn3yN04GN98Yo91o5j4Lo8
fpkM7EY6hmyfOezGUpxvs6wP1G5GiGEFzz0wNvEA0lUVvNeGBMOiHo3UFQsSoiOr
UoevhcE6zo9fhlLslg8JRwtEqBLbfetowrYPtt4E0ponBUyHA7V6KkpC1/E0H4NT
gAPvIQ84E6WNPUeZQ58xrNHgKW0+XUpOYdFM9MmwFSadEOhGVjfCbMDOEbjrNqSt
oJcotEG/YdFIjCc31oCTkk3BgGFifkrIYr4rw2mEg5XYbkgRKh8D/95m+YV3z7bP
ZacJWnaX0Z5FcOlRJV3mKRGuqySO5qYGrxfc7Sa7BwwKLvkJVOC0/sSUAZHfQRov
CJIRNVBAspcJWXaoW1UPCR66BBRo5BGZiMHrQoa8NUHxxVKLn9oBwJJYcIYtHL0o
flOrHPM9HMhgSYD0q+EWG93lAPPDvX6TkWem7VT8zjgTZAwSHr8TI4By17O447O4
gjFpr9YKy1XTv7qWYkriSh+tEfd+ZBxrqhkbvJyNjJNdffmRVTfWyyon2yBX473N
D55g0hF3woihjZXadxvf8KBdZJsLl0Q2To+J6T/7vTcdiahzFhtynbbV+kzbI2/I
q2BK96F8JZGR7UHt6MNRw4CUd+vH15vcuckILRfUSYqZojbNJv7uVvFeqQmhIzG9
c6on7Ngo4yvgBQyUvnxClidHpo0ymGBH7fAxESEfbDj+UJYlN9RmXEu+e6Iya9s3
PV5exwfrNkwuJ+jwyZ3rGdBChQlYN4aflrt+aB1bnZjFE8dyf1O2YxYgo5NP7kgS
ryZhR+dvK3DDoRlhrPJupz2gGcnfhYMpUmoIToIEjyII5lWe7pi4cT6xcyvm4fo+
vbb/CgAQYEKb3opOAvqrhQHmlGoCTkhoBPCZyqe5JNfryS45OUbMBgpGQ+rwQotR
6gxYbD8gFhu0nDw2Vq8AvY5ErkOq65Pqa3KR+1aD4JMPpEFt05UTx6OY93JFdtGG
dAHoQJiiZIopWjYvwDYhwFMum57VM7aW5hF6MYB1wAFiFkFPsVAw4YA2DRn9JxSh
/GarwimUjggFoJ+Cdu5tpd7EXosOwuGJVKmpFBE/Y/xxfm1uUTLhUjIas02SI/34
lh5dVAnCQ7txmGEua9WuyQzbdIP+0GWg0iWYRcwwGciCGFTCETrFiEip2fllAhBJ
Z5T1z7IeXRXNkK7pLlkh0MLJfFNtnl4VurMSxakrh6domq27sT/OIekzOFh33PvR
CvtdHljnAuliYZUTOHZRsPzp6iFl4bjQ2Mo85OfENuPQMOZfjgB3PV5/O6w346MX
eM/XenMosttp1b38vjbdDc1MZPGQgLlztH2Ke5bKRzzQpU6qeSB3lAzbqov4aroc
vzbqNEGTL6HYrHS233Ka3m7J2awxbXFUBUqrPcHVSWmvsqDdILdQp37vofWxmMGD
9DQ+NyPBbnRRVk4149HDbk0ZFSKowxJMTetM0XJhRnXAe3w0hgVLwbu4R1skWiPC
u6GQCuA4Qbt9lmbDmhWd+ncV2RZFnBYEUTMY8motiu7Z/Foc18a+iHpZHVS6m9lt
rC06NCc1f7ZeesTfcmhCZKR7Y2BEx4q+PCukIzqV+s7DPdNUFcM1cBazXq1+xTK6
8dj9wQeodsJX6V66sF1ttjQoTSnhfrDQWBJwUN8/4F9dz0Mw6luhcD2qlbkAnBwq
6omBdzGdd62DdXXGTlcxoYI0/NSa9xZtcd6Xci/qfI6/3rZOGbhl5qcmV/5qWX1t
EA1qL8rhRaNxouDaP/3szpej9uUuEht8ZmgtUF3anPHjb6vNFGit1glPcFDDMtEZ
rbT/EjdkoyrbYxUJz3f7ruugN8/QqNFJvWLtDE5WtcgJazoQPFNNkto1jWoelQEf
0cLmnqmzUNds27Eyz8oCXJGLi02nhf7o2yJF1jFXw601e/OZ9YXXXIxp7y0xg4//
taY5NrCukLv2ESDcaHkM5sjER7ldZESSg6UebsDLX1mdZgnLiQMlPzuZaA96bPRt
glX0wfbTls4AqiBmVy1h4GtpAVNKa5t7cSbOz1Bwv4FKPqE65x7nElsYn5dgFsLs
PEX7qCGFdGmbzajIeNZgB0tSgKG+P9uBjrge/e6H51QMLFiDtyY9aEXGdNRvXNp/
x06r0xRwI5Xj6L4RsA0QR+sfPIvwdS2h2EJK7XpALChzj/kZ32Fh5SHE8KfnZRYQ
bMpKDrJ1inOXcBg1vCLyckfBQWVqu8noDB74RhRnNrPD5BVozwlr/CiAP5uH9yh1
GjmGo2siioIFRhEja8kYBypMHM/zhxJx2e0fDhOxOuV0BpPhlKYu4GI2FtnWY+ra
eo1UoXrb82jk0VUfJL926mPaoLR+CkbOnp3hn1yOVppgh6dilCgbMkGk2LtYrsi8
ptap1BQ/JurCayQ31p9JPzFbmQBCd+6dGex7cbG0X6sgI9ZdWm39L7ySys5X01iL
w0fsS31s8dLVWcHTzOq6JLG1AsWo3yXJeYsuZhRUb15ANfIwvOGMce+ZsZLq1YYl
BFwADW4lXyKyc62KJJ1HVwcjlpLscUL3rlwIkNUMH5KdSRRxZ9AVslZ/Nk7bqfkZ
TFI0y2WMvvPdvjzpBPFd7p+0F9wzkBtmGsULcmbxxgUJeibsJaIVljJeRSlhqs60
tE+KVVUhLlcnyleDr/lnOhe4YzNDd/LYHAXsvDnyFwTmUKvDvrEcjhkrEUEmiva7
2qdLvyg4MdkKifra8O3DfQTDHrkzDF6KXNelrJnmxyL899KGybxnnaO/mv8LsxLm
8WUkKYXrBRe+6nIBE/ZbP6IhFKZLAG4oRNF2XFI0KuNxM8/yWKcWAhtaV7XOzVLK
9Yaod94fnyK7z+7PQITynhN44vhjLZmL2Io0EaD3IlMrPgpWyE5u31qpmVGpupiz
o0Eng+Cq2Gi6ILmNrFijdqch+k/wkwmcFzpjcp4sWuOpMe+A343BIhg4/doW1l37
5CUeKkaTBBzHHeAmAr/h35vY4vhOHvL815EgGGqQnWSgMIQAXsvdTwbyLzbCa6iD
1mGTkbvMCE6vC+5ifjQoaeiCaicPbYcqETK5/mu0IJGFUfIIAIVsAQ1rycBhdGDW
hropcg7um4Z0nUAml5K+OPu/uIJ5HWQD1/ovDo3DdVDhWhdGXFyPNoumt1fxzIt7
IJEaJFzeSHCbvtF+LBlLkVyA8ehpu7xoZ/yBFjcV758YCTQElcOIOZytx3Q1MTd3
aqWKE7Ti5F5iCkbeyJz4lkLuHCm1rCgLWhSWepyxgtba3gI4i3A1bfwB4vlZe5zr
wZyphByJCtQ/XpT8MvPRuALoXOcV4+QLnaRX85aBdka2Dx4gZWZgc/3shFJKwSP0
OcSv7hIfYrkFo5rWv9QjLp8ZT6z0SETwpcZn0injoTrjNbFapjnFciFjNMj2yecl
xNdyZ2IpvAggOdjdvYHKMzs2PApkM6u7sbiczw1Zaj5svT0xpJwXpY6z+6ygIKEG
z1Hs42yVI7grUXHRGpnt1Pl6NVvTIohpZwwAFJitgPsZeZu8/BP9RRTIKiXWhQeI
Pa4TJGLcPjaZGEjC4tVqcDRPN4hdnmOVb68aNROazg1Svju/DBWvr++gDnISefUJ
M/mFnxMzoh25sk5RxZbGgybJBi59dIrnRD42QF09bqwODZV5VMLZNmLXUSC65aD6
oQG8mkHEt2x/76O+LchrnCQ1LVZn3ibSTJtlmr/ANhm1wQU7Pw54484ajmN6HEal
p3pZ5NheMv2VpCcRCvwngBYwEtjjrhb5Fq67gKIF2osl03CrXEzOw/ELLjfv6Sjp
EfjZ5kXX8WOyggfCp9yjI22b5Zp5JL/z+ZAfyoozMBjw6zkskH48DM+ye7Eb1qd9
ILF7C9NVw+ELJIG3OkuyJgdZ/m2VCbb3sZY+hDZWMdNIC0h6BBQIYj1+P2q9yaS2
hEkZf4nd3PVfkV8l728CUMGcRoEZAcvTjSzer2Ot2laOOESaKVV2hNfSQLjeuQR+
SY8Ug8JuceEcU1p5GVIf/GceHjt4VpbUY9bOTcK9STd2BCzJx0AuGVhCETqsoyIm
sbnAW76hpvV8bvaIynGzBAEO74UdFxGwhzIds/BO5uZkMS37NQM+Io/8ue4uP3jB
QikkmyG+xafobAq+KEZFp/Fy8YMEpuJ+BndIRf1OoA8kjO/S08DqHMbbwQ2c3tir
FdxgPqVvMF6m2exYo2Sn7gRGSdXHmwSuopAOmOy239feY9oNLwX4el1ulTYM5Fwq
xBEtHyPVyRqBdo6E9RZh9z6PeTBtHW4+8ct5ajUug8NoirJtdD91TYJU8NGE8OmD
1Y5PrJKAhBYJ4bcglSYmT0GafVqqHD985Jb81ctQ1MO6opd+i3tb47moiJxPEG+C
8lcUqwzVC1oK6/xObkWsWOMHBlB/ZVyVH5CdSiUuCEGWdzb7Tpc+CyXLSZNNEyIy
nVBjcg0M1sMK7DcBJcfZQ3GSAUy7/VsluKiVjQ0WpQbAd+EGaZfnjiX1RnOQyu8i
+xu/aBnnbVdzyYPx9/qpngO4RCf5SkWbJPxve9nfPdQ5w2jT1Mzu4fY+6Temw65d
gZQVaYPRGWgYB0jRNuzkn1J9Zt/sZkSFpCyMy9nAumSPcZ8A8/dlHsokcV0TGDmE
osITgE2mrlrnXsIWiQEYZQEBjG24rXIL9Jv1cX65/uy1IpqbhHKUV08bgcVrjwAd
YfFylAu4XdZ8ojghtQQA1xPLgNlY9odPBowSpg3F2zHpK//QQNZdQsP1AUcF0dgV
tmRvRtYK2iWje3/a20ureR9gAF39Ozm+3iffjQy1HnBis2ss59Zv4tqRu+aAK0di
Y/MeVbKqOe6bc5+e+dQXN54UuWu65DnznQU1naJOMSqNNXydvmNaHgMf/MAsZUE2
qZhmUdHHmub6CK3zXjRMZzzyBq+N58cJPAM0U1KkuFTdGnACWon5xS9nJ3aBsoW6
CDLe2btz+lXJDL2CBG7TgEGgn5ZNJtN5kCeFKLPGqhOC5ZAh29hLyNMvdVQcnIlX
UHW0uvnoFBFOouZOyCyGQUEgSdvin0QnR4O0mie861xBn0ardHR1sc//+CzzN5jB
gpTteNUDnzkIXPEgke4S/2dFEA0nE2cl1fA+FkdtvGUJ3L4mMu9FC2lPI3RyhN5i
AnbC4+1NvyIskOUfGPYl42xS+Kl2WGkWjCoEY4bEAbl2A7Y22Q0Bh3kniW8qJ22L
C6uLIaVIktgURDEfmjm3cv8vQLbA37hORSxYIVleTGauDA1gUtOZ3BDCpJSx4y6R
0GPaVrfVlYUKBG08dsz2kLpqXTkRKO8cBtOkuTCdK60U+vMEhmZ3hd8KHzHbSwRT
ATW0op5AZnQMIyWWKCKlCYBt1j2JABaoPcCjygij1GuvjaAs9mcv9AMW1RGPaiBT
KnTkXX8GvLQmH6V1sefIRhg5H0UkAP2oiMlYYuWuf+CQwVKyKZZBXJaE+4UdDTX0
Xdpc0fq5sJ+LSjFrlU1MMuysMMSJcsrntfmlVCVjJFan/aqUuq6sMutCmbTRY37g
l7j3iubU3yUCdIvWsZdppzaYi8RjNCrqftYKlGsyqFliWfgQD2Bbj0jNx4tvAEfi
ZBwNd8xca5j2An3HKomEHNrDF2Yt4SCwvLx9TlotMCog0PtU0EeBHEvEkIE19lbq
imYzI6vZnoqjMPyQbSSbozOhQN4ffHxId5BXy1xvR9XGIoQocy2ZL0V+tr78pNvQ
HzO0N8DxvFX0NRd6ifK51hsSurs/vP03MNddvMtQUOezKjqZBpG6zgp1RshWGicl
V+PJIcsGulG9dD6GqQA5yfd6lgFy8aQTdHu5hQ3MVKB4ge9tEPl9g1+x8U74YJDA
jb/36vP+xBx8hRDsxUYf8Q9u5mHp94A9e8jE1IpiV2WK7E84p1wbX+f2Nngtys+D
ADMlsrLJmHHpdp4no44LQedljuDl9Pu4AQVM56Tgm1x0AA+QcTRRLloym1Oit5ej
MMyq3ukby7sZEdaY3bfGR7RCcyOx7ptrSqx8jI4ip9CJs+jWsTv57WsZ0zX6Q5rf
d26qq7f4GxET5ElRAthy3RBLArEqultEIA7sBcCnVidOGKmIsgB7Pym55zYaLJT3
r9pZVxjbHwQ/oApt4ta6oBlyCWSvsiyARk4D17FUcSN6Ddex2wkEHe2/P63Qwmdx
UEsBxESrVzaW0gtx4MlFxuhpef/odAVZNVOfgU3WICh+oe2xj8ib8xNTykAK0cko
X8vQkxMULHUBGgepEKY9BOuD0UgVwW0I0ToB1+st733d05lGdCdnedkRvxOw5Z/O
k6jkyypPHabZnwRSsF57TI70n39KqT+bFcKpASOa4bXK4vS6hPItmCJsN+g679vh
7Lr8cNRh0v8pixlH3FqvIY1G7Skz6Ao9E+pP03eR8JR7HzanpNa/lpdhZXqEITi2
qcasHQNZv1VOX6DHje6vGhwtiwJHGwT1I9WOHr8juyaoD8QIGvXeiEgztrrQ3eSA
xZOZRKLmrYfyXZzzfuzOH0XxYIofFeIEz+jUJlaZbwBWsYYYezHUJtoV/vki62SC
+03l8BOyMl1x25Zr0kx4Kgt5bf2JCUFAY279oQK8nHYWDtGMZqazx+cT4Skq/oBk
ObKQEiZtkgpix25Zi54s5LEz6PtFcQ9J/Tu18ZF04DsAMFZK6oPo8lyW303A8+JT
H8W6RRzuOXgVrM/lY+HUQcGXLzMMwnYG4mkeE9rRRd/Oxz/NFynlhUJU9B7XKN+J
8S5FUIflgwkRIIeNe7bOe73BsROwCOsz/g8JK/OtQ5F6BXdn6gxCVZCXyYi1BNiq
xd+GPPCJ68jPVnoCv50V+bkB4NHmqyI2YtcE1VkV6f9GbxItoRYYPXqFCUNhtZsl
L72BEX/L0ZrbkC6aAtrThsf+cRisvter3+w6rD+l5F0HKEInk3CqHF/jd30+qL4C
jQbRv9Ysbo9ZCwM+nUek1cZFSQ0CI+s/CsQB8yGrYdegTzug4YIu0mxVWqbwXS6z
R7f8Pa2p1CKeJHEidvpJKLN0/PhSBtQyIHqvpc8K12JqTl951yWCrPd9bFKQIFmZ
BcDS4a3rElz1EWHDwIhPAnisBw9o69AjdW2Y+I8f+f+UaKwrsbktLybL9nz07Pbe
UgSbmFGI1+AZzo8YAzadfHMqdFYp4Qtji0lSzPYm/qHuQ+OuGxwzXPC3Z8MTL8k7
5hnFFEwMafUYwvqF/a2YPFu/ae+fS51bRsg5sdvh7Eqq/iLus79kA47PtwqA0xiE
iTV6nlAjXcNxbhOGxZ8HBe8jK9CughQSE6Z2yWUcFhbFxY5f4L4EpM7U4xyjq267
qtWoeXKzfs5r5wsska/xX2bS6Fux9sbIzlonecYCIpcuJ3Xp5n8y08BvicyTvDYL
qxLfQbZntYaMw2B+vHII7h46qX/i4LNzz33LTkBj8k+LTpfyLP6pJ6WF4kyTdS0d
y+/w80I2jJwLXFIVfowRfmgBghRELRxZjkUOjociPQRmnMCnvHPFH72ZkiXyN2Wr
Ea9mjvDUAhXmmKfWQEKgEKvEGVS3KFxBMLZdbVlXQZmlB2rWnEqP/NhQWNynygPo
8kV74Ee5kt/3mvGSqFfT1uXbZb23t0JNcmsiTQP/yvtZbi1UKtQ6KaAXV1JvppZ1
/bGieSJLDWbe4i1xmYL81HzNcxkQhrHg+VN3mxxtMRJgcfbzRbVcGnKFRTBlWw0w
s+RXQMQKSuIZoAhBt+WbdB8FbE/ypDHi5iSNZ3pc2Ic7xuxWmWrGHYiV9wytrvqt
LGLA6mik3Lb8JsYr416wrKLX6VGrSeNOTTrTC8sl/Vp/GPBdgEu/efN0JlYooqkk
S24ZWVTPVD+KchwbucWtu5kU3jIIZGHiTVavJm204H/SZk/eSNQqyiAsWo9wtwar
6yGZjh+mZxLoEg+sQUir6wEIvoopYtKRCFj0qDDQfh4Q0Jum7vCbVoaI79EBt9qe
JsLUMIqQ+PHQFgDk0Pb4b4peCtn3MyMxR7mYb91eIYAG2urDyP1ccGsJgRoKzSVl
0B10w+F678DnTYhs84ZrGRieYZUOucjPZQSGv16LH/cWmzDcUHCrJhyRq2r6jKQj
grSfts7KwXStOa2JaWEbGiN+rqY7r6EiWVY+D/M3FqNquihguxttLgHGR1U87JWF
bheEjzFmO8T1/syBQKRVdh6nl/zW4BGVZzpdWKfytVBaNZ3ls3mwLAMxFAog4JZz
sYZ295MNv9ADJVuR3E5RtePFNhOH+dwtukXdfUpYyAnVJUekuorid483KFr22k/s
OTApYOqaNkjvjB16XpntXVRONRQuRkJACUZIW3Dkg/E4MGcdsiVcsljS0ZBl2CrX
F5WNPLvtPeTCFzp0/S10od05IPIfihr1az+fSPTWbF5j0Qs1dMUq8feYtOvLYihF
SNTr5i5ndZIelHEIMvc8graVHkktQ5iAyouZ+I9+LCix6gynOpUAF+oGpYDmb1Gm
TI46njmdkZBTxJ+qMFtHzxogSCN9hNbqZrHOgw+7lKmfVxxdwu04a0YMJ+vV3siQ
76Irmw1CVdwahW+Z7d7UXM84RY6EMZD8FmKxzUEtuUZ7jNO1ewhtWDLjIWm/ll7v
6oj6QfA8WhI6Oh2nqhsrL+QzqnnRHroHBYF7tLzElN/Pw+tLLJ5vA+34fvn7XjBg
0E2mTda2xC8K6dHBxWlh3aWxSo81o1P6un8teaEkPIoMKv6tf9j+pGadBuEKw9V3
idtiC6gmTUAZQON0Gf5hOX6bkh/yx9mwdX0fYj5S9pjOn2epEijCe9wYsvDuhAJ2
62BjefUja1ZB7w3hjtGKlqOfufNv/J0tINasMLOyk5VlF+HpG7NGbDEEBgyBiJ+p
P2Uy969PtMTYeMx3131qKFc6TGtn8sQSm2WIfPc3cHu44MZxGNK1syVSVRgpvZ4e
mCRJepvLJ8cwbVOuUxkmoVQZqYy09r8QrHGGXSzhtRXQff7U5vpNaozsZgP3dVLi
YMes5d8NqwKmRa6stHjv14LxoIrP4BfPKxRtCV1RLN25lddmNSUI1fhvZDek1HIc
U9fhMhAZCZVy5L3cjo+yz44FSidzT6Wi1/PMP5aMlph2KbgDXEQKvrmMwurq8yXS
rvhk7Q8NiZ9cF5ltuOU3UQvOhG7RQXmlirkEHx7K9YpW1kye6r0AH0cH+RE8jWPr
goDIv/9cmppOE4c5sDI4nqZMt3ruD+NVuU6QEtIgGzpS6rBHEPSsnblBMUMx5zbv
xzPRHWpcDoZU99qIbD0iF9Aqz5S4ljWkbbB8q2D22H2l2XRx2ncFT4qWnGMaqPFt
zorZ+L6I2iv5kNEciadWug+68zlzwNmsw59G/2pbJ68J0fRmKFhOUKJOo9MHYoeN
qLAYWjZTsRkTsJvOCTYJSHXIGnSSk1L5iA550Ihi1aOjL7hp5I9oF/8DeIiDhvG1
vSsO6xTTxX69RweBuSLIRbvS4H4fzzXCC7d2kB0LJyN6BqX6M7m3W+xPv8crfxBc
7pytyF4b9+inWM5vDxfSjj7019cskhscsvSCIQRSMYAz5B4afB0Kuq4SLjgTMPok
+AnQRePj3VkCVYW/bU5mbyULc1aKGcFmTuIiQ0jRjhJ5XS4oSMz2V0WRI6mQCEGv
z2ZU7p82MxC2/Kt2pmH42VVcF3vcvxcILcOvErmk3G1b2SECrirUt7u8lVHXtjwn
rrTGGreQrg6jqktQU7uRtYNeS8YsXJNwonKF5m5BA22PrEHf2OKSON1H2iycqaL6
hBzWaGVvmXH7Z6ZKEEDyc1bJoxRM68JWZ0Mk7qSUuP7DPS5TtY+lssgIzbn275dH
jK6z2SkTMECvX8jNL9D58lh0KyTPqqPXxl/rqIE54mRmsHmg1501RduABRx4oq+1
xBuUBd7VKw6lSmy3spr4na5uX9CSyGbr02edZ0Y0XFswS7zsJ1u5yRmFwxYPAvQZ
XatUZtrOWZvufcNNFBcJ2yMTdN8eC6ZAAgj9IvaaQm6N2waIGm+NENe96wJw+3bA
Lx9unDmntBIdcaBuwZalUuXqzfNfQ3W2XxMEG1oWH7qsxkr7jwHY7QziIdX2+RNz
RCkLAY51umR6OtAjOH+9x94ku7KzcbgZmGcAyIe+x9nW3kS4EYNa1husmXUVtzeY
OUc/nv0uTRwwIXk4DYYX9eZRf6t609YY43XjNZcZAwEFAzEb7emBc9osxGdJ+KOz
4X1tHUHStTECSg+6IkAobYgRaiBpOEIHGjO7jgrnMxJt/FkZldsepwswIJOROGRa
UfxfHmF8hiSBOBNbuoEbfqMFs5xZQKyuKSj0pBfuXstdTjXjE7w4/W37jPMdTSaa
Y0i28tr4R2yDomVtcE4gxBYmu7J49J8H0Vu1w01TAFWF/jaetBRnYh8Jg7M8ECIE
+t17d7Fl1Gi2sBmxlbU8mRsW+zB1rrAcXpWOvRXxoLrXC6Lgml7BzC1ma5dFCdNW
55cb475wmTgrS6dNAbxxiUpRmbTkXbMuOfCbXP1LJUHO6IeX3+zUTsg4Uala0b1u
n8ICNdxS553b/1Bm/pz4+34UlMz0Lmf4gPOf5ZE7XXa9pQJhwubsglRsT4TUK6xw
4WtiwpvVxm7Gh+BhPzD+phhRdcnjHarAXPc6JzSF1q6NajCYFbnwfYVrFOBM+XbV
dKBLXvASFxkKdg/4sAPHFOy5qelVsXFAcbPNiKEPCRvrfuIugVGY6VpIXyMWRKH+
C4rfhbna7ChrtWl0Lvt8dkUZ2Xangvw5NkVIg5ez0eeMiuJufJS3hKUDhKF5DPj7
bwN5Ry2esQYsZotJafB19OWRwqGrGXYUjk1Ai9KKZgry9GvdEPhuNW6yc59jk3b2
ZtxfY/GTEK6zUQ7mEvICdjLpU5pSHTCn7wttygvAW6qer+lWxjuhBT8VE2tLRJmy
fLG87ZR+hdkdsAfgjDJUP5kPVZIdrau8v4PSW1eqjsrKSH2MFekV5Xf5bvq9DmpJ
UqbPskXFhQFwq0Q6QN5MC8mwOErDcD57mMcn/bwi8Q5t42NrATeJQ/E+I9jkiEUy
+WoQ8cQtEl6x5NYVj5AdALuu/y4TWvSsQ7TdPTeK/DAOkFpotQPRAv+3Zg3O8h+i
IBsx8p+eJXqrPeRtcLNuuWsiJDnCQuM9UAMkFW0hejZ4uHSF/l1WJzvNhjx8nz/N
g+3P0cU4+Eh6ut1+NXqoSyYru8k2WJqFBwqMa94wVBFQG5BseFk5SCmCEwfr84Gg
ngdUc2+we7d7HGOqZcAhXRHsKurd5VZWY3mJMp6FNYVWaW1GEKaC5D9XV+C6iKv7
i5+dNzx/ZU6PUsoHH26rVoNAjB/vN7fNg6LpHXgF8/7WLzxs5KOdEs4r+5VQycYI
nrsmhg1FyFuV6s9jWz5R7+XDuX/ryhqbAnpfp3Brz93qJrTdAPEqJuz2eVAwpOzV
JK4tks6S9jMpZDWQJ+p7VHAycoYgZNMB1P+QERdF15aPcmbdR+j3hEqPB9bStGdO
BzbRQGd70wfcRtHwTYmT+8XKHjEhvjvlU7+ycB1WQ3zMfiZy12PlL/zFn/OPD2Ft
nSZH/dc69dljWkzf2ypu00MTi+TyIbTJSkBpxOdd2j/T+D12ZZ/Djwta/T0M5aQf
uN4MckoAU51dINuUegqCE7Nph/jT4wK4ih44T90Es5KIS23LZq8qUN4Dnolx8oMu
0Q0xl5ib9j4MJinP/JS06Ya3gT16+YW2rFWFDlYXMMVwqAJX+udAjToss2O77HK4
ObuvNDWAULErOHe2BcKj1H4GlFOfqleGjcwZ0xw1JwdcS7CUXDzXke9fHNSzKDjQ
y2XpO037YezFPq5hsWL/PH2zApuxAd9i0tUAsrDj7AmKp60s4/UYpKrCK5TiqIPP
h8wQJ6kj6kNVhIQsPzkv1iAyJ7Esm+J3bIILHJ2KrfeWphs8pjH1FC1UtxH1zrMR
qieRjCe0EE8TLaZmqBpkcaqRb+DaUXpHXrJWbgJ+NQuq0tjNeAFRdQKkLKTqlbZL
EB1F1svenxMFIn5r0i8aoptUGjte1kOhAxvoAaJUskwc1VLTw6n+fJ6qXen+ejVl
lsETq6mAlNtYnau9Z16rxDV0rTNooJs1tTqhLV+wW+QGWCC+51JFBE22XPLuB17V
PQyxuhXYtk2itMJAw5Px+xxP5xc+SfleypkOchuPyydoWyxhjPyxg97BGXbwb/j+
kChwEErZoVAh9IUXd9VzkNVlzWsL11MuUHNwY4nBR+dlZlGRWITQDQenyYZKrV38
s2TtrLUOc1VKHXcUBb1Va7P9NWzaOp4YLugbX+h77KBQuFcEvwmkzUYqFaKxGPyG
rbMDrq2IHm3SFZqt1/umqTM3tDXZcz38wOI1S3oedBEYY8Lbeyenzgdn1l84SznN
Adm6+kKOTHGstbwSU1B9QbjfnGgYTXilP4l3d692kGEl6v/fKmPwbdZZ9/tCg5kS
dXgMjOg/DPgooHB8ZNHtjB8NdUuakOgVAXDFI19PJK8E5y3xd+iO3DSpEUyOf9/C
cr31rdFuWsydlLRgcUxXp1L7ZHtMXRHM6SvSI63Do2N4uOcqDwpOQDVtJv7+Q1+c
BLF8WvP5yAvlqZZgnHT1xNJIrHswvMphkPlidAvsYpJATfHFddooSIprckI4UK8f
LedhSxiRwD8tEvZdvOtz58GE4fNFrqPlxjSkLndvF8Ku8ALYlzcTd6csN704mYZ8
IORcITHwdoi+s+hcLwT+7K+x45io+Wm7eL1Jg7MWwx3LEfS/eVyCSI/ganX1OfiE
b4EwM+UBHT5EFwtB+oq8LI7uNp1ExNECzderjSSoaoygp7MmTl65sYmO9WhpRE52
LTMCiydP6MM69tmFbPhU7PqlRrk+1hrJBVg2Hzb9bVki865UgcBvAVP7lsrG1nMH
finPG3XmnwpnW7F3W2xL758MstrJiBK5iwa8Z5WBthASVlU6QYhDGBvtOtrHIsN3
UGmNi6A42SoupJGsj3gQWAlJV9qOQwnJOetWMnJw+bxmvFZ6WlbVUWjIAbS0To0A
PZsZp2dl+xTWgWUn3QGQKvluFcfmhzNFk5AmaioJiZiX1tO0vMLeUxRePmJ891ct
sbBU1IxaHEh202N+1Lp3d+mo1Fut2VUzNT4e1/BE9MHWQqrFZWFjSBjM+ND+89Cz
7jOPvHMPS47tlT2tRk9Z2cTPcdmf9QMi5YrMK904sbSwElSGwfrgd+WWb3IZlkWw
QfoMy2B+0fDqqFqIlqSwKyrKr3qlmuETtI7B3/wfVjacPhTmdtYEjnxQLcg5BdaL
VofjVRIFDltpHz5r8NBtjReV7aTeT4xRCf5Ft+Sg1uvwjdN38vaTf3kHBUd9MBni
Sc7At2cyarOuKmxBlX1Dv7cwl36PkJ3iP5Bt/dsw5jBstN/A1xG691sM+jmzN1CP
mg8NhYIJOiY/bjqXjsCntDuKqdUa7YRGWa7C3EXL0OsHglvltG03cNgAv+4ioJPm
JtlFt3tnA8C/reSLAmiT51t3+oyDZvAdNHcfmnix5/g80wqvcj71r6w4IUcTSkpK
sl1HKLjRbyTSG4dqEOFtza9V0iT+aYGJ/LHyg99LzuD5JlOESih72Ie0vOQVLSBK
/SsaGak0PEq6GmIkfWbbni4SrXgneezNThPZEwd7F6GNeZYo1tKkN3Rj0ztLxWY3
n9uLeTCP8IY6RTjn4w3gnH81b1r//ayqAx/BF+UyoBRkWAKug3IFuCh+JOEQCrJV
Bn8tnkyKkGDyBww3AJHrPV3g/4zIaw1zqSFRJ3FlQq8ssq+1SdOX1mAyHn8MrlC9
1JjHHb9ilScWqdGXOv28C/kuO7ccvUtdYlAQU5rZJrYD3hOL6N1YjENWrt8KBswL
qmMof0w1VoqbCrobyBCvb3zCZbbZnS1V1XxBJyLrd5DJKdIYQ7AXVDMGuoe8Loaz
5bFasnWgVWceVPk71tJQ2e4MK9u6VfFC8bLvFDm1RXGA2xRRR4fN32GHtgR80HlX
K0zpEBHYaC3DZE/yPqpg3XsQvjZ3t6IE/Iau8wn6uq2SK9I0Et/4z8lAQ+91yDE1
JyuhCkOE/wCVCm/M+h3ImO1/Pi+Y2JpE/leF3eawjedk9OUAc1DWxF+nWvgaFybF
gGogcqGtZdJxN2wI3crGTEFM5qMIwo9xuPITF2qRqdHDAQZ6ClnuIUWMRjlxy5ci
a84o1Lbp8mIuc3QYxBDLRtZRdv6V5W3+3ZQYaArY0L6bldj/EtmKxY4JL6JX5ZvB
W+LzzQrkM7Wwa471v0PmZZHfWCGZnZBm0oafG8s3gIndM1mGWOJiYOkpQJ2C6vGc
qhBftamqS5HFKXugW44AWkmj0a+1EYSBnW+kGIOqS3yt6y30EHgZNtQoEEylNA+Z
rP4UNFNFTqbmF3lgYFV1GP3APpqMyPqv8ZxN691+yjdSiH1YnfVpjv0hzSxS193q
jYL03gfrMCOCMkRv8YiUcS0vNd0A3kCwgpSM1kq7o/dlmg5huBgzx3R1bHnYpYrv
DfpuGiodnr1nXpimfLQhrNfq7Bo+F3P1zdN+98zGosaWemcsxXjIgQv6aTMxCtWg
a8VSxgIiL3zKC9+cHVB+vDnQMcJfBD2NRbRlhkf1gBNo4uoBFwg7tnbgP6o2l5j2
4VrC2im8ZhWp1kx0xS1hxaCvM1GuiLSmCm31GlY0ZZY/kawYVNqrNfAzMQmtNuMp
EQdjp3k4BFO8I+/04k4G+dgqKBH3c2pOYn6Teuzq7gXthTL+0+Rxz2/IfxwKiK8P
BGyHVtIikcu6oW6PT8sa7rg+a3H57W44la/cJ3EbwzG5gQdcjtncI5EAoWByfi6G
q+wi9aKUk0eKANcUIqSRowBhY6VtggFPvNjwx2nGuDgRNRnNhZHCQSma2K8X72IU
5PCnBAMkOKl8oA7xpW7RiN4RXhlBYckB72XSAf8bCrewPQmzADlbSLd6YnUvwoAd
1XwceaQUXfxuiOvX7sXgc2aK/IcIrU1qT0jMO95pJIQnX5Q08e58Nfa/iNAIXRf5
lnVyIftTs6jbhhd0midvCmv8spcTbhiogw9s5z0Hrmu6UUbIEe02xuHRmYpGYo31
5GOrrPgFNOa2Dq/rQBJi9kXBIhSlxgG8SGofXAbxggTTBhwNGrEoQa+ZgFrMzFCx
oqZyu/Lk8ddVL0EnHPGh7cjPiLpV5neUfTH37+1leM6rZtBaz1pYnPrx6+myxnQ4
v3rjR+97aQf91BSEGfucGWFJPNZCG5v49Q4SzCPoQe7za9C8svELiBgs0wbeqKcZ
JTq4xtvwD+PrnFkOjcfD2AV4vH1y9W75SemIApljFswioMQm8L7BHveCUqdmyFB6
TkRnDTTPJQpIg90XMtqN18T4mUrXiLUMB8BBVTzslU6UdapuxXpz4LAzl8IW+3CO
ZBPX25k0mc3qCpeMFG+DNnv9/s70pQrKh4cSons6pt3JjMaKojvoqQu3Z+Qb+ndG
0xCi8Jb1u4//2KPc8amvoa3L4jnlrDm5i7yzFKROOoJLQdOIyFIe23kOdNhuZVeS
1I7y9IqZ2nVuqrtjfKiD3giYM/eGVZ1ld+vxqA8mB7uC56oJoPvFq6hzB3vIqbVX
AmbAoENHfdUy6l5CMlUmjD2JTpQiPjL+WAtxrDHAPrEG1nAgb+GwB7IkekCY1hQL
ishqgAT/iMOvTfS6uW/N8O28pyj0hROFbyBXGdqfAX5nM2Vu61s+TFv25m+lE5U/
ZxBAZDPBRwXy2qaKFa7I+z6dU+2x/clCDGkqW9pnUHwbzxkawgVvYOdUqCoKh+s9
ZbaEgy4APrthA1TehQ2HRiw+N0OXa/BAv1JvPxzYk17eUSZTbbt41KSaPBSrTdTS
pxgDE6faVMXov/+Kan2Zjq7WKG+wp6cpG38bjBzT/s91w/SZeN3QZz11E5KCySP4
voE8kQnx8OSUCpdrnxZT+t5PiuwvLtVjEJyop0v8cSbFSMt/0mE8ysczXw1Dj0ji
g2M4ZgLyqX7o9LzTE7VemfclAsrsOVa1+/lYkMSP8khgq2bqkZsP8dFA/kYVH7ve
72jbSQH+sJ+JjFFfSr4sWn3DhpmGupsy8GTk++qiRLdNp72HYo7RH1cb+MZrqXAk
PzV8MRB+PJVZ6miMPlO222w4g6OKKYjcyaSpwGoQBe+2cGjDnwRwDzGJQqDUx5e0
M3tytr/AilOmFMmov7Vwa8WGZgp3Y0DxNN4L31/jtERMVLcPlnFk204gbrkpg/wx
32iRmXAEkbhZAtUwHRxWTxKI57TwPLybJbD5xbTtcUF9W58+qA0Ex5a0HI2eh3PP
aEFJb0bkWkMIQ+Oafa1h2V9tO20CqzPokVYRO09StU42OxqS+bT8jD3xgHNffh+I
d9IA/ers34AcxGtyuhuIvxuWmNbCuPCtWtd+QuwTc6i+FhG/MefkScgJ7z6dbkG8
6kpRKRlHpIMaBUO8+zQ8SZGFGO5BCfO5BuPYtYeOfEDDNWBiI0LysiWQImTLwrKq
KuXFeorXXQ2FyAGygK0oYHOoDdEQwDnt7pVwINCwBJtQVFz6/CONF7gvf+MDcxNq
1FpgGITW7I5zwk7EzBlvVQcLu2aH1wk/11wOW4d+m3yS+XLKdWxZVUbpkHnk9mNx
vWMrfrs2sotHRKMU7kJDV3vDkeYmK17jlbfiBuBgb2tKlMB9wmG6xLZ/ATWDCb/Y
0v/+DK5XKg2a4MRDf0nV8yJumPOKhxkTjxkK7TVoJHkvviilHYn0P8TiO6ic0r6L
1tNxyQzv/CFHIhaD8E1HdvCH13nccTTyKCY6ostWIZqhDCUOhoGH4svLGz0t5jJI
HWJ1S1H22nJdxXk2jc8kz1axoVx3xfBblSXcQfoD/+kKCElOm0orz2ESZo3vZIbt
C9jg53ej7Uv3+NhXKM+w5liZeEcc0kmAzujZ1S1yL96ESh1XSGKj0ILctOUkTNLg
YMNOccJTMvcEVNNAlNsaaMgFWSQVH5QiEDNf+ERaeyEcbf2FwnHkLsVXgXuEZUwo
htrMa7KMLCavTBuwa5ocmody34NJXK40eVYb/VGN7smq9eDQ0vlNEihVkltJC5u2
1Jf/OhQzq2LGrmYpnSl4cBmF0GY6U2rp1B8D7FmLeasfYd9e00qGc/z1GOSJ0B31
OKUEMp0ypYECEeNhZ70aLvfNdt3Wfvj0mbP7Fivpx4YIoTXC8oYO/DzHl+7sf8U4
SheY7KYUPdDYOgAh++k0IvHVrraReBWIorSh/kdGNqP5VHpjCxCr5iXJsU/eGrQI
HqlSIiiK14Dkv5tRQL56sLxcvLwb+oIaDf6JQtOLPvVq17ciQyoS6DUJwKxsnZM8
8NNN+0O2M20xvkxMQMsyog7+iEZYqGFSflw3a6K+ktslxywpyUfvjUuNe3gc8Edd
e8WePFXmTsbuA2fVVrlFvz6P8Xh+mMT2sQLx0wZMH+gTkaGKxsXdvstV2ADEKL7G
T3j13YQcXiF2tXyz4xczOPsgCUdRY5hxAUdOFlxi/w/4fSCNWzDvJbAY72uivtNl
4l7I//0mEqa+p6oBw2pzsQm/7WH8mWV4HpVaj/d3EH7Vo2A8Ccc98YD8baRUce90
tVAmB4dewGbpZNpgf7MZoztUSQoyue7i76kQ7WLt+zIQMQhnydQoCKWZOSoND+ms
1NLHm0JwSul442PZvxadnE8G2xMCfzgnSGP9yIn+6Ka9eZAG4GElfILAQWO/kSV2
kYyzHHjqlEB16fayK2yXGj6pRDDky9f73QsONptA4++IOO3JMmprt8UqPcL73WzU
p+0o5rXjJyyw3JbipCZmi9LSaa9YR8RtlkbiO/f8rLLo7BUkyzO6dVmUcfqBtSUj
iKMSD3ndyWkirjpyAYstiuWT3gpCfoVTPVItuE3hpNpxeD/xVNYXyr+F98sD1bcO
tSScxkgVd1ibXIFpop2/IlS+cuaVi+117sKIBZ8Tx7z0oU1RSQeN3r49Hfqj/hEk
LFPoS+VxGzcY6gLtLF2cTyJH3FBtSXtnYXZ2UBAOUbNgKy8s1zfzmEB5X1sk/Zc2
zJqRNF9ni/xW6AJrSwXVonE2FP6hVnlsGNexXw2KxjTLrjUwG3V5Ze2q3Y11/8Ho
IsWgnJ0BYlB+NFp1WP6kehKXqGxplJpIpkmCf3o73EHDeSEAeusUlIaJoldTwpx8
/pkhLlSiOMSfjM6ed5gYk5t+BxXb57kKzgbcwBOcPNqZhOLCeqrqBOHd7CexYdCo
RnXLfMpli7MxIIX3dljQ9e3LofgiLC3ycz/Kifdi0Sur6e386cjPmS7W+0mzZ6Lh
Rw4320W+28M81rlbfuXaD00kX/c4MgIRa9msqms0G0MxWXey8qMCUnmsXiTPvEcR
lSzRhN9ilkRvMp1eagyVJ8ljUtCjh9uzGkGipybCB2HFZUHYhXxyfHHIcbaDooh8
7sluSTDvGyjqRoGSnxIxbvQrjEX81ZGNsvYI+/nVkYGvVenPQAe/Eza4KV0ZvVhY
uoA4XXGOpVji3uk+HU7BuqMnH/iQrgW/U1g0MurHgL9m6WPIXwveu79cZLAEUqHw
ABVSevXWwyYiBs3/YInuV1HQAVyMvyK2pemfWSHgZ/jybb4N69M4R9l5Xffyq+4/
f9FFO/7mrORA6BEF/cJqmDZAfD7RHtw3d1NSRYzQ56vs2CIT6Iy7cfysFdsWya+e
R2HcnkrC/E2KKn1LPnL+rDy8ZWTHk/M7Zt6uhL+vrqKrny1yYxl1zOYsPEmgWMZ9
HoQJWPhwr8jL4n9sEiQr5CzXBNxNT423vCpimU+H1/scFCKZmZrhLb18uG8w7pp+
ObUx5TP+wWCwa+qMMlu8Mc6kdjMOhXLdruDauynumvR9u3GOH91ZYpjLZZw1Lmnx
szYT3EMrW1aNFYHEpf9CUHtl00QfxEqDwwL8FBF2GsKOwMB1cK68y4+lMG2j/tiy
A48MYNNGCBCdjHVFZUWwXdjC1FYl+eyFGHHdiLB+oAvMXVovXVqZiad1uwckq87w
jXUX4kCStgEy1ieVYxMhJMY9lkGcaAE8pom+1IrC0kRRW075a9bvFn951hRbvWeY
36jwtWcj4LcLbBXCcPV4l+humKDL/asm/etSw7O2zFCtV8fFJIzRWLytfb3Fo5OZ
L7SSB7xpMiGnZiDboawdhwMqmURpQG/H2AEvv/fWrwIRC3+m1lIIZal/9dTX0WOY
Tio0EZlAmsCbuML8S20yE28ZV/GTRZHNuWRxcEcnBFz+VsTaWKYMbTx8gFfW2yA4
yKzcISOuk8U62+o2zQQiWYQgV86tPACV9rXmz+VObaYKi9/YVjY/cAs+gK55/GXz
Zam72qyhijOnY43nrA8AuufETtBi+M7KVJZGus82QHezgHC/mjMhcBMGsknP/Bkd
vaTo2HZwMC44qvdY04R49rMbkFWMqc6iGLpD1oWkZ+5msEKacKpicwXNyQ8cURzx
Wc6GsQqfXINVjuZDip/ejBjVSvlS0QYxu4MDlevAxPwBnY60xB0s4Z87SS/yAmWS
6+iS/HV2WziZWfjuAK2Xm6WMRjYROUF0niYCbZITJWaKwGocJfpEKgtmLgF5f32p
ig5qmpEvcuKJz2lIxeuIeJaE2LVEH72Jj6Uy6ux5zOsMzOp5p8pNL09qdJGqo1+R
SMfJrjvlsmJKcGq7EDi88JJYKr3vNQpI2wwFdp50aH+O47cAn71EdthN0IO6qWbn
C57rkFTXmYxLvl4tSNVOImN3hT/Zo55pU/fvxoDSCVy8MV/P3UtZtM67svtwSc7B
BP6pSIGPj4qrrIR9+eTiSPWpG4mX85QAHgyw3fTAlTPU7U7IlyjPT4wntGva7P5H
scZUwFPvsNYgpJKUvmjzxqwiktlAouMdUAQj5nHXVHHtoXihnKkKdDqf7lOZtJV2
eRf+vCh6fgKxMbmFvIRbBunxPr0Vlqvok/Y0Azh1EWy3WCfXDeJWJkMb3foiOKl4
B8kImoxErXIdWZmxJYHdrVMZRSAgaqTrwCi/HJ7lotrDWvgvjFDpjXUv0HwwfO8h
hrsvJgeJawXyZA3CX/+/b7VXrHA+aaOqIFR/kZN9J9/FQpqArA6GkP+qySKv1Rb+
j5uSeA8+oFAL6X/cEJIrd3kNjLJX79zN5n/5xnVMBigQHUDEi6bcO8/bQz2AEg+c
binF7qbEf6Pg9SQ2QLMdugQYF+hyimqMxWKUwlzuzf+MAJsO3eu61TA/I9oHOeAe
+Sqvgddf+Np5ECWYBniZbnvGRaHxLcUj0+jGEeDB33uizEF8o92N16OowRL1WaqR
fmi8yNn36Wyg6xfHzlyP0B3tEInjgl9XrkYjdF8urI4Z4xvizughnwjQ9SVvPzFL
vUo3dMdL0BC+TnDdEw3S7gfIxFkk0MS3Puum1FnNZTnpyRXMP2YEkKtAG8SWc1ih
t1o2EJm1OGVSea0XFkPQVHQHXcYFMbJv++PyeSuVUQm8XkSCg3WME6LYKZ8oPewy
mW1cnHXWOGHsrRf8QDrG1cqGmSj8eR9cNehr/cUB/S2OU68p7Wr+8opwBTW9q7mG
4nVh9zDQeIDIZmPVr2gnsv0ovsWgfX8EnTkz4ZGNnzmQpkIemp4ovzEl8EKIEDCb
s8CcvOQLrBX2IJ7h7QTTrTDx40YVlyjksEPd4id55ZobUknv/gGYMeZK8y6xurHz
zVs4N5TAz8Jqdo1axmBskulCjzDmTOVsUq6FhnCjwpDfsKd400eAgZqILWYfH7Yz
PIu7thAqfSuxcXd2tD7d2AbxsR+/7DD13KlY9LywyxWoArVkhbSZRWhoVAy9sg8Q
HqtQiyixgnIdpH69rLisUI1qGLqjpr6hdDUbO48DAvQVjvqEWq6H5T4uMQP1wPLu
vGIa09wiFIXAl8gYpCxqMqC2+QjC2H1DHT51QT7V4Nf0NKGw0xmGi8TK+LU6dNft
Jkrfsrthv0ekxeSBf7STzSKxQ4CPaK+rGRdfKbJb2qQJ422xjpu8bHNV+l7XWhQ+
OwYRNHHiiu/PL5LDvBJhZ5cVAqne93mOdI4cmAoixUHyZYt0jZG3TdInexaCwl5d
RIxQcX+LPfrnDZvyOFNp1IGwa4nqvguPyfIcQl3QdtOgWl6U8Mf6fjXXvikKWleR
YVfa3eR9pACB5pAWdNQI+X5fgUJCrOgNJiB8ho5OoqP2p1cOX9S08GFQHZLrNEn/
tiqkEbcmtx2kojE0yzerkFXevJehPtEpWNp99xVwle0hmLpFWyyEUSVhVjAXtoJA
/FSP76EQB4HiePn01ViKSz4m8fZG1o519QE+tvimkGh3LhegPkkzG6QwiNmvsDKC
v5+VHEPwGwrEPJv8Jx0NcD9LE3VkCPpvjoxnrJOeJrF+y7ktfh3ydKLiK8vuE5xD
NJs5mOCCbDJjB19vVzAN1Yq0XQ4dbeTPfmeMI3ycg9B9T2ksxrwmRVsaSkRnIfEB
9JejH4ssC5zuJj9IcrSKU+rFZUqECepEY9+ohnB9mj5mmf7AacL7RKBRsBYSpFrl
lmGiU4PUhMKT+/y2644PaIOiIhhI+DD3mfh84dE7kjXxtk1CpAseT2MA0+REIOq6
Uvr0u4GoGLx5ij2M4yxm5vYSb86zLh4HqwnGIXdgB/tImxVnzJMwtibEb9gVM3Ip
yTxnctXMCprPAeFE+PNsyg0Vc0Urd9BeyuxeHMIFMguHZ1srs0S7MRio0/Di3IkU
Is3TcKBgjzv2Yh7lTf2LYSN9Hk5r4cSAgxvnvFUgeOxb8Ru47dltmALPbCDQvo/F
QAuq6zp8VZSZax37zax6gGkONhm/zQiq9T4OWk9Lx7JBAffDjU+8lZxuVOr8cuAZ
T5XoiBjdUcOOLrMHbrSDfeLK/iMXjDrciM4uDVZ8goALsITZaTmdyorcYVzo9Zx7
JUjew5FOXamJCFGWjRkbBZ9hCfqWIouBIZnBAw60m27YFminSVDbZpuDBHRMOWbO
jrbNjLI05zdQfb66swLzoEJYJFcgsTDDXaIkQdWT3kvEW02ZTg3p6hjss9qBY75J
mCZ79ACGH/Hx5Zvon8+PCy+AeMw3+l74b3c6o+s3waUF27FX80s/sVvDbWyWxRgU
SGenGso5gwZjKLZwcCP79WXzSOMiIIphsM2UNPVwUDIp5/5w4Fb3ZoJE5aqw1/rY
9VoyD8NhIj97/fHzynqcrO8P4CtbqAxKLqtFNWMtFzSsSvglA7S8X3bUWmyQYGKa
fkPS6X7NlEteXIXpbA2ZsYOFns/y8V+Yj9fMP+3wu/i++ASukJqgAoR2gFa00zV1
BuSC4CExETn6Y9szTi5cIbHwpAZFMwAOgyvOtzF0rX/oOO1lxURpZ/QKRh8JkuT4
UcYJ/v59pVdc1E9IdlcBITLtZHMB/OZ4Py9Ne6A8mIiGrqukfjVw2q7CB0TMLu/f
dpU/pHyN4Si4Wuc1HSsHzPX5eCmayemyi4kgQDUccHV89qMf5xao17AUZNTMUe4l
rPqRqBWNL8mPxx5vzYdMh6SMpws+Shn7LkZHzw4o2X+ikq7Z/WRtaX3HoFnuvPyq
mnuS6f5nvQBaY5zVWTBRLOaudKIyWyBd74dKpUY+JdpKMeHwSDQMNdx+4Dp2fKI+
cBXnvpDNpq/uc4RjA5p1JxD1y3LsgEYI1xQfysZ7OOyBl+dxKGmcSUe2kWrR+SK9
XpUSlgdI7fJBQSk7xkeugIGVHcqo4SKCaxjg7E4kwMxhMq8HnoTqXWfnSQ2kk7IB
pPML5V/KsCL7D9QHSdiqHSNRDlP/JqEBQkygGw8i4NTokum29TPdImqQs3x59c7T
JyOGjzvk9miX3rPjNWFPzsDgvt360wsaTSa0BTQOlnAzwtzQ8NU9izXlnwDfpfn4
dL+KKaAtgxn1884BwiAOr5d3UNEUxMIEvEh1Zg03jKRdlPyb306L7Gf0UtzfWh0a
XU366cV3wA+JQrx8H+dWppC2B4nqtC+z01b1icUtHu9paCQw3yd1aQbJyzQ2x8Bz
jtI1crEjsGHkADR9IqdB6A6xPI2rdBKMX/fLj6IfIsoDSQ3AkqWP2RS96f0Zx9e4
XSwqBtttDwK4d4cCdl8bUc6XWFvO1jjsmqO0FpT8mqy1E/FvoVzuAY0k1NzQZ+NS
yc7so2iNI4mVGYMbZLuEmh6W/FR1iuQsWOD2Zn4HKibNIySgSs9kKekA/xRZcpCT
Y+PCWpv3Y8je26iMatR4HbQaXoUiwin+T9eUQu2SJfbD9i7I3Prwaw1oSnAJUkHu
+oXIzWCH8+WyrbOXJpaICHfB1+9Ngm+LNHsXl5xNGSkzDTqq4N9nBOShyjgHQfW4
y+lrtrVUDKgHwKId3kvWlDfdw+YPvL5Bpr8zvF1eyrxKDUHxhJTSsdlRjyJR6A+5
tGy0K2z1EncykKojEldsGC8xC0hy4t5/ymaTcmxXzBimzeY8Z1ymSEKcBJY3yjHI
cevPsUPvTJzuSAuegz9KMtQPO6S/EC27bYSQtKRpKV+sYh/Cx71hFLgobZsrtSPR
1eBaNlCgxoWT1YZKVDK8oArCs52psLm8P2Hixp2M081LkfrDEolRH7rcsqfGGWKI
upn/fVY2kXG0aOsBcNub1iHUzzsF2GTjEbJSpQtRL4tW6LGV3cHFi0P0bVlN/6rH
QsUTZfC294u5n0V7f++s7gSxqRmI8dpIdrbkIRRn24H9tmRblI3jT2RuZl6OJhZB
E79DOc/oN5OKr4oodx0PE5cSJJkjp907T+/Es6vT0Ku6/e6zTReaLdrPiNjA/9D7
DZPWCKPz791tvVcN2GHpNBmPH+4sI585CoTsCu8OJnUlpR3YTyBsPiAcMiN22Pfn
7YscMYMLYIak70jH1WRHItG6fXRe6UR/lYnw+vld73+YW1FJIPWD3pBQXoL/KAgt
RekFggv/fDAws3WXDaZWprtw3RmoozKgze90diczvEHF9e6TQyrA/5xPN3nvttOi
23p3NGs1TSd7yp7unHbkClppKIJOB3IXDBapMpNHujL1jN5YUzVGdjNZiXXSceek
jCSrDSkDrmm5qHSNp4zJtL7656cRIu40UI1o7VICWdQYwsVwEsVjJd3NImbQA/mW
2pqG73Ym+ibt5c9wtxO7CKbCwxfmW6obOoRcE/qXXKs0Qo7WsFB0e8c55lbIeG8Z
sSKb7zauj6ead/zL1e4gP1GPK1arrcVvAbdHKDjx+oD3x+enrhIrxQfD6gWrAS5M
UMTC8ZKHIakldKLpCEu0L+DkMrKrp6WGxyF09Gl+YFBnPHhuIqqxOrO3Phet/APS
gL9UKlm25kRX07GeLelmAEY1LP3IhKJDpeT5nGLy7gVJ8NKlULW/jq8QJhl1/9En
Y8trgI5zCttTzsgaCk96r+HP8HzbJEwUSNKu9dO3SD4dwMyhwkep72F2aNlOYeCC
bNhWXFsDVcgOKR6AUF/Mtok2sOgpG7Fhx+0fIQK5livGOlbuQUa0UMmAcIWDPZNo
yv61771z2DxvPSk0i2Y92FqkxKzs0/xCZ+HZzG9sRlQM75nk/oeGzEdGvi/SC1NG
ApQv1YJVjNjgF2FX2yz7d13GPuEWpIcRMv+EIikwa+lcolmLt3KRpuTxMB7Aw/GC
5iiYOolemAMZJxYfWcQZ4gfvrdB9+AleoHH/T91BpY+8oqmEPtKoLLRNC5aMitjw
Dd88/jgyPH/1WcdTh/XNoAUe8ThFzsieG5ZR5r+9uOQQY3gMryqFF4ldUR8BBFOA
b5PEnQISocsX/X3fNVr77RXDqYe7r2J1vuWb2Z1vmoQ4wW7uBEeHXDjhUUKN1Q3V
Ug1ErUAdLz13Lim3yjg/36lSK0RHfepZjh0cvq218Ut8BmIRYk2gEF8vkYvmTj08
YPSrkllwkGqCU/gl/ZUdXL1PseThsmXhyaV1UouRBR8dwlOKKcFyQNuWoLupRAeI
ds+jJeL19rtdXXVUP6HcEV2ME8P9ilcior+I+M5J5dAskTag2QGA7aH0ChKCkFcz
XFNyi5gmYlUEKPT0E1wVDuk2LJJbjAIeKhIViTHOjR8hmh6mnHG+c2k0/5yBIfCy
h2TNZNWPArpN0MPbnj5jqR38flEjQIb0MKWxZHNojbDtV6nS2Zx1jNiJ53r3Rwnz
JWZFUsp7SQHCLRc2aH6O+xlf2QFzLh284qEAdZg07jCCrr8gpjw0TLA+IpYQABWq
O77Hpso4sHgS8z48AAIYW6sZEg+1wXZuS8BYp7Y982eJRwgWd/Pmup+u6ZMwXS+j
8PtpAf9pfiZJfvLM2a8M9TIfuQ5uuTD9UWQIdMyE2kKiqQwSRVwp5JA++6YsZTZw
6OQ10v/VWtqK2PHqkaddWWh4Ov+rWBqcnQbtIfTqtd6zqnAscQsrAlNYeSOLHl8J
+exPGowhR0G6ERBHWY1NxUKIC2jVe9819U/3X/EDUA4cB8W3wvDbe84LiH/zUJXO
f2QcExXz1lnTp+mJTqj17OqjggCUytx7PNNmZCusK+pWLu8p7fKgmsICVM6pxhEJ
9dMimKqIwdZkUXBxQ44XGwwrSgtf/IdbaqR8Oxzp/YN4tRy9c3lJeseLjV2fQd7J
SPLWRy2QH6c2HdesNJ899aJ1lVaI1en8JgrfUpneZVxEW+wNmO9wF4bSZVW2oka+
/sxirkkw7s4SuamQIU8paTdCa/UWhu/v/RWaIvprbYMpKqKslnfnLYeYWpFh9U13
Y1asxfC6WIV0p3tNupYvjV2zir+5Z7JMosAQNsVfqaadAZc1/9jcpfxxWkbpRtGf
zaHtZLKoF8Phw4FFARTMUNCMUENqcpRpFMoRKFG4/3y+SRpIiaaHQ3rUZBUpyrIb
vLzOF0VELEn5Q/voRt3XHuOhGyWd2ITNdq+s44pdctlC4Rc5nB16nmxGHiDNPgfx
3Jg5OlXGzol5FAHmFbLAEPHr1FKoCy5ChKtAbAlQF/Q3oBYA9j0YFodL/ePMvEnc
0iPfpVuS0wkuXq7P49AgYhVEmcxDBB6MuX/iiPL0KK7Z1QlVmoY25R3ufp/wllUN
CGs/bsy7mg87QXtTzsI1pxwWofrYlSXo64i/vHFCOLdgi5N7dEnT7k9wvtvTxsTA
z7r7sIE6V+xigvhi1HfKMEZNRMkxIRvOV3VxlSdBOkDaYOoctpVIu+V6oANWp+tE
m6g3FE0KsQ4QRAAWiHGdpf0vC0ra2gmytPfRE7QJ5We4kWJV8CNKjGQ6YG39WwTu
ioU6QKbz8Jsd0nIrm0QDJiZc0rFO/EvtKHLYbIPLXHHcL+t+rsOeN4RSvcrsWeaz
x523qGG8WZt2gMFq4/E9N7mxTDr7saXi7Ceo3FLL2ABskugy4fhXTLbXwR6eJ8Yp
QA69GKu9lsXwEVSey5Bd6u7CEUh1ro7WjtFi79yGZEaFMcWq1idyYj1qMAiZy7xs
ILhiO31JDMbULzOYsFHo+i673MjjHYI/0EjxirV1i3Lt59WU7QwcELa4WXxHMSq4
uqbG/nBa+lSRJISzeshZqatYv0K8FKDxUiKnD3aKqwDyyielbmKdOG03hdXc9zWv
K4OKSWtRqBtNwqfa3N5zyuJ7VbExyUqwTej8p2CYNq656xOY48ukPVsdwSpbtD2D
fghaQoiWuQ/sXK01LBYcvyn+JTmtM6qXjecu7WgXq40wGqa0CtQmIlvDaZIJCg0X
b3iVl9nvzz682l+mv14Ds/CSu3VxuFp3eUUN+4RhINNprtHpWF6OfYb0IWIWTk7a
GIvvNh6UdAaW1rM36Nk7RTeaFGT3bwHFNuitAbT4haYf+1pzLG+2W68FbWM0AXne
K+RtuGIv8O/Or0KL+XLoKJPFurEwrcwBH2/jSs5+s0MpBey/6jq1MSVf3CAJq7bJ
cEWlfX03dtHJWYVTwmthAWNSD9p3QK4yXfm5S6hRqUEV/GtkcEWrc5K89PirLnvV
g5RwS37G6p3kB/wT2yAHgrrDSUDrqXTFq/o7F7Vj1RQYW05H0iBPY/sCBF/a3uw5
3ouq98kvVEv2W0YUWPmIg5x5rZB7SVEqSMqKdiD3ihvIsoqDMATJg6vyjs9+zcIU
UFh6nxrCnDGIriOEt7dPjP4Yhx0SDsRSMzl/fm7VIL8xeJ+W4GrnewqKtC5PdRc7
MYdrEibxKrKZsWMu+F5Op7jY2lZafPkX1ddGlYbzOPWiRRaMBL6YnAHK4WKNxtIQ
679hcG94HnYORQJhy+vy5e9CG6lc+Rg9IropeXhPox9Ddh0jjjVKrwfvq6emzyQN
D5DUpFMrnM6KEZR/3QodQnFI/k7CKP5PvuPQkVS1w4SR9fTA/cym0VOs8MaKWwSu
t7tBebSwcCNkJJp0rrdH1XfpoVDxaLF3Q5tDV8SYbg/P5Tk4sj5fAAQvJT9xHX5K
NO4LU87qJNKGVTfsp+rRzYl08dzo0bsDIGbpobiWtzGs9Sk8Lc8E9GmrRPHLs5uC
M5v6O4syzbl8HXV51K0XFR2wuC/jmSi7BowfSNCqLUUvSaM+cE3F0hznR5NvzwaU
QFJEjHStGw0mhEdcdgcjF54i07uJsbaLaSSztlgY6Xx8QukyTgSk45LgxPyMYHvh
auiw1XIo9pOs7/dKEjganvV2GSzfztHr4DXTUhHA0UvBkKJiYczpF4RGX5EwxYpu
eTDeA5mZsbXAmrRMRwWM/EjyfYEeBCBXYpzdpVkCL87ltSgMYwBhP4z6+WspMdnz
OUxM+aeZFBIst+QVuSinOUinqL3PvrAxH8R9x4+YBpqT8F/3xocLWiPYITS9yiwK
s0xJsHlb8dKL11U/uvGnw4C+fcm4B23V+dVmE3NT4p42oWrkRAaFSDwI/9CCMhpJ
nH2UTVX3Gi1cRLUQAgzEr/7K0G1q+C9fOFLjGrCu/M3of73wvM66ThbIz86y7vN5
WqqpG0C2xZX08dcj/6gjk3SKAkXsUmoTknujAF2s3w9v8tjp61+sLESaiAAITLl3
G0IpUZrlop/zIgYq1h5+6A3p2vA91D2wCu1ZSO7q2dIl+6DAWClIeo/JESE40Jzx
dNDw+FjmmcRcM9UfNTr7yWSauemOF44+UHx24xriz5DUeEodhHv3p6khTWIUzC7z
QO5RUaqZqYQevqz0wJPV8x312Qk8L1mRlB5FVpwoaPAe3S+eRxxrZ5lGUn7T0nOl
3LJbsFsSw6zmvy8vGx8Fvf//x8eIp27u4JYpwapwsS5gBhBD5m/6HpZuu2iYQkmL
b0PHUB7+apoeK9SnqhmKy3CfwWfbLzwx0vczX4Qh18GACvGTncihs+rYtw6Tl/s7
9jA5171ogJKmpOOIgI2jSaS4krwLnz8WLqLlTdxT60KBsiNzd2wlBGOWUAj6qJHU
GDImikZZXutU24xQNHg76/k5qDWedXt+IbJJEfhHfKqBKOFLBPb20ugEyNb5ACpG
Mf3F/+euekZC4yNRHvwrgnkNVsL9yOLxxndPDK2Tq2eJHM0KEqeFiy1tzEoL6oOC
zPAWpge6MuthBQ6ktQOH4OK6ecj7Wg6/jznRRpEY5tiIeCQPLENvlSMFKAYDz2Hu
2ezDfCF+Bhv3gckEm3J32mgqn2BoYBPApbPBkHuF5NAuxH9KNMgstHcw0cchb+7q
hysQF8q+NfZmSVadCDeVhe2MwAS4wcD47iLDahmNWAB8Zihvpc7a62ucmemQIzv4
FMO4DWjKWZrYTjwOEOH2yySF8jWuVWKJZoNL14yNL2TYzEkRve1q/1ZCXmb3mdMR
rYiPNBgnnGnms1OEfVjLac9dl0hqa3YJtsRuIZoE/ykgWF/LP1yhR6U0QTHaUQHe
8rLZwE5o0LOroWuuRhrgBiscC5kTy8z6qxtQjuXTUc4TsrRMpG3OvVfRn30URRkD
UjD3F4fs3V1spUKCq44o7OeJ/N777dq7Xa90Egaxy5R9b3TPJ8BlXsI6bbpbka7u
As3in9rEODhqhLZFkSAA+GRnkQURtntAgyGgnAFUAwpjNw6czs5WVwockBBUPFVU
2/qIToLJdqJrbZ2FTHkqeEQtWdnb0lNXPboJ1whXllNGrYaH/3CnwXivBZzQf7+U
0r49Ls+QlW+Y/Zu4o86nTQA84UbMxZhEQTJ0lfxG9wHNvZLLyx+SHbNRBSWsuD9M
x0KVrk5I/WpI5MHa9lsQaAgxwBh+l2MfR3TNxm0IfJUCiLSqhaGC8MdW0VcrCiYS
GMHMuh2qPuzJIfV/IP+QFYBy0EdsVz3cRJkvqFJJFbicoiDaa7p8jn6oh/ao2W3b
DTUa0QMk6JnOqFR3OnGTn5NHRlEkwmUuD3zKgl/u4mF6i4HUn2W+Y0T3lVE47wLf
t5vHRjSEt4QqU7KyZe9ofTzWFdMZPOiKX+5yFJzmzdlnWcvb7yi1KH39w87/JDSq
43KvNOVm4AYjNEi+1Vrrii2DjXGXXPf5FczPhanSsQdYL2am5ycCF5b3RCCNtoTX
/KRF7IZzveLFtibbHsvlV9v2lE+ulgJhlP4NNi25EIYoURlDTNQz4dYMX9wEjCd9
gMQH1AEQzFFy6hweMBurmuE6MelAsAYdLPbI4oIKwGIDywoqKuimUjxd6umw+xDA
IpldbQwHd/yhFBS3O5iuYykZuKsfYZSGvZXSdmsdmw0UZao2ggw9WKqU3yqdr6Cd
KNidJZNX/w8xEuMAiF8zWeZO9T9WkqjZBtnsuJU2mNaSaVPcrFqHggCragiNxG9a
3anGmgDCvRAfWG34Z3cFks4lMB1jZ4ZFENk38+ABNYa+/x6b9uN/4Ta0uDDbtIhh
J5t6d4MCKnoqOEJsqHL4UGnsipyTY/GzwwrX2iFpgYL0TQ8JraH6Z2OxbmvQMNnM
7swaeL9ZpIdBPmAFI/TQEzMBfsr+8M/1YvIb579yZxOWtQPtM7rzaY42NJOKkkzU
Rc7x87GTpz1461Etsw8OBD2Cui717D4KF2hglfAimY+q/RMKvSraurKiEGmt+c4S
jm9rAfKZT3dp0/1+TBIuN3e5x9ogd+VjllqXz/ZTt0S5/AOviGZyEr1gYDt4OyZM
IksJ5+z5XS3nzGZPw4HHFXIV0ioZIDCxoJI8GsArjhe4VB83Z4Yfu5hUD7fqytRI
MwneMTEQASW+l+b7aCFXAQFtooth+wQbJVo8RaHl174BmB1qqVGX+pQhqjBjKWaf
Lv+NwzPkiVeq3PDPissjbgWyOjgtuTmYhP+VbPF2NhtCDk/lVndm2I0psIqfrged
dwAQ+hGm3D+qpkbDgNbnDEJnH0QmRqENLRL7Nt+dkF93MqEnqQe3vq1y4XQ8PKyi
kRjAKYlZ2Z0Zv7nO8shVMgoFaKM2OVYO+QfPbhIja315etVSAJAMHZ+fp/OoYIs4
8v1kcKvp82IdiziedG3XeEBwlghdO+JKf4b6CwWG+Xg82prr670b/5hr0I1s0NSS
xO9QlB2cEl8rqB5sIRvk7LhI2xyH4Ur8tX+eduRa+As=
`protect END_PROTECTED
