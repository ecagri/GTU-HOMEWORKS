`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UdBD81Qgj3lZ8ZEp9you77d1YnzZfU2C5kDIJd9uKBdgngwHj3kkTGcbZBsEZIoq
sRRqlr2vwxKnkCKdTxMlb3ck1B6QS3+dM8JVZjm3MDfkhLBSRjzIbaoxp20871mL
CWDVEnLMJ0/eusuh0bzG2JOOt8zK8rVaFeQv4zj1DnUg5A7n28Kgs7svjHs5KRuO
etfihxkFbyA/ajwUXio2BGsaTmFc2FA1zY3OL8eRqsntfPthqiYKg7ZtSkBAuARM
ieOg+xgFgo1+dzAYIGgsZLEPS9xoTBRleIeOtiovqH01QMmxL/cY+LWV0u4fjYFA
6jmb2pI++zEk5/4A3E5ZOPxrweYEIvC39X0Ntl0uHLr/7TztBGUjEh5bHOTqxOrg
69YNO60rtyDnG3oNIckeYduHqpj7gYje01y/pciAfkKjHulqLPXzP1oJcOQMZ3w0
eP2WSd7laRaV6iqaKVk6zTwfdgHHQumkUdhUXJr4I++mpBEkIWLemYAq75snyMOz
3uXZiXTcWMNnLD7EHoVULtANDM2dgjV2T40n/ru/1mzQDcwTgaJR/hg1kmiZx3zv
qZSJRkA2zcCESSlbictxlkbMML2Ag8VRsAeZ5Oaj+QQ9visEAcMNF6K1zG2X4Bt/
NJ7BUpIgfFC+EEFN9Ggsmg/K48wctv5kaVRpno3oZSyl8TFQLTa9s3Oqv1CcoCUG
Ypb1VBRPhnuT4LKRYQImM+N1hBGrEudlC1DBBkEPp0f+QtjbjLyKxA7h6X/PmE9k
BU+SG8/e7Y7t0vdQOzPx9aP9GPf5qmhnxYrF8koItyJFbGb/ity+eBBHiuWrm8JZ
QarPgcuZaQWa2WtNh7DUCu5t4ncMRGCemTBX4sGYK8GhN5q4mrbf2HH2/1YkQXEl
K36EHJMKiDqEVrQW58hBpOrod/a7BLc8FmsdUB4U/oObMaC3GBse1ieT7VKMl05h
f/sita6LTa2nkOMXAI2N6StsL9kWNYI13XZX9i1WXdkC1Wc1of6pu7ZklkJ8Tb+y
4OnEoRh4K7+fOaAyLEgjn7RNrbfPAzOTo/DZLSwYHCPaDBn1Mep7sOwjGPqmto/8
ANyPV1WgNwnwbvIrOizaUwh0ZYWsBPWOzPGaEu/HHewebytrBH65pUPWrIdrrtHc
F+ApepYOXffue0RDuE3WRZv767p2HEpks1yAfySP5PKF81CjqlsZby44DttB66vC
`protect END_PROTECTED
