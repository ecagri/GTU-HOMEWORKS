`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3AMRcyKfHkijmgqqgQAMJ1BeubFaxN+ygBHw8dAohNFtzbFjDtKW7WH0tEW5YnRA
PhAGP+8C/+1TIjXxxFOL6SfKM4dZQlQPzyCdRlbxeMZTbyZgQrtu6vJqC9rs+vOv
4g5oTunxJAgjxTL5hyQLGGS133paWm2nzmDt9SIlzxpOaLqJxDtCgAdrVEHrBoJG
z6R2+Y3oEyyu2Piuam1zOg1lfGSWsbZ4gNMVEBE92gBL7GmcPsoXLj4WmQXcYnhA
L6N9rN4iRy1uBN5QEt7bEYdf+FcfRycSkAIJgvc+LpJ9HYI6dPF3s6FSJhFJXSM3
usOWdxyT4eSSLGpqIvDxRvKOjH6ai64ohbxaiDK47WftC3oqvETbIUFrmL4pM5j2
kv10NUt7iDBmITd7wIgPbpXXQfv7JXZPWxcsRpADLbZc9ub4JazRrk+1XMFznLC7
g4ZgHAb2jTXM7qLWLeSsUT9/bnd1zuQbVhffflyeTcYL0Ns6YivU06mDLwqDIbHN
oX65O7BZGVChteeIGaN6ELJ9SwM9epCicNl0gLmJe1KuRWGKMOSj/CqEnJTWgvI4
vvJDny3+kT5BfMeLVNxmLQ==
`protect END_PROTECTED
