`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sdoVBY8gBr5tmHiBMSPp7wospF2afivicVbLP3omsyVyUp4RCYZk7bCBybIplPKX
PDAWperb/h/bDRzsJOvRMdyPRkEE+vP8FhH0DHDJDM8VqY6Gg93sZ8tKNAePQ3JT
vZ2AtsAfXFOR8+XAG66qF31WP4c/h5RJMV3SVlhHQIkDWyagew3XC8tTHuG5xePB
14TrtEPs+Y8f/ifBqORgPIDo/i1TtBQudiH7zfqZMxlCet9InPKfMJ+UaqO/W4aR
hZBqTgj42KTMS+jDS4N1uIOrLwHZhzKwyl91zHxKsKm8ygekqWoo2dTViKGj2yW9
rTl3+hyUwffA+9z7+JznM7jpc00kK/Ysp9rC2avTDbI9a39/UiWXV4eDe/1QCWy4
CSgQKhUF2YlarN+Z7xJR+uFHpIhYwfxJFBcdQoUpwRCUg77kKrhdMAgQkRF9IQ2f
NZQork9d1sMCLtYFM/I5B/0+BP66y84E48Sl6zRg0i2D0gJ8wPofynDo4aOIar8z
uygeaPmsyagXbdNkoHWofvy1/7tN8KtJqyf5TtlM2+z+MbDcei5jUNaVAlL2MF24
dI/p5vCZgvlY3eSwm48X7srYfxDClbWqJxOCtYX3kWJNE4NXSgi3aHyQRBxrNVT3
tgLdqIAktSfmQ7NlPakMCNviacdAmmet6aAd9ND3AScNbeqKN+76FAgd/NU+I/gF
cydGD0MMh6ciitjk4xxx/74XX9A6dN8QUuIwRb9IAuj6c4LOodc2xPKptx0jjDve
gw+0Trq7ATG6m5o35278Iycln08JrOW5V8brPptTRitD/cuVBhFOEH1WmQOetdhV
9wsGAOQ744pmCGhnY3WDvQp9VBiGQIZEp/qX3wC0xfr2DX6xKDBdpaCkHj9vGdBV
8joTxQF1pB8ioO/pfNOy/Cfsb3Vuz9xkJB5WnsE9P0orFR3UlACAfmlMx89OgSaM
LPkJS2NCdggmb1fkL5NNUg7k2+EOU6iFCJWb6ADr74PpNbdCRBYVzuXVbysMIfXJ
gVE5qzAuYzz1P1sfyJ7WeLLqAj+wlKpxveGJrIw4j8Woie94EqFhx+dJmIPNUJof
CdkyA75oa0Zmhpuju5ct8MGm5/2I9T/lML5MuwZkBKJUUsmpHgqGSxdIroeb8b8U
30QXQMZf934nLu7zikekSIoXU9ii8kZM0BmXNRcIGFTD4G2aR+RihvYdcbp1eUAb
zycI4yC2G3LxbuefcB41BccJQnPQ25W6Mi5BSo9hgCgBfhUEl6NSgt3MFpQ7ixJO
v6PSZCYGUpa2iWmcwHUn+OAhIysj4uBjd49igI8YL7y2zuiGpdmDgOkjM4xPVTYZ
Piw2lpTtkqcgalAZ/Qrb0DvgK7g/uGC1EjMxRTIBneay2lK+MGEy4avq2KXfPjjR
2ZgmGjQvR/QVPDGpd8Azwx9K2JXcqScsnCIojTIF+eWnhQQBJ4uBdIJFSUVni3VR
Ak3jEUPqqO3psrNMn+AboZoRzE63LfotG2EC7wnE24cPqvy/QNqPzpXuGinIYK3y
Oe1rlOEJ/zY6pD3DROl3sSLsWgZ6YdJeqvAz3ClqmO7UV3cNVQfTZ7TKJoevRKmp
GjH8lTbwJ0TA6Z2rFmWyDV8sKRvbT/LuwCJIRery5YGtfB6bpUo37v2Jt812WhKn
JOKwF78TodvB+KKhjWvvOMw0B2J1ZGWSJi73kYKzn9f3qLyTXCkTjGUYs/Ur8M61
vbXjdFyzzKdNqiI5eMl4SOzYJdHn+YvRpvBsbcZyfPqThhOql/IMhS8GorPLzDvJ
lcUvb4XbmjRQIKhg97IYIPsk1eEGnTrO7uD5pIYinL+D5cRLwQRzBqWdvdHl+yhi
dE+PRREVnzp+JcnIlVPBu/qrTN2tdsymtmuDoH5EjQj0W+RkEdI+UzdDse+add4n
1VNFLGfpvR8sV6NEktPH0B8gpPyNAFAM2IOlKX7NJmU3Hni2iQlINZDwxb2P0MKz
wr8SfCMnIUEjNEql5w6I5T6FyjDPzuzER9p5uPrXsDIM7EDj9/HUYE2R3L+GaA5P
QMD1cQ9WMupsnGxikzzwVIUiDN4V3dDGbpOSTagjKUlOcQzhiOBTGgtO4NOeDF8c
dsJ8fjyMaKezpyjKqbkYOUxtO0om1ZZxaXecezreBf5wTwZmWXolC7QlbkOFpiEA
WV4ikvnzatwF3GKU/DiHrL1A8qhLChzaHWXL8+Awjx1eW3nzhlLiUMbHZGKPZZEC
N7Iy1rs1MO4+dPyHdRy8g4qcSq6aH63jXiUZvpWhUykY6mM+UMUYZd9B29TmPmMb
WAZwI02j5fR4+loObbdXPPvQfFhwtCx1pWVf4thwjnBFd3wpDa4fN63LLXOqEwIc
2EaMcsbnsRXwei9+Hj6HJ3ftmhFf4iMjjcoZtDwhBY0jlYhtYLcviD6AFL2VUtaI
A+6C5KpXWJ7C/EQdZ0jVWgTyZc2eCazMBChhFmSfQGSkC47Xgf6cd8jXjt0UbrFn
rPT+QhgcXSiRPPoNfC7dnRo7GGT2kqtMepBZC2/wiaqCllyUcXx+WqK8eXkp/XaS
4ElTi0DXwfncL6A+ngFMiSqS29BPQktft1AmkZSAnQzC5SsZ/80FE/qn7wHGqyfG
m6zZZ78TMPDBpqthzAJOGNqXplBqWWwufDPowyj4TK5wV+erSugS4jhg0KnPfNJG
LtBaCBixgNaIrkhs4f8HOTstYjC896J29NpdE0bE3HRpZB+V4e9meINz0E5FwcHq
xiYBu32m6bl207VTOstl7eK4DVNIoXIM37OZNi0OO5nTsjWMoXx/M0cMsVwzy/84
EJSzO7sZSvu7D4c2fspNBY5kr+fjrmarjijNZKEASXERkoSlM9XbIGfTUO40DgwB
wgsnmalPHHjfI3kDsboZ0G3iI/8GixodsfQ0rDwY3bmRsjCm+QSskLs7VN4C405F
qiyg/8Z9SA/ZoHBrA+HJBCDArrAZmyeswbzx+m8MgD8IuYn1cERgfvFBwMGeSST0
TTakc8MwEOXvcuIBNK0YpTkeIat/lIA+su72yyY3BrzevZB0BHU8MVz1FRryy1gc
W++iPmC/xUT3+7hOjydyao7XSY/F/gbk629vRCYY1PGqfE7VUtr9Am6DwnrY+HQs
IkJ8B0VfpXNvXu5VmkSHiQozs/WQz4pSAy7NzH7qu8DCu1OsIX/u9JpZiH9GORQB
1eaLVFR8uGQde0OJPxYvwyiCBVuHrgeQm0WGQEJYTvyYgglBXKh3cQtu/a9erXNf
rLKscfnIcpTnf5xcqhrnlQ1PLvMIQd6wNe4ztK/dD5K+OSMzLwpsLGs+V22fEta4
cdlgdfBxYK3j8ERlciW5EK66iecTJH0E7O0BnQNxtOgz8dbVuBvFynsZRbNOfaHC
/030RP0QvJ41otiTDw/N3sgkGGbLqyuG7UksfV4MBDaV6KC6YOxhWotiLWQR/qis
Ml54pYvT9vmss9T2sMJLy9A3QuPcpkJ6KuhQYvRaHxiPDrq/2Nbq4EeAEoby1OG0
`protect END_PROTECTED
