`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aLz/luOtRrwVwVR6iP0+P2WQFl2nlCCONyP+6p7fVMRwJ9bD45FjaPpX8UdJrVbQ
3EDh88d31Gmf8O9EWSYdyJEoPVWw1Q02tFmjxxmt8sr0GpLevtb0oGtOMoEVmGtu
h4BDXOB4gBFDERKdrvUDPR8Am/WlWDSQNpPrVp09G+0oMapecX7tR3Zf8u0Bm0Gn
gXwkOdXQ/ezy6oKLsl9xiqy4bv0ziDWlqWfay2Hvsx416H7WLRsau76IRGnrVQNZ
cmxm/zeuqTOzzZefWd+D0au+5gCyw21IyVXPE3j1oCz08l5gxfxcpRrZb+GhS1MQ
6t0IJVM4n1Dp2saOdm8J/H0vs+GtZbf6FMWSc/lGM2XcbYaXUqwGCENA833ioqcm
XkmNPSOSk0k2V34yu5BQo+Ry33KXHi6HFmeulx9Fd4VpjveA+VRqH1QjXxMt0pbU
vCE7kzUR+aXtjcxwAyj6nC+XvU3LHlfeF4VBmKA6QH0=
`protect END_PROTECTED
