`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JQh/8gZ+tUhAzplYG2yHtvHeT7/XoBAheygIVuAlwpEKE29D2I077WoU9M7kDVip
LEtE+T1UOxeuCNnPo65THUBslOtE38+Bfm/wbiTTCNPKzANGGloZUZbr9xl7q3mL
JLY7WmDiXxYnD8R9CbQi+YujbVmc+iZObHXPpnIr9g2Ofbq6kCmITKQw0YcKKX7M
CRdt5QNck64Z9eE49dP7UOs8XlIpryyf5qCzj4e9FAWVD+IR3d0Ldb9wKh4m5rXt
pJFCbJ/ZJ8GS/e8sBWEjHw==
`protect END_PROTECTED
