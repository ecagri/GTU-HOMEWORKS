`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q5k9SIHTrZzBUAcaufq7vdvbrCX6LDM8b6O7ciZrf6LpR7PBzpo6yGht5lBN9sp+
gSNx8znPEnd5iU0LKRvY9zCJtmAahcLCtpysb5kuKxbz0oWHaP71tUNY2I+WHaAh
bjCZz7jVIreM6BsRZ/jfxeKKF+ZU0y1mT5Uqsp74+yTLYalQFejlX2cr2hjWerT5
MPnZYhoi9iLrVjKsaT9S5E1WrZt0laRBlpBWz3PHfzdJk1ZMRspMYUP23Ls/AnpD
Qk5lshZpUxR5kp9j4SzqLtvD5F3sxv5sGAI6O+jww8t+KsSljk1QyFDZEZgXj+s5
IfzIdCYdVg86zxxzxwpC9KVJ7aiwdbHzZqW5OCulp5Xt/+Tzk/3zzFb8bESneNF0
jHR96jdI74IdoDoOztchsZRBO0zyt09WtMLyshl62gFiOfg5vWlmzdcN1n2Fhj6K
aGc3YolC4r35Po7NNS9NxBcdBnwvpkAjo6B2mez594AplEt3mtosq0irtILsPv2J
9W9peuhNDR6P6Qk+hlrxOiYNNOZALGAP0HeBa1dpK5ZdXBb4N2tFOnFKWs1WyuUj
W/ol2H6yfa8HaggtZFibJgarvbzHUALSufbwAU/avIDU51qPLzYhEA2JmTR/ZuR9
c366OUx1xk6U6k7S+vgQ5ZZq6UeFUmyaFxldI/Y/YDIrmAXUKT9tm4MF81wmgYQb
oAT/hZoCcTS+t1LuD0l0WjbZnSGIOEsAwga+ipZ4JtjKTOfGX7S08XJgcJ9i1qgA
3kySL0AxounSRbsYR+BMihVhkIQJPWLRp0B/MDD9PjdDmwFXTe29ZS+fKg9vOLRD
+4lhgBN29VBx7kxhAhSKITKXITP6hNUMP+FxCyr4O6SGV5f+vqSVFc0+DEs9t4RZ
w9UOXKpz39xGYI4nQef0TXHhMWQ2yqSbn6JE4QkWU1t7YuEnzjelFbWXC4yBm/To
FwiEssJlGhDmKUwv0/4vbm3qDGL5yLI6bbaeqz+9yI547Pl1wxDOpdtg5wT08I9c
bkzH4K1vTdAFG3O6vaisjIGbOtplzY0LvjKm1A8pjQAWmfvYQZ8XK7vkBGfFhyyq
QDl2IdzOI8rMd/QNXsVP+6zdh45hv5lBT7F3Atc/7t87OXG2TDre3c2CAl7nMxkd
ziKjKaksHqIePhUhIZ/yr9zRrP7KwpMUJCpalWbEV2Y=
`protect END_PROTECTED
