`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LSSzRrXTRVnzI4XJ0OaP6SmDM+03U3l4SbCM1v5hdAVvkBQw1qbua7hbDk3fFoV4
rR+cGz1yXPFcMWZ5kC9Bh5hhzJy5G66Jtg1vXF+lgTgtYKA229RkCxjKBsJ3jU4C
VEwF5AU4s2gtCH/xEevmjw9pZsftcDUVssvH4wsRC8C/t/l40oVClVGaAH7KJpj2
NzN5/S6H2aAeuWieiVnJRUannAAflnWcHtg3VFjA1D1Rz+zLta5lC92Ki5wBGrsz
5xOsBMLVoLLX9W5EuVf/zTTBaoBLqwA1bIHSBlHl8qndjYx1exaGQRAf3n4g8zgt
0Dcwa22HiRlCdczgpWKAQa1GWhcySHaqF4ffm6EaU9NUmQjO+XBD+UaKGl6Z6ytm
O+lvbFfHPQ+s8BHvOib8F1rutNVyKa0v7tNyURtHk1WMpYWCx8VNd5CDlHEEoS8J
f3abKrsb6RTjTUuEcFBTQaqb/Ek8n3q2fgVefuccHcJItRm595xL4V6dCqpalXw9
8oeV/7vMZjRthzcntkG+WiBVlCrOCHnJ6s/s6w4FYK1ZOvDuAgQSVFLYlSXDIAi8
+rILUFEqHo22WCq1/6IFRjkRacdKPao+9g8lzhDHCDRIMpqQdbgq5jfjqmvtg5Y/
LZPyX/FqmtYXDTYdD70OyJpK7VfAIe594sJyersWmQ+QThwl+3AOQQVCI+PTV8Hu
ILraZ2DvUb7/1YfC4H+jCOFLDJznRhLAThOq3hQFJV3sOL78AU71Dxpx0x3OFnYe
zG01qOWLPcC8P94uy/rioDu0PwkZnZYp4OWieKYWukSkfEn3SvIXcO6H117iRE7/
us16ZHWrJxlkpAEe2KXeiEQblwa4iwkHe3NT6IK/jlzKN2M7a6wZlY6wp0GQ4W6C
DgsKmcOc/YmBZV0weK2vNP1RSiESRqoXJVwTxXq7WdUJkJzL+HBsCsOEiiHGW0J8
2wvT4ZUvyfGuEGKgkPfEwPgdwx/ce1jumcPjo+Y6LDRb/TEUpnThV6+bAi7UIyNu
SW84fj/6q9sOQZ7wiPYhmLgAwSee791E3nmnJBWDOtUp2Dz8q0mvtfa7E5NwztOM
ELlirfBPJaQCaLg4ywCGR0VZzW58jKY3qBYUMBd0Zm6lC/3SLEvhkuMEfR+5a47v
VnUBT7i6wHo8xbwr52rgDU+WVo2QVCDitRuiDrphHCrva4a0170Bndrcr3npCprC
+4uyPO+J1fKPT3j4OaU2hqzc2O7eZ+kpXjmFOhlEIzghll4RfIExEwgTkbQfxNav
aafKjNtkVF3n8UR6JzcRkZg+pOVUW0qBLGsXbogwsMTDe/Rx6cZY50OaKIwM9o7r
SfsFufdtIlcoXNDe6qxrVNml/bhmfhb9lnufxR+zCZ2X1gXzoqz8c1s5CEF1CN/O
EsCx1SDEIZTW38JgdALvLoNBn+9yw2kqAcOcSzZNVkswGga75UKYzsysC9iH/cZo
4zifD6hXhjGH/zpKefH0/+Pw5qFq+0reEcD9+xSVWRan+8RrUbZoUaNNi4/Sdwa4
dkEy1XB6XpPo7hwbC2ravXQFmTMNjy+lbQP2MCRXvsP4Z1JMQw+TLDUfAnkZmKpL
bS9aRkIkhOnm32g8qyjkjfgMcBP7xLrE72EJuHK/2j4sA4Jzz+rKN06ztgEyMTRY
rTb1v86L0UL7nairQJ9N3fFWwcTCqusWB0RmTbVNycpq0pIhk0G5mbVnKBDGzAEA
rOcn/JlqGGclYRKvXNhKijk1zIY7caG2hFoijOQ8nUJK4ip5cGMwLJjKeEtFooz/
CqQeNPi1cmw/F+DTKPiwiza77UkUhlqXEyJkhUnvtq6oHnkoeCH5lcieSFyeuFV9
/BwLs6eCrWSHHDDzZIq4mQFIBrBxyBdt5DOOqF7GPJycl5wEeyskDDZB/kYKhsqH
xsP13RNINRaS+l99AVzbyw0I4W0GJaR4YTQ3m7JUaLq47EQt4nkhh7YvHBkCdveW
VEgfC1ortXZmLsV8ErE8wrz5vUo+iRjz2sxxAk3PYa6cSHn3HOWVvJGiKIjreKT0
Xj1iDLUxiG3UQ4WPwFnVs0DZ0gFlv/ESP64MxXP7eP6uULxDBuvnPGhUMp5SIeGu
am5J5bAUWJwYDWoIM4KErvhYxBotRcVIKfb6E+P2zzz4tdUPZvw1wOxHQlB4VU0A
t0fxT1dLwibkpVK99y2y+lbDBJ6XID9ks2eQmUYI5FroOM49vRUBcke858k+ShX2
EJpwsTu1eiZawFWyYFtKgSJARs81+7ZWK+1KD/cXGlWemxc4vVFNOqxK8XBUnDAv
Ij3d9rBYZXxD0Ua2s+UsuH7pW8QR4Ery5fsUIjWzc5I4sOksn5XmTcSHNk/zGnPi
kGdFmFtrh8p67YaEFV1v6SkjkMqwbe8BWeyrfR+qBa02fVk575PDy9BPXtJzhiAN
YgMmCgl9NUaiiSuSGvWpgdyXM4MlEPTiCs7zB9WtvoiETFsqVj//01yQVKyI/Inx
qSK50lAeJAG03fnifhllIPhBGyOlMWyMVtM3JBiVow2gypR341pl43QRMLImsBUy
p93FVmLb3DAQYFSvyfKHK45Q2JzuPSc4S4uL3b1XU4DyUjuIkcJLns1dW7zqdjt2
3sW/d6PQJEl4niNQEyckRMMydszC9lmfNHldsWLk03Qh7o5rQXV/H4Q56hHNuT1d
NawdeISFBfqsbDFtPTkzNMQjAUOe8W3AIhiKnsnq+SwhfHC3q1N8ELoMjFde1c8p
CwkoJdVCvFCKXbmfsVGl0wsSmdEGMydJIygGF4WU6EnaLCC8Vy+l9wVR7PUmtTw9
0MqwI8Gi/LkACk+0s6PzXv9F9XRCKtB/NfUfFhEg3W9tkHD8+YsvHOQeMdbNBnD9
`protect END_PROTECTED
