`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L0H3ob72rUfMDrApC5G8yjdrBIkP6gosQKMEzMIBbWVqcNtd9r7ZbFwZ6spZWfw2
vs7yod9GPXo828WAP+PRAImvNZNfi6mRsL0+87TrF07Y36aOpFsTXmXV6N4abTGw
QOQJGS1ncNIJppDZdOv8Q6cJsA1H+YSuRra6l/0JLQAs7eUKsvSiwC+kPJVDQDe1
UfCh7GLs6Ko9aO8L+kKLokfKfw6KGJ/7Le+WGOlLWogYFYfN+Cio9wnErrHg9nVv
k0ChLK9urMZmMcq6rn5fk3d5V18FeA841gpt+BRkMeQNlVV4sHib7y16nM8cYYFf
hHqBUCfhEZfhBf2XGfn8AJwGB82541ZB/qvs/rd4KIjiZ8EMrNwe2Jfbr/wC1IMB
Gk7g2xwRXl30DCueTTCUwOGUsKFddWI9FcjkW5FzPgDBFcTy3ROsVtK7QEGvGu8J
tK0mYxvQ/5ZDLHsNQPk+r51X6xwrZ+rODYpw6wNqVhDqxiGNI0wZ9T2xZhF+4v1z
Fps/KvQArvOZOY+AdQQSLQncgFNh5wyw0m+9fggWqlSGb5k1g3ZRXnyPCN067Xui
UvhwSflgo+FLu/JcyV0Jby8NKUeLxwqdylEdA/mOYBjxMuoTrT9r3xl/3ZZgFyg9
sVH5UdpnGplDxhMgcL307k/KCh9yOap3ZAQeUQ/iM4KtODUPntQoy3sor/L7Zz0M
mfUs7dxsfVDs1eCTpCvPpaxND+pHpacv2YIJwBKhLOUx01wVi53yDVMNR86PM8P/
yzWH1FXqqaX0TY9lOa4vkFsLbyKJr0KqXr5myRXTGryz++jNv6N5mETasSV5IPQT
1dGVC2RskCdyMPxyX9jH1pmedjJGP8oq8H9pskj3E5AmfpOZ3mCNIOaBzNMdLJcs
ULaUilnaCgEtRa3lkibO472k8vT7L4tmidegY5fO7H5iXFxQMrN4Jr2cHW30Qa1c
1L9nyDItYugCOKnXoVo+2HcBv4VJOhOOvtu38z/lsaXBcZyNSAvHQWTAIHTMkYUp
wVzB/X4/aaGPYUSExlocFcS4g42a3faxHzWgleBmmpjmzrPBLJh5ZlXaqaO+UO5S
A9kZBAulULc35iLmGngmJdjourtKpDGaQe3Hd11CkKTwaKpY5eXtY2g7ryjKBUKo
mbMUCv3Z01ecgSFTSYbinhzGQSpzSQmHy+1xCJfwbAckyhSz0ywNZDleJ9SJnuTS
t4bvurq0Gf8zeHByPTGgGeOUfCENbG4zEvxi7V+hCLgcjacSSxZ5VE2+OCYu2qpI
rqYTqtP/sn0JqGe+r3tzLn9BoW92rMyG190cltvJFVrm1txoIF1DF4KzgFL3kCJG
sYH3H4FlEXfvH+/U+bWT18ftwA4QXiXhjAXN8uxCXHOomMKqNWys6gkeiI4CrOE7
T03d2m8MTz/QnA3o+KChch58tggvp6T96jTrUW79vU91lgffcMEv0VCpId+Ms2UP
pbtT0tisJUOSNFI5AuLsOXizTiRCd01GKIE8aIP3FwVztSyHEtr0orq3g6F4/fng
QIC6GDBpklT+30UUkaTZwLSWnTcNHkhZEEWtrn3d7po+hwN4XILjz9eThKI02Aya
/CG0ZwIWYy3XxZY2XGI6KTECnSigkFhfBDtrgpk4wrRxzrkTDNe6e5ixV/DkuAGz
TFUNu8rg9xCEdhAtBwv8gQ+oLVt4tuObfvaYKaHghwtoK6096ovs3OWF8fQ9AsK0
RF2MOa2E7OKH9wOWBCb/TnIUaW+k+/8BaT961Z9rr8DhoBPhnyZxfz+jPnVKVb1/
UtQpgX3u8kSVU2c4YQT9O13lSbTxSRLuBlys5wvVbWrXKqAD7WJIbMoKUO51CqfE
nHNIZgPhHg2KxGfuedXofkSyBIasZLSoPQ0ykDzw/UQ3B/8EBjBYgbciJcPgHvGK
2CF4chOmMOi8xve+K8k5DL8RHsTcq4KITUZ0epzIJnwxugvmNzFIVBtMWRKnPluo
C1tWBspyaJqsEKO7Tc8E5VlB4phavJs0S/EDx7HOyj70Uc/zMyPbq6PaTP09U090
MIDDwNnI/puUO/qLmLNHZVxcUSzD0CP0RD4rkHhPOZsXfLRX8+rk7ofLc0iRQeE7
pP7td75OLyiGwVKsqXUBqEMYEsiYrQKCJhpcDO7WST+N7w5dIuDlmKkLMTws83Pn
WKmLUZ8kQehJrNsJKqKNjiGkzCWdtB9wlC85HggSlJhEkrHba1togC6YHEX/Kc8n
3fqRvv+fZjpFFAJmpmDs0p2mCKiFDpeJY9ZmcPY+nnOoSpOfUREAPtOS45dqjGL4
lrI1blJpI5Lr2Ze19FUWUYSbmW/xPrtZhz9xKM8hf1rvuPeSjoDw+3p+OwsZ1bEv
fMOpI0kFOT2PoSsJySng3bd2uTPGUtuJ9LGZpmGlRYRTS4zvOYDGDNhsIflAWMv/
261n3RGz3r8V13hV9IR4/yCFGedddoMgwz8STJhnDBHc+FKjLoZmz8SPqiupQkZK
U7fT4ZA9YcNzQNYCrHAXR5rZ2zLe2Ni64XT9cA+E6wtwgLF7Y2Q5j4IAchKH7lgh
umb+YsxUhlMHhKjBrGI4/xrIvnelqpuNMi8FTMZkVxtNBT5lusl80GJwFPztl2un
W6YTiUehSmpApO50s2GVnSzLXTAB9qnE5qgq3m8Q4k5DBA7AkIq2yIJzgEgcwOqz
OZtINkRgKb9dNICiU+jRjUA3wEfQ7cjqjyRXu88aehxUL1x81neCjUjwhVc5Lxdh
gIXEusFKzOMWNgYipYuJMFsy+eqqk4IaPQCJv2IkD9oYYzL95jg9zRIWwFLDgqjn
wYPpSbGFJlIi4hdYLxACvtMqxyHKNviEplfaSKMLZsZ0yh4UXNDZK6XoClqtT9Jz
2GW2K4isOhtUG0gqIyVNEaTMdBvLqed0s/S1uM1xp7X0D5iZ7fYXG3GUM/ABw7dE
Cti4RL6O2Kvb3SyHUwdUpBc/D6XoMGMb+l6exebcjobcU5qV30KgLFGI6odnfnFu
7mo9h34kr7b22o5KrtE467sEvQKt4u20QBw2RQuNji62bZTe1KxsMLvUze8deQz0
qlw/a0hnwYbx/r6Nw9D3fTZMWdb6XB09V0Y0M61i3NQT/z28vpiTw3OgRIjDJUaC
S/I/aCqRM+rZiJubvWte/QnQkHeml1QT1E+mFiRP/OtdymkJJZQOQIwkwb1ht5b1
nPQqdkbkYE6Nm8cZ7QeiC9S+8s7b4pMwGiNkDyAKWKa/jv9WJuZkqDn3gVdj6Sau
ExyD6Ya3blRmiopZpHrinZYWIa7Xqa7sJ97NfiRWe+6B+Dd0PHd3HfiqOtGkBgJq
+WtyQrm2oDKY68SNoCjNai0C17Uls0Pj0oCnDUHBXcPzDkP36lyCto5/dG+dTudt
+GKa3dFWT40Ap8nlNPLKWrtksJaoNhmK/Hbu4k1JnBltci5wb3MMjknvCNZijupp
X/XIGY9PkX3lP2wqHAIVYe2s+e0aNyLKXyWqnllRQux8BfTdf7yOUgY7oyvdHPsm
AaTfhF3o9KbFAjGUli+5Cl1k81Q16z5BHGuJsKx0HS2SbPb/1byw2+ionr6sZItx
hdoaXUWA94F1zXzvboMplkIXCT8vadUVsOQZSWZikMSUAzeyng+d4ydGdPA/tRwE
yFYTrjjsjcIDaHE1Jrp5953HQ52xZvtvLvC3vRst/Kz1ZCz67fHRrni2hfdZyMHe
Q5tVv0m6Hj3nMhLiMIFxz4LIiOcv3GiBP6S9zRLc184FvTTTXNxcooQ8UCsE8z96
PpJazwzwLrB3UQbiWqXLdqtlZaBxwsE+F4lauYuakYsCW4E7KwJA95A3KlezOVRL
eBVUDepYIglG91MKiVVAq76MTNMWpVUeswAq0g37625Fa18kjStEhYslH57/afuj
y4nXulw/L8H3yAZMa91tUYwFBTB7+/NlVGZmON10NEYvYBIHkrN48Gi/aJz5h8wL
ed32Gz1Es8yv91wBihK79oy+8yTy0GcxeEGCCBEnHcKt6auw7CXLV/6h7FZctlbc
y51j44RUMZAgJofWJneh5qvfPQTjmjpJc1KPA7962bKdg2zvAklCOOwxY0LKjLEM
iPGcvm2of9Def2Kk9dff3jH7elPYPh9OKHWOlZq7Z4uMMmqlaVdV4+9lrSNvRsGD
WLZ48HvennhnLTQMWoqDsZnSK+5KeiAwzFGL9hwZIx6uCRT8TL5LosQf160GwaW9
s+kAjRtqtvkpzbC3X6++E+hH5ZqS6qj5sO891o5M/SmRsfgOfZ+UOPwZAoOUVNJt
dZyni+cU+6vIbJfWSnYbk5Za7TlTSPgThJiySwSn8QijYx00pUojVXPnWn0emSnd
H3TwVU+vT3dgQ2dNwrPTTYAGWX9RzOhMgGoojqQskdy1hy6HYQK6c7QDiQJUTAqY
hgWAL5RVMocHNjzEbgX8lty43N94+nS8SlHn936KV5MJpcmJi+S3MYINM46/CfIt
KqkW8SoJ5FkgMEFEC/VG6C92lEEKfRwNbWgZQDJ9ttMHvUF8BIRgv6oSRi7RlwS9
alc+c1+4gPY7FiKF9Vbh64V7XEnYkOwJnrRYCsCl+ENO62Y7zuNsfT6kMLgWrnXc
vt95fcW1zDjxVnbSGsd9+D/WuvtPHugMw7SIkkXHu4WJcMHf7K5SUg4POzmQE+aX
r6ixwPGFdzg8uV2yOPmL7WcR/A3BlhhGFtCUz3YSb6EMD2lXGfV4Wf47S4YHMWKl
lQKRC3kxEKrUIri13Yp5ugZmUlGJUaC0VQrMuxc3yA8VBF3oMQRsarHmOTZy1Kfy
38Mx/YESuNMyXYiPB1HXozxSdlYlWyeEt7eQKvXGRdAp+NUiZ/aD35B0IfdTack+
MuLcGnk40jEA5ZyFXKr0l+kgNFDTSjGXhFBYm+tnOGvqUkdmVhTlmJkkH3YLa+rm
lhqcdvOQeazLf+XAluGIVNyrXtoef1DKqUxUXOegr0CtPRqeoG+6z/32oPtAz1z9
FrET/Wgu2oR9b1nsIvHMqfnFlp+PZ2B8Vun2MF6Ksl0VYiAyN5B0lW3znzBIaH7O
A4KLkTu0LwsEvfeYYzTChwJtaE1+FUzWltRfudnfpC3iNDWxDWWJK/D1lk0naoUM
cVq9zJZoLF0OKRx26EevADgCH1KPoavD31R3sJkaJT098jy/lkvqwuCcH5+Kyu5j
D75Zy+uUAyRU4dNyoPE0AWNAJsuzElS5wbBnCPMCg+9zqMG5FTGkhi6H1iqQ79dJ
/vkWBq+0E1YXP3zN2BUl/4fAb8mDoEDO2qnjYy7sQw2F7ONUiZv43haZrHXHtkdM
maOk16IhHcj7QmzjMBDNRwMIwRKUIzkMt7ymY5Ybg+si7znDDJaqmloGvB6uIX+h
kFeqm+8sLSovdZDjpTqzVV1AJEmJFCoDxBAXd6235ukDcpS38wO17krqWwk3AYui
OVa4/vXdnfdPo+kXBVKFfeaDLH9FmmYxLL0ebMmF7L6QE3jVmQRVWE3dt+RYhuzH
dJFaYX5M6pbYeUcYZuiFqouQ2m0WCWh1YvuAHozREvvxYNJG/tSzyK4KDI1JuW4Q
zzCaipaSKSkVyNsfhzwvqjMl3aBLYN2JLw3pgdAObM7jNnUD6hEbrRee+x3vFxy3
PnPdUW+X5jf1BKSOhnyLd4FDhdBnYHjEh3ylsHe81kiNV3k00eMcNrI5QTkn7R7B
jS/k5tBXxq+OsQAvdegS+vC6SipNp6+78QoSnHb1ztGYbp5DNMloNSmwOdwsZDZl
vOhhuxIQbpYFXGDpa6S6FP0iqEgiUIPjmpxuiODtlF8CIEJLH0ZSF2RkV7XCfdw3
2bZmaGgEdb992aYNViB6R0kY8NaOnn/D4oyi+wsRz+9deR0UT/Uw9Gzx/ScX4EWJ
xUuaZb4X7N3+Y3HwtFcQLKukaBJco0/iISmNeTLOriF+jDx6cROACY7nI2SMDiTd
uHKiW1ujW8ocRVoOImy/p1Rz+XSiA1X6FzRemNn5IN2eE/XUrXmp8iBro32YGEIC
bC7BH86PeuU9m9Ms5A7X10WSBKNuh2Nve8G2NENj0HgSYsTokXlZsY+dTld+9uVM
MbAdppVJhP72yCpcgfvE7GJzhQKglWGrfk3eeOEuejlIVyOJVZZAhWIkw61VT31Z
NNezk7Haz2EOcTxBliGuOsls8R2Hfq0o0dFcGAxZkx2sQVpCrCcfli8XDJHy2iNz
o433ykFvzFCx2lCPJtjDNvmY4zzpT2pwBsxDCcBaaChrhVgSxQ5fzFRB+4Tvz8Bn
UApyGYbLM4zlgXMNOpx9B/L/Qfmh1+V5j3chMjRI4C41dd8pKusrzak66FxWIcE1
R2VHCwVZdq9QUMluWdtpA1esRFVNx2lNw2bT/LI6DkCvljYqK7+F+vGwAtDGDzoa
m9UViwneRjC/CLm5JwQ1IxLPXDtHuGNdFmas3jdxTSkXHKEg4bQ+pGl7d6ePwJsI
8xGvpDpnLpcOf4IQwy28XVFY9OBUi9OcTtoBUM6idEXohRVpfR0mGfuIlFQyb80C
rQ1AQD5riWBg+cSQq7SvrQ3Ra5Bkfu84k67wnCmSIfYRKlr2NK5lHNYXPAKs2yJL
OccU06/Ho5pFO1KOwQ2+C6vcTnUYwDZzohz6xFQE5SgHsF5KJOu2U8yZFHP/cCTo
5GighyVlCN7cNg5RQx0H7Zzd/qz85M26E+92k0izJwN5Uv8FHVl4q+/AXUk+J1Qf
+KD4ahAvYuafcH85xsVAz9/BB7CkG0ufbPBvD0B9I1UNIPTXmyGesfWwEjQjOMAi
pq6GOnuIC2MhaGQT8cmnBrbw8k3GIH/znge34QP88WO/c4aHczv0Vq+xpUXHNAlv
e8nplVoIjER1BhQKLlJnWDFyuz+bEPearVTflRHMry4DRHTMU5XJX1PVjUcwq/3l
7pE2ZQWoV1PbcwN2YiD9SvAyx8EfNw5slfnL2ZIXta5ggMdiRuu1qen2KSNskC0u
UNF3uMQkq5HILiB9DjbAvOeZf3ZhfQvauhbT4Y2gDhSFg7KRT/c+IULGijErpouO
SsyTMOwzQ5ghqIpbiPYmlCl26PYRWxyl+2YPlWMAHDBrvAw7wZhKa0+fMAWT26Nx
8LvIiL2/Wnx2bd2hYpqFZmjTq6oXN1VUEY50EfHBDB3182EAv5iEP06wmuNBNX/t
DDWlRWb/ir2eCKuE6N6vYsvSpdx6V/mSwDEuHj6q5FBjkcaZOacw5hv7jejEoHov
mNnY+vNjUsMkj0cJO887tM6KOuxk+pXhqF+BwgWTTXIFeZf7yi0ZraBXQioh0Rkz
f6F7igezApLUeEtzQWLMYvr24Ss9zkarPYuoFTWAheK0ShzjjMiroVLFL1o0QFNg
dQyVC2aweDdrn3vDM5WlUyDRSm7DZEkVDleDkdqL93VW83SonL0XnRsB4WTRC1ld
vKe4Y9UpeZwxWM4tOEK2frzfiLij1AjQGKmbA3R4ot2C/vmkrv8kotOPZvKOt//j
f28M/Ds/INBB87Oi5gYAmDeKFGeu+iThvtu25x7GbDQrQYtMmBZvWBYYqCeM+jh9
8gfLoOpg5l/Yk1Jvq0LqVTCjyS3YWhyAi2sT3Pu3q2SkQVshJsc91iAAILboMtyP
FtvcFVal3VuSmepu7AhKXJUN0V1TaGWTRxVbQR+eNMhJhqnxyX3KNn3thu8OyUaA
v7vPjeUMkzO1Q4pWAUZu3dd6rqWT5Nbc3yEnyKx4BFiD2gczmu/uoLvadBaKLLDX
W95yKakFB2AkV1x1vAzanqpZzoGaWcFETr9QLFYRDzzfq8JRJRtkEamUbYPSbQ7X
DxkffBLQOB9SbBKyRxbHMQj6bh6dinPnV36rnu4xyV3lCrF+MgYx/ercenqac+Lt
I2To63wBPS/6CXkFKuhBhfk4JCUqao26NgbS4heNyi0ScG7abuhu0irvy1qi34hH
TRVnD+o2VImyR0KCWUQt9tmwiXgXu8Pj1jy7ioZRjR7crnHmDnt1BqMr52HRpHGW
5GmN7ls7fSGT5aT4MgijuQSE9rJjcji3ZWyBF1ub1b9RW1/Z0HCcKz3S9wIBRP8A
binD63VvRHvAJ4vUjVH0+OGV9N2hlkx51TgbfW/6O/9WRcCg7izvAXfE7NFlvS4T
QKACcmtUyE26hT5ENfMJLfFvtA8XLQ4qhFKfkHZVOsfy4bFTSBwl84JRSbARh8Hw
gK7zEG3rOhlcpP3g+RNJVWuoGhXThUCeAEpXViteZyQbE9xfaI5Nfzci7z4l3Gy8
YmNTqrmEmRXzFE9kcWA+Nc1eNWmtbZcpzntxXObnyO0AbG7ChdhQBNqJWsXG1RwT
ADizZzTzX6wGE+A9TcuS06rsYxYXcaLvSj8pXj/roAEk35VS6EocHE7wHhAaabpV
5KIbQdMwLYv4/ZrGo1oBYXCd9sVJptPjkn2qrqYSAHQJUuv/eTspM7leGzXZqxYC
raXW/PNQ4zMUZfq1ImDmFERe60Tj6v/utt2NboFg+8OZ3e7/gw4g5nevsb0bboNT
a+tP8a+2H4fqR2MgNVul8Qu14FyvUJ8v6OyIAv8TGgjGtNILmOnSW7v6rX9rQvX4
4Wb4ShJl9b0xDTVIC7P7Sl4px9pXuddPWtjD9G+zwjpFLhjeGzUpxrqMzqcuDrmO
NnsDR770zPjRk/s3bI5TjH9V7wwuhXbZ3xGJe3vl1QgVQEgb8koxbi3gQB9NJMXK
jOvbNJvrK7ZF8JKMc7gQiWT+M0BEmnNvJfPcQ9fX0hik9OS/uvPitvUdHj/7rHZ4
WecT5CUuaFFU+8j0u32sIQcMr2g1ss64iwRH6aHoEPbpkYqXz49rmp/GSZ2ttwo7
3igaTLVTPcXlI+VYtdezNy2dCMDQer9AY39bVKn4e7rGlXwdTvgxMzgM/fu3cv7v
j8o7IUaM0AqfqmEFZS5HKU/o4qChtzNOEburEUrjprStO70th8sOZhHRbXBcqZG/
LzEkqfWxMPAx54URMGw/UrLkwKoh/csh7idlNA74g5iE5wGM8ECD0myMI83atOqo
W5Y5jSCBSyKjT9fy2arDLtViBl0HmCLqB38lYAVHrYAtYQHqc6pD+6//DIeFzO69
Vycq9A7iF2DFoeQtHRQFaXPKJSJqlRjICxZLT+OFma4AqpNafSuFSz5tjRAYMMWO
JL9+1e3hdDtg2jEd/zun9e1PmDxPWN8iIZjrU6DoPKP8NGPHvLrpx49PcYR3Vc8v
NRBeU7z22yDWDKE9HCgjlrxFE4zBTYQniqzxntgxJAct5doMWoDMt/D0xTcpzInZ
jXOeIf9PwSPKoddfTzbOBJTjJ7/RjIJgcT6FUj1p8pbQV7B/4ucgiNXLOuYrot+K
5pQflwBVgvzAARHQuPKFiDVHDEG1JK0DXlWAnj1Tsa4IgTAZprvABUt7/uaFaZyJ
UdsySkkQH87EBP43Lvtqdh4qfczdquUqhjAcuAVun5oFMS+RTeoQHj4J3qh4sFNU
qVEn/aKE6uz6NKWE/4x8tgApk2gu6QRNzwnZkOrjdGrE5ilFAdX5RZTE0QDTL54C
3Dv8C47g557ieWrz1DODkmfTaK3yqO5BJ1GiiLOYoOdd72KiGiDuCGz1jKD7hROL
VS3Wdxpl9GRlAb6w5Ye8enGLNq0SBpZ45KK8n5hG8/I36jCDjO4W67u7mEvG4BK7
yFBOr/V5BladbIOq7p+txmq0gRjDRfjSHMn5lz5eit16V27ePkvu+H6q7N+kSyfv
L1UIvrwY8gfqn9qG7uz6vNyoDogx22iL/jaOviTm7purnHWgR9qmbQVMOtq1vxkI
6DDN6UGATlYTVTCyL40QUwToFm28we/88vfRL1rwWrR0kcJlWeyeO0XNUucEqMjt
JPgWtfcXI2wnw/vhdF3c/coEYt46baSdH0DcMCAZ2bx4q+AwS3qk/NJdIDHwOH7q
cplJD5sS38Lb851H3vM5h3LBfBnYOZPVK7D9JMeDraIABYUtAPX6ErrwNfIVqSQo
ap77XgLQGbshC9XHs0CBjWgbTRcBS9/SKZJyHNVWU8v4ov27JQEkm8exnjM9duvT
V4Ge6f2rAtaYJ3/kzlimKpg7p0GWL0QsBQ+6WeghSWNdoFJ7lZoYANrS2jMrHxBA
2BY4DtVeV4z6f3NBBx+SnEMUDRkr2tlD8+ohVpLE9DT040yrtNqfvYBO0fwyqivj
dd2LKAXhX0mODO3hzWou4h2ge6Ei7+csTbeotH5QDYrhOc62ljAq4YCccljb0MSs
wboGCfm31PcsbVuldadcb09fQYnSuBi51u/gvlInOc6vyu1EZ1ATBvnghLp4z+52
wqZ+IJncJsCQYIdxh1HbXTdXoWILpqwG/m6FTP9cTrQ+bdvWUTTGBd9MbJVVAP2N
RJDLIoR927SBOPZobfsoN2DYlnMt98aiK4XTs0lVCP7/5Vxkt7pFpes/dV27lZ5q
hVzY31ZVVIf6HOJZBvrpNN83czY6r4hs1URdGHNAF8Oa2c+ExI7TlvJFd9wCKc0H
9VNpVGCG4kEvIHzR/QcPCYOrLrmqejrpZbjM+oioKMYMppcwkuFzjkQzQClZb9t4
SChKlwDzGJ5mRc7uSeGKKCmOi+PUJJNOPyfjUIDci2RNNo7zQTZf4D6w2b6FIWSd
NlY+Ts0o0THGli781dRBiJ2nQTDSM2p4wSBKLJRXEckQyZjn1TI+oa/rO5TjaCgf
j2ojfx+hhOj2+0awb2g6/jRnKfvajQ3NamMKdrh7jb24WZA57+aEfx/etneOwds8
CHCcUPj3R3X9/Yoq9WHi9McQ05K8AtSa6x5CYCosBMt3GwnVn9iFuW15Ik/saYx6
rOW4hHELaSDKJeQSEk4dSjIZIiJZ6axCYLBvqESUoPf40j/KuCW99b/XLLDaQKbm
9Z/WFQlnAez6hYwgdgzqEH40izY9o6Y28ZucU3rhdVmHAmpGGqEAkJi0laxlFm9S
NYrXj0xTEq7i5/I2k5F2x0NFVgC+8jI6+dYy9T8rxKFwcsnLqLXHPQXahhUVQKsM
QCANEwN6y2ZseWTqWYY51gTIVVAFo+oMkVFfXU8YFBwrz5MuT+dFRcCtPDim02wb
PqsklrvaX28OM2/iLhFJxFfL7fSVu2E1gvXq71lpt2VRcAEZ/16UepT+4M1u4Ogd
JB9PRB+nhLWU49Ie4GDMr2l9lhSsPAgpI1QBJa7PkrwUblGXXHf89ZU7VQV77+7X
MHFqkh8LI7j/s/Rjby+zJuvU7NLs2VpZ5wSmtG6+GyMMKi/9/8EM8qV585bUSOG7
KRQcxz2smlN7+4kuOPJ3TIo+JNm8M+bd2aR0Op4UrFHk8Z82Z06V7TvMJtPVTwzS
bVxSl4Mh/qf/L9kbRh869WQRGzjOuoB/jMUSOMxAPN1MOlZTRKIn1BKcfHTHwsXT
v6inRGRwU5YqmXk5OfnuksuLL4K43pivHZGI52wekuLiF+90MRTaiWNYVpOCTRm6
QotgyALxHBd86mtoFhf50cr4KufB0Dm46wnxbiLNNYa0PNy1DEuzUiiezq4D8HkK
TUAcJHTPOqrC9LsuBFkhb0YoYxVnttd1rHYZv8equscRpmitVvYL3JqKjQ5YvHjA
BlewGbTbOCXIf3cV3TZc0YKLLVaVzMMfH6GXTToIieMLEvggIvLh/xtZonlCQmZR
0fUxzc314oESeaVTGqNboU8kkCvQSmd2NhUactamnMkXC+7XVgwDwMyHNy2Xpm/U
Ez5r+SNf16KMlWtg3DUejK0Ln1ne4g58EjcxVzqqU3gr/LRoPzYult1fy+6PabSK
hXjydaTz7sPJAgZQzPnbOqx/YfC9u4C0yA0X51/bQvDUHJ6XmPeCS8WvUT+/8eLg
OgRRYneJJs7kiZ/tKxgIFR24l3r2+ZHdgUqnz3OROedVUUJiGeLk4Hrb3mpNHTFB
vCgIdRj8SwiSMrSRUyE/MG3izlCvIgGli3K3DuCrBDjCFRuxI9xbsVRYJkbpL4co
dmqmlApkFfQSCRpfgnyhMnMr+0wTzoKu71wHPqdm/RTrTA526ffZIpBpPq8uphNs
42ksWT6kctVEOyU9VYK7NMjB4v5i3pHUvDyhXMlk2aZOjjPBQOjeNbkLunBsXxDa
0warfdVT9e0sz47FZOx0zALimjOp+oy4vEcb+nh7bPMhAlAFGGIHL4SalnYWzTMi
/1b0iTfdf8GGFaQcc92J0/wTWBOHr2ZGEEuE606WLWhpcG5yppSGFh4qHW5MMQQf
9EuU13c5pz4mzf9eOm+m18AJffXGJOHV8OrBReS0N3NazfblNHeSBpPhx5pQSWr2
Kj+6zhBR9YQpjQEwkyrTy6TEA8pMs5lvZJklxdpdJCZ2ICldeAP2Ewt2fgpWF5WP
mWmWBJOPCGrl4lSxQA1jBIQCInGBgl5O6FLeGC2vkonQkuJ5sSgo3zro9hBjpXcd
2VksG/Fcd8jY6OCVRo6cS+Svl05xozhJkcKtFBxPptKKNol5mQp06AJLqDxQLTwA
Md1kt9/X179T918TpNYEIAqqQCtCxmUCN23GqSCM+aU/f6/Ei2sJER5kMJrhFv5M
mUuv/jvtTpH5l9i1fHHxopl58jD7iMfHt0Q1sK2z16X0Cb2eXR42IW7m5i6h4bBh
Dx38ZKt7f2cUdpQGZhLkaenCEMdHiZXC04eg/OeG+xi+8axDZzMxQSlf/ab2M+k2
WJciSoaO9Ig1uXvqSjis8g4qfyKpZOA4sa1Pvj00CUtyJyU5QQ7fgHJMiiq3wRC8
S0CGdjHRYVh2lI0Bz87n/VFbZVYIY+D58vjVTlBPHlnOZtaY+tfkXwduvBBNKaWc
MLGK1NIqE25tKBb/l085y4rLMYM7w6gHmzXd5ToMxdYFomXOpaJAeUrIa3b4XlJX
PaWONDSiXcDlR0aitB5RChgfA+r0/bIf/RmmMVmUEITr9ydTtWjaksCDuaj2Wi4K
QW9cSqjBEdHBz7D4P6YNiTM7OETfq30FgydWwjt/l3BY3cdw3jNsDO5cMNytkHJh
S8tvbqdpIQFG6utyJXGSY27LrUUbYKmsL1hvHqIc/W/tUOieOx9zSdkqwdh1Xelo
Kwvzvdn8EHc+9iQ5k5IBR/kReH+L+dJGBkCyyHdEIQ/n9sSdBAF5Nw6YzOZZZ5kl
K4Ym6lg4KwNXCx+naNjbzRLXWznAN0+UORBDskOGamLRkLvAfS0uf7UmThbUlKzy
J7Oa7l5ljuAQsznLvFHG1sxkU1FCoQxZtK/kUKwOplhZk5humSf5ICQEmp5yXsB1
Hk3oeGWbehVsXFpgc43twYm7TT4RpX7lqQwd8Ez7sM6z2kixsDzcbi1Pagfo9HoC
icbspWt6BfNEj4unbssw6MtXciuVLrw/tAqmq1uGie4YhtMZ6wYzSRSgaJlDddEz
b7LCFmLLHDRQ07puI1epzzLUxWdjB+u0moASA6t88ETX1N3ydISpN1g8it6nbrAP
TY/LZd5x3iLDLLVeBd0qoeJhE2VkzeaWxM0QSKzRc/Tjhsns/soUFqGHtau/kWi/
yRrUSaY4CFljMmQ6Jiri4RA1VMp6ZTb/whOBSUp1Qh1Q7QlEOuFSNcC/2KdZqela
3abWB6ZZEnjOtWMD7JopxtF0uBiTD1n/+jQ3lPQUxWR1TRagb+p3j9n3XlQuXUje
cPEeKnOIMc9qBIIf5jEb90kp69dZxIHMpN4DiwyJJ5ZFjTxuFKrh1AWnqoQbS3MR
Rsuna/FNd+eTnw3qIsSPhxx4OM4neUfUMXlU51foXeSDnKgl5GSsZ1KcMwPwg7/z
YZdvzueTRat6Q3oK0O/T35iV6P7Ni6ijfCPLmRL/cZ/c4JxMje9ZoisM3sG6dVko
iVN4hjYq9+aSmQLaIXfXvYWMRZMQdyfj5ndqxlDczmPTpdX20Ub0mIDLUQGqdnbn
HIVrw3xkevMVFOW7WX7gtIbbnFjzpdBXh3rl5kdiMVlJYrEUSXY2hO7Vq04SBQ2O
a1hWV00j6wNyFV2OxAXZCJdFstHKX6jrSPlaLiilZfd6JrUZ78c1QcQQvErqMDn4
iK9x3zsL2gQ24n8Jl0pT+Mx10XuaMij+uP2y6XW/1Yv0e3mrNrC9BnnJ9NJr6NXw
s5it3eGWzXsmjGWxzaozQYgrYW//IaPzi8Vt30FxyqKe73kk1ou5WtXKerW3yDfe
3QNMSywmqZ37s9mwz4UOY4nG0BMCx1iQVjUiDhAVS2mYoHLor3g8hA565kuCEe65
SQmNg1Fmiob1pcSutZvzs4IUa+3zf4ctRgEeCTT4spiEwPg68F8KxAfk8wB17dft
4Tv5Wmg+0WimYya/3IZJW19kjagKVn7D1sUsSxP2Jtez4ndOM+72OWomcsdkBdcG
gm2qcRycqniGx3TlJXjOC0pxzCKmkl67JxjtG0hjQUXu5JuZKFEQhAZEM8jB36Zm
qjQzxyfLkxCyGZeG8WK9f2bJlvdmadss3cELFxm1Flh+SKD0WaNXelffgu4vbAsh
Kif68qz5H/MfADeS8RGxehpkOsu1jxA8xhg+ZG2dUBfFg6JoBXfgQ1dSUhm5pdmy
/ribjplhzaa1Ham7FrzAttpYqznVtiChOa/1OoNeGJBF1dTvqNZ5aQ0WLVLRODPe
XAOwNQ8Vx0rftFpkzlz4Mfw/8FZnoy8QUKs2KkwniIpRFZzrT8YC/TGyn2A4y7HP
4hICjIk+Sxo2sX0QXHOKw2FqIhgnGUVdTony9uNruDtUYk/+8P/vD1YFDm0vFRSu
e7ZCT0Z/Udo1KQKt0dF7MNjCKEsE1Ijy3NIQp55X9cigmdCLbkenZDuexJGQTUaN
K/F39HE/N8xdM7hBu9HbeIv6wjuuk/10h2W/8836wTWureEUtWOa8L4mYPRvlUOg
WmZAHFWmClS+XC0pIWEw0dK+nH0zyUsUG+7kXBEpaF7wUFbRfu+kVPu4X7hjtIsd
ezLwZM7DW6jkw0oyluLRoKpBBIkIXHBlBzAgPK5lpsywnclyTnEy7DIsR2FlVPI9
+OPJJP8vVMKZxLi2VWSoWuJQqyv10U48e7ky69+jdb5zWX+vWEmAn6klv5oesb10
D1pgwkPEH40Vewa6LSF+X6TOghuEiEaDo53j2is1DVnLWiaxuCATdOGLgu1Yhfgu
0FP0g3NJOeF/kyny5gtkS+qXY8xCmF1YNXdrbgKq4sLSg1UezBANZKJciCbnbEDS
Eh66NgTs3Q0yEYjyqt9qWCSG9W4clV2qfttnynrTE2CqQ7NQCLSxQ3gzz4PaBmTs
e1WivBS4X74KxSSWwRjmaRCCxxMFJd68OPAYL6jL2Sx/HnJ6Fz0z0Fl3RI+T5mzu
ZsKrBj1u8F2f9cPQv5LpbpU37LmBbKZF0CzATO8WaI8M5sHL7+N2pwYbNniQOJdP
5vlI3whZ0b/B5CUAUcMqevKnrkUTBF8pj9ZtlQUutQlNG6MRLwwTXSM+9zi0KgjV
zAo9Edpv4NSaoQ2oWXt9QKGvdALuQ4KnCJuqkKac6RTqvoed05PIdCCzy0OUFqfb
zmHNxK/mMIPGYDTg94zdqZR1Dm9BboKVfRMu0BGU8kZQ2kZSr2fbQULI8Cu8etSU
AfwNkglO8wW2EWI00xT9FmR4moF1PedrpNcH0EH6P+SnT0VkrqDS0yz7epFAzfBT
w5QXfqAMEGH012mLmwrGG8H+Zqaz061OYyGK6AWseU7lrleN0QtQgR6x+4Q2D96m
ohNyC5DFDuMCJkAWUlxvx0MqVCuQfopt2h2FUu3TDI9kSDMgBrEooyfjZxqkVpuq
0t9fSqMeiyF+j1QMOSmcR+dvg9ROcbq7ouq7U/WihO9IMT5qfyAk9v/d/eSf8ouu
D3Je7FeuUQ1IIwMV5pfDEhbWhdHDJ/Jj1R3QqM+I2WOadtmEeJUsvYrtBshv/kpX
rfqEobW/d1YrdOJmSGbl95UPQRHS3WmFGVBPMv/uRiu6UZ0/B9shYCpyosLaT1bu
AKpsUB6HRQH04bp+YnWAwr5yzXf5sVUEbj3DWeftwApyrIK7WRSasRG3aUbj7URq
pvzFiNR062taIzkS5UvhwYMhZpLKsTOzI9AwU2rHr6uqQTMIip+I5O8W7sEKsUoJ
wwgPcqEUkQlIJurroLsshUsjlq1VSO/lNiqgAN5ChCvFh/AGL4jAXxFHACmKWExd
uIH3T5+l+LglOXxrrAFe5T6pFn0JUKpze/MRMs50GnwYNCRD0VsJDxVEKvuLiXd+
DQCvdSmaMwfNPtZxd1ET5LenO1G+TC8hJIdTg9IEzjPyXl04ozB7GN/v4ctE4AzV
t4UsbG25oMfomAzZlY0xS0qjDwPeAaOvP9ob6MI9A8G4fa22AMhpECTBOdrR7N6c
dV42Ha4h6N6jfS9fk/KcxhwQ1eLcIxIk4VU3seZEd7GJX36EMLPEOaT0jQvoMBJB
Kh1nNvB1FwfdY7eMx5tvxYrJw9jdKuZ9TRXRBri5YltOnEGY39wBokMezVg/NHAo
rrKKQDBa/NzX1fzVjIRW9Gg9QO3XXs53SFfl+pE2IHROLk5AQV6lJK1NWhuRNjck
k8IDJKFLT/fOBv9rYDf9ZXMqyfl2tIwdJs5KOrjoUzaGZvQcWdYhtdSJOBHhmeNh
nNGh3e5J/e5GOkxreOdQ0MXuBCWIk9cpVo0CIG9yBZGzlXB+RFU/eMuewR1GOQwg
B2yhrQA4WEF48AzudrOHcqVshLATmi3b1crug5lUf1BPqM8T07/Dq3zR50zGe630
fOLXzwve0NFs03mtKHOub/KE2n5a7CJLhZHG1qz1WrcFt82ZZZ49jptGCDELb8yu
8PmHZs/fq8bs0anX+xOM1R4Iq3t7fHET6zxcPIA1BU4Fq44n9aQ264LfxtaNIcen
qMbwf7jLdssbFY6qcNiypdf7g5l+nizL2uerYTM5RhwsVMkJWytinDCYOD/FNApq
EvCRxdoq4GCFLTmf0HrrkHcdLhut79ReA6TD2Ut8L3JP0zuclctEdi/YETAsdPna
KQg5ved75Mu7szUDOqUEe2ac97mObz9KkVs+5bcwyEvhIyVjrgllPAQ3VNDXo1Vp
QcYHFK59FRVLYbnDqa+Yij+RAqqqiIzI+Yr88/RzJE/0J61U3tjKHac3yndBM+IZ
pUttkNUY2GieX3Jd6izZP+0GKUhz3DJdMHsXvI3aIX1/hyH0tj4BeoDvxgG2L2bA
SjVIoiD/VNzKmhprhZxMwzeOSd3C3NJjH9q8EoMS8f+n3Zs8HltKpe1XJRsjPXxc
CAPhYtbCur+X/VfVOsi5UMF1omcXAcyLdpu773ss0sOSnzya77nY72BGU2B8bJzY
1hvWxPrQbVvr7p0baSVJfM/ZTZjj/xDR8ZPSLkRlV2Yb/ccTqpVAa760Z5rGwA9O
GGdb1Y5lnKbHsOXOW4V84khvThIaKm/gX/05NtCMTVOKqtVtYiOkNkAYpKzf/5wG
R+NV0trEcLfUim8NKc8whBcWmPvBaSSuRqrVSvtKPVorniG3niJ2OTWlQF/QI1Zd
n10zuPxiJ8GV7f6DMv8T47GXOHGSYs8HgaYUgUzmVeCds/rUpdCK4fSsT8XmXaLW
LblA6kKkWERuST+3J3VKa1re6IRI9qJfFioBVmL1i6MWwWoI6KV8+6rxet0IWyi6
Z2/6ey3Gyv0pnikwGfjGh2RgAhIHc04lH2cLViLoFgf5J1dbn237nfuMcCgvVa/Y
cHJktGbJat4PIf6a2K2xNVVnf0WGMjPbYXy/RJM1H1Mmw7pSkvp/kbZMBBGDXh85
TtW8mbF1HCULn5v6R678Gi5e42+hqVqABoA3DZKHAHa/skHwlfUy2na2RDn9gN7y
wUemGogWnmfbLqIxJH+2y7aB12T12ckTHK7cVujnBwjNt9CeHm51X8tvsJ86BCrK
bumpNj8IdAxqMGREOguMclKH4q5R+XTgvLXJpd0ZcgxruFp5wEE03dJhUGHsXPFD
KR3eH/8GfPGJlDhU2J7YJWP9gJIbajG703Ct3F6agSYTMDRBde+piHuEvqORx8cj
gNp4KemEveM/iyeMyiFlPx7cGUA6R2ovV3jkNboNCr3TGMw1sL4u+ficZZq7g68l
gkpXKnw/3vGgjs3iNNlbUZJqOmwX5wzdRQY+KpmBJCB1nRdzuJZWjUk79gOqifiW
roBQkML2d70GWAgxtN6pHbNUTrfqHfAb11zxSNHreAvA8xDehE8ZTHTayLe9ZhD1
ziQwL+hZ9d4akgtsiz5hbJoTCg1n5CRP6gQsLMkGLopfXzaMOCE6L/rJ/j2yml6d
JnaQCxNF1DaYWnhjYpKzX2bXnuisoNvxlz9QzF3TrGFAC/lvOwqH1cFXAYh3tHn+
crD4Vbtrf9a5EG6O4SGPa+SYNcJ7CVm+AF78fWexMY5L7T28w8fiuGFjlzGENxFq
3wKZtLSRzuyIodzmY7rEufQdYNnUnknZvy0egD+FqNTllS8QUYpL/e8kJJC7ZLkq
zPeeJDJujN37NlhTdfkzljO/1D5wOJlXPY3bvReLqvLw2MAThTUrLirw5wKGYha/
fi7ia3g2cBmt3tHI/yCBsi35/qxKVbo0wtlhQQvEzz1yXGl+FLjdw3R8euwPbZWm
NFlP/3IFMQlqAGcWUY5K10GVFVbTMdDX2Z2kD3Dy/KzOEYHuk9Qa0GiySoPFL00O
P13d0jTixLG/9qDwZgWP5HwmHxZW21Rtqk3YR91J3VbwkfDXyBh9wYAX766sPvbu
6vPvimqEojysRkMX9T2/ZaNBlyqw69XBjIOtpH2+M4wmWZ0Bg41fBqGgO4+J79MU
hMjTCJEbUlHGIJp3gBHqZjTDQqCb/GLI6UdW5BWIZhVWqxMpXI0gD3ZoqtV+VN96
1gVG9Y0UslvvSlJBurL1Z2hf6SWtY5FluI5AdAkaWNyewGUmemHxMVI+YK/esT+n
H826Tk9eCJFxIBcXeEzv5dml1OHaawrwy5PX4xP9YMevCKykqUfnPt4C8O58Q8dc
ZS/uqDurRKwBWd7dk7QzmHurc/Th6slbOLcQ6hC3ju+R+WA9mXFmUutyimErcZdw
2Ty3VFIrs6tPxGkTCtxQVeCjStEPtJE2Y+VIzHus68nb4dUBf4/mhWGdHsOcHxSx
YVakP8pw6fLrneaj7M9lutUbq3QBdBVR5ifMMcgY1BZ0o6YT+vXyn9VFepzT3ut4
+xDueDNfmjq3850fvZjUpwhWRxDAS3Kx6R4/gXVGz14HR2WFhgHou20T2Q4yWJI/
tU3QYQJI8BzQV3Okiw7nkwV0O8NZces+6xX/sbMAAMSRbNlpvzlLgbz4ZxZ1Jg87
GGzBdZ33h8NA+OAT5DF+vu8rX1i2XBzbX1zOor9UwBNrd3DsmD7NhvK1G+6AyVP+
VtubRJfoNFNYJfHEsPmdUueXLnVqbPIR1fdF4qG270fDd5yt5eNGcU7cxYaXD1pM
4VQovlL7QGLDJVQyifO2XHU7tF37LBjMbk2XhfxlfFSNV5+akKvbn7l0+WXWQBm/
BPLzcP1piDugbqCOI+yKLZeyoCA1Su1IMqWystVwZoiIpMp0GgKnTVQ0Nb5utywH
nLYEeHjHpcGw7seectyFiepK3fEnrDjGvcMapBMyMqqiFerlygClQNovka3Uoj40
Mp6SYwjJ/h0rrYGD3OrgmqMwMZmExtlTdDkXswJSSFHKFFZMJ2qOyZ4d8akZny3V
TOHiFHC972hJA27QN/hFqBwkOEy8Q0Wn/sdOARn4F8AtEq2mRjzsr7PZ38NcTb+f
BFL0c2piaeBUeIBGNmAkjhV0TwR1CTBtUS0Bmo2Xm6ffQF6939kpVDwcLXrgIfyK
2W1CDDvuPVQfhec9EurzXwOVrYcdMkLHJU0OcM7mkRPOw5tQlIH70MLkeXf456My
bmhJC/G+NHwR22lt/cCzPmVadbElDA1QvLmy+29OLtAeZNdI482HoN/K2hDByyxp
R7p76HAEl0wdhuhthZgmEHxTkepUFV26ZwkvJKg2LSO+P+QuJD12J11+KgOoVjAF
+IYOWlKa8dKxdgsCH6tNL3wle1g5kIymjqR+HorCKU3OVOTGwwh0ZDRhrxfufMtb
VOy44vwMOnu+NNyzL+XOsBdRCLh5MeZUtMlYAiLynmOyFAVNia9qnjG1n52llEkk
5/cWWnuFC8gM6+yotIlzp6IgP5z0vdCcIwWoZOOFW82M+c2RFpTZrgcbqObCuZVZ
Xq0iuKoHOYnItY6WIHNKQnZid8/UG2zixIHe/yNlVIFnJCMCGNFEj4W+aQVEXy+T
ukWcGX9wRWqsBHIbPHxdsZ8/e4//+D5BCLB0OwlX+0ofuSNny6sFGvboEhHoBsYw
AmGRCzf27v1Avp09sWlPOzFOgROLMHsU2mtabFqN2U3jo/2cpAZ7g/xsiOa4uOKf
vTSrdRhq1fZrCjDvwOrLsza40DZyGO2QUX2Cd8c+XNrzz1dpPaps9DwsPUEZaUZU
32hXcYcncynzXFH6r0TlTsEfozRw2+39WeEPZr4jQbhrO8m4OdiY61680OpKo2pO
GWrTah5vjnZUptHScpPuQxciuxO/oWQYj+l301P/BA1V4j3+L6RDDziPQdfJPEfM
5i8Sj1Ek8UHLY4JaoZfuHwNGFAv+HTufdHJul/qTerHjAZtCy9s0n6y5km0mLomG
UZbPrxx6qr2pj0PLh9QYha92hCtTzLZdqieco+GfXVfxIJYcUIl/kEbFhUjjA19T
tL+qw/5Bmy/Yyn6CVUMgmmY1M4o0h21t/wqPEFzQ2zaKXteiHNvM/ic7tou6opyO
ig/2KQDPm2hPwTwy6IDxb2mFCqqQn3VucvGyUxLLWnzMr2LiOCKooVAF5l3QACJa
GjH4UvhJo6PjvFxzb89fLM78V+z8mkANnG0JN1ivPjU+SJaB1Szk3ap+Px7G+yI8
G41Um3qowPRr9wnLIg+yEsuKet7rDcpfSpjOL9i1XiG7mqry7tYjpA7ceVoEvZ48
flN6qo3q+iXHCaO+RMPknACqbehf1iVDPxizpbDCFw7S24Tk6zJezwVa8jj9k7lA
57T8Z/5044DVeihjL24rD9i37HdVIb6YUzIogixZRy79Fikg3BM0mFL/gd5bcsQR
15vpIIgfDXnQfn/PJwi46tFjQEqxoScQtZmbFGSM4vxiFwAa8SVRf7clod5z4SvA
ILO6apU+2U0ADZUn32ix93eaNZ84OstQC8vEGwo02n5JHfNDiqqmI1MgEi7K6B3E
/gDIsrvitNUI+yAJy1FeO7tdEW97Cpa8U+xtdirczm0QdSpbF5bzunV1pc75mCpb
dkwtQtiT5aXc/nFdqvl7ssfsmKVBMhwU/eskt48JoD3x6X0oodCI1CrV1ZQe/Csp
pBonaqWQr0PWlhmFiSzE2MDHIeMSK76R7X4yDCBw7x0RfBpDb9ehdDZ8kfEHpuyQ
7Xw+bWDwORKsEgxXzKzqaMvKJZJKWSDdRnEe4/aHAjKQ8qFuiSvG9U15rTWVPnbj
1Hy3kGGqNZW41mg26XaBdRC/Ud2M645irT5KIPPgL4oqNf6mzVDtIXenhAR50cTt
B9IErElembPsJnrnzxNo2T45tIkAKafKkMEeO7UevdigW4F9f0XBmYi8enPxgooy
O0Q3gJticiBM/C8H2OUTnCxfKMp7cHfcHioHx49PSqgCoy11gm7Adg1yf0ml69GB
V+W4Pi2Ml6lGCugFj6bM3jdGbVgfxW71vsjmiw6rH/SIQGQdqT00hZsvUkOPpkcB
UWP11eVqD6zx3uQY5PR+zYlsrXMDxdoHkaku58pnUV3Gfk/rYgLoLPfXgVfOumQw
T5RZJ2O7dI2E+ED3aNsIL9c5pdUIssimPphQXSV9Hp43/7hXEuyaRVgwMGcCoR8B
qN3Fmn/j7fPP/LShLIDUJ5jsDW4XnPWJzKNayUOYp7RLDYb3bcgjr+4UFXZlNYxu
SQ6lhBgZGAIEQtQWJE5+0Z3ydrqIvH4T/URD5PSRUv8JuUiuA0HxVgnXn0eXm0RA
oIVBvy+ac8aIyJgWs9RSAD4ahJ05RqR7AjmpKlt7wH2YFK+bNEBc+rh3KKyVltdf
NulBLHhrvs9IFnxrZnLzkYEhKTa1Tu13s0GuslKRJi07Cb4k6THM+5hLg48iMdL0
ym76A4JIJwDfnsWu2xd6C8defWwBm6xCEopE4P7zZyoHtAyCaiy5XU1LwnZDdbmw
x3Dj9PRShBufEysO+3hLxvcDXSEyyaOEiFpiLd6+FTXKMgrEUcuL/eIoDvH0H+Ef
W01TaNAquAv03TUH2ySfMYZRJN8yuMgAn+aLtdGhO4ApRfDnOwbpJ039wdj1p+fV
Mb/CvuwMt0Dt1QWZe12Wc0QjJl1+GzE7o79Lz5L/BIj+QiPxwYPnaDBx57RAZnkI
tMMyFqXqBFAtzHTBi2PCOyH2T2XU6wUQgyfF+mh5Aw8u6I1igD0sGfZgfBBtvu01
E/7FWlJpb3/NLTzqCsBYlGE0j1DhexN+Kx+2kRV9YvAef3wsHQ8zg3iHzifjJX8n
UKKvCDsvnnRBJWODX0Zjfph4Z27mwP0b2wdwP3a+h7bE7/hAl4FC6fBYdAP9ONMS
e/FsjyaPDpdTqKh5MFRBTWjO5qJW+Bxw5bT6+hBcWC+ja4lupcHpQY3IIhwlAbca
7gOSOKHtwZ0T4yTyGTXYaOWPaDfMQMwe9X4fc9bmCbeUuWkoYKRQiXgquldryVmr
SAHk/1pp4i/za1/8Q6/h8oAOqrCGH4JpZpPt+x6Qpy0W6PTVGyrhSfBuv9m5N/Gh
iHYUv72CQ5TlQv9DMt9Qsnbcl7XwMfpUEJ/6oZ8wXcSltWZDaIr4q6C3ALlgk2KI
i2vMiWWumUNKNLU5cAqyGUYTzSzzCpQxzqomIyIZeLDbatwTFnirZm5Yk5t+DETA
hQKgEb8y2i2ho/h9vWMhalwRT0fFfLnDW6bLIbGL/GfYNmtv1YFez5yR4oXhJaU4
Wi2jsFGyLTLapqOAZnHCP7pj2kyEIbxu0k0ThC3k6NP3Y97NmZwn8+o5onJH48ko
7z3mdcYA0RyOMzXL8mHEM6Ds+0DVcNcqcM2Dl0EiVS+ksGNSbYtOavAVPlpqxd1d
CB1ZdjK+hY6u40HRA4f4+pE9W/ShWqknYQ0kevL6g6Hxp0WdBqRGYSrIJer/q5dG
upajuGq7WAw8vwjdB6gsctnDReeVUmjlh+vEY/VMpB5V7I/E7taXtobKHWAlF/FF
bbSl2lx1+DWoOC+QW+BNuqM1OSvEYuCSZLSxNHfa0iqPi+fkQz355O9PChJooats
Lll4rJOldjnvPGbNCxB7sLWeUJ3Yi7NqwHDTsNHXdiWSZVOcgQXNuCBUzEBwc9rB
pVP9iyceOD9KGefPeVvqhFFHlsgwPDvvfUDrLB1ULufBraFJPfKhbcE8Gr9N8CNX
LK2byb9dJpvEB5drVgfHzYnZnSFR5I9hLqv26fiiQss6Ff9WIqY4bEuNOeb3XKNE
Bz3pixQPu3SV54REBFDVJU9UVdghMQpxoRR0IrEHCjXiHqr2al3N8mQ5M4PvEGHA
hRlk/oj3DegkN3nhwScl5QFj5F8KXVHPgP/HIQLAgn+vNa929YRK1ZlxjghktfMm
wLfUJj3BxSZnacLrl9UbD3hiPzV45evOKDLQiyUnulZ+x6n//X6wy02wTkj+bbgf
/ZyosXn+SkKo2OHuvXtBXBGYNIPGFflByCDZg0LdzSct7EXpk9k3PnxCTXhaIOUN
If0j+cBGJnhl0q0NDGIEOZHEkltok77Z7b9o8sItdNiOn+f0uCqZgriZNx17KR+E
MYJaKUktaLQ6jSM+9n5PwOjZMO2GhvfNG1gO15e7pQIGBuvwBCTK+274BaCQYR/Q
0yAqXBE7U7nXMT38KufbkOAA1yv/TxnPjJ4UYf5L8tvbAfWDA1iF+txWZO8OPSuU
TVwbnWklBtkbZuO4+njNe8OkkzuaS+RbWyuexWmwCvg4FLTnFf4G8bXVjvwEXiUP
c2PuGzGcYe3Mm2KlzOXNlHhxEck8mabXbrTqPH/9MbQ0XgRmQSN+LtymCP+aI+L5
izDPUh6ga0kfIiPMNLVu6KutxJrsCY2bz24Ao9MFGTmA8VF991g68cvxvLzFajRN
y7Gx0qKb0vSqomhlEbhSixV7u9HG6z7jiMC4gFoQXnYdNj4WdgpC07JSu3kz2g2w
8ncdsq68dg2mPZwgXcF5cWQQixnt3bmYqBM67rCM1ExAEyWXYklkJE7lHSfP3lC/
Nwf/9RzINsYRreyQY9/i4XEZijDxubji9AOSDo3kvXXm/AyJsBJvv4vxC28oqu0+
38X91Y9kvgKbI84fZDry2HXEAVURp0eJ+g31fZjTYGUU0ibvHiS6R/gG0cBTzGUj
FgUDCf1d0GflzzsaPkjyumGR8MlfZRCSZChdq/qzniBLISUa3LvKOqZG7vdySCmo
ya0paOKMW0lhBL8osEiY3cdDeIMcEdVe2bmpG8gORM7EzEkE6JvBYoqAbzQ5RTjB
1+jN1R2GDNNrxcLZtmPl3t7dOJEfNGN+W3vk1vaqpOzvuIfmGd4zn8vHYcPrBPEM
tYw5e+NugXq2ZAtVUUp8bU5bSOkMwVm4HCHaWy9Ce9EgFtVcCquNlGktMs3d5jC1
x3shoAm7f2uTwMj1U9WShGrfxxlQh/wV1XcHNlhhEHF8Nlt1TH7adCvyTKsJejew
fb7b0vrs1im7nONobFafR84aoZKcTr+0FXSqSnjA9Xn3NxoTRJ7yqwOLCc0DYF2l
LD/tr+4Ij3NO1gMMarF0lAGzjxyNhSShlgIATnsCYauHD2dqzNogb/CtK6te0hhL
VDW9vNj5D3AywPxXzpiYKt2QFLtAEneS/V2CJGvwFopt2WDcZKNIshfT4GtE+y2M
4NFL13LeAezfldTYbN1ka3VirsITGHnpzRbIjcO8L/f5/nU0kK2gCe1bAe4qyQme
GbIdjx4X4ZrBoskSaKLeg8iRLOA5ACs05T5B1utjinpBJ2P0lltsYfPkDNukluBv
WuMR0+IAgFzTmiNXXNK3wDQBA8N3z8FursQLQXjjngVMGxs7jIkptKxvK89U/9CY
7Pidnuw4t7gkX5c9T1dFkukbc1181JZ5vBSQCCOJ5VxliZAFEleVst1EWaMF8Jjh
/O1puHswFJAeUDjlL03vqYdE+1X2X0dObA9EHV27a71CxdIfCjrWI6nHqFoyZS5u
8ZNaQFdR7fyBOSh62do4qSbWmNM/kLHpw3N+WQqOqTZricX6JXR/43QEn70oG0WT
4p8cXBhM/s0mNkiWWtFGsvadlpdJ2Gf2HBpIcz7X+ogLrGpvbtg33yglsNiTfSW7
tRQX34RjofzP/J/s7LSkCBh4pWX0oVDF3jLnRPPONcKLpexYMq3yzsEaaI7JhkQH
oCQA+moMqsSzwtkgpY3Qzxa9XBwVYb9CBoxHYUHwkLkhmsOZSdFJnzhGXV/OXP0v
AFDmG0gaRH8j6rgYzOXvbuv+8iBF9DnJm2bdkr0a+1PUKb7Zfy0D+Jq+c8tRSjKN
whek4UHuUKJaRkroiMpR5wSauz/6OdHuaLQaKwrg3FQ2JzPGdwxI2YZ8R2+LoJaq
LwPI/2idcJqHEMaw8c/WjyvuZ2PN00fQggmQ5/fn0oAflVp0T5D+yZpI8XXhp1px
3A1gR6OC5djvpa47XJSu1/7LtvgcmTXPuBiscRKFbQpbIF6sni2fDlYxNjeJV3EO
5+eZ3wfEp+jAH1uZRdcw6mxwa5j5SKiAaeyTDMxdQ7Q+EocWeY6Ye8xsqD6J/+tu
NJP/mNIESshSsyVMuRNsm2Hq/NmltVTev6XoA25IHqUE16LjzpfmHFAzh6HtvrCU
QbmlynNtUY4NqLvQc8cYul+wSq4+NxIKLVny2omhbXrHeDRlCWoKDx7KZ0+dtgnf
/JBqlMynXo9tv3sWX3InjoMYbbw/wJStLfKwWL6Rfck2Pba+uoj3pGRBW5lEUMk3
AhRTjKA3GCR25+iXwM1cMEWA3VlRZZtMNBDkeFuDkyJF+WVC4j8kqW+lw7peW1h5
jnX5NXuAgE5S3GIf8tFb7DfDeWflWHqI5EO2AXWQr9giC+yPQpkd5rErZ9QH0bz9
WgpzhzcVkVKHmjrrp+4CMxfQ0BYdX57WkRmEwfJQoP7OIqu8H2o1IB4muyZVQ2bz
CxCZHa5Rn7JmghzDD3IWpMeHMZmyRgnfpeCKZUs3g+IK9nhUosUibavMPtBDjP24
rANXbnR07vwCqeu4gHS3zMyhhYuObza2TdQi4gLnPX3nT7LhFSfViowe5pVnvr+L
l3o2AnQWLno+uVgOZAQM5MTOFplysjt+OGwifIo7I/0AZUNCUwx4P2YfdaSxwAU2
QosEP/mhl3lI2drVh7xSKmj17E6whhPtCtgkAZK+mx4WBbBf5I2+YjiLuSbWzg9w
Jf/vI+o2oBFZOoTsnsg+5hNxcKwy5Cf73Larw2WRqmt1geJbBIVigrVb1Kgb3VfB
dsIdvqD0b6d9WPqEgTM8S2+5ssPj7v+DWLfYfwpY4Cix0vqj/la0vu8XF3GPp6CX
g4Lctqml4tlRmzwrQPnbSH/0jSbvgoDvHAZKGbKzhHc1J4xacGQV4Ecv1Sg4CM8g
lZOVW45sCXkA/MDXI27EpV6bGeE2eylQ7/4jSypUAkktgF0toQ+OpDRa0J2UWqU4
fP95jfbuKpDFZFrqPqlL1rfi0uJcF5VVxVCq4lXWQO8eknusFJ1kDc3LOzkVjDfb
EGr2gtnZhb1j2Ge3ONO6AiNmIxTbJ3CAQdvZtnakofaZ7JMfkg3tabwYDAHvcnKs
C6FYqv2kRM7Vdl+R4ggqR65ObIHUMsRosqE+8RIKqe/0q98D8lLZ80q7FT9bkF1t
TyqcYJ/71IX+DFlbt9NHM8wkTvtrc1CiXdAI3aGqjjsevSsTNgUiZkR9ppUYert8
1P2NZSNO28YQFf5Nh2dxuplKrIVW49Xd9T3TQZQ70ny/dq3EqF9ZGPN6fQ61dfSh
Vd7CuhW0fUXA+dZ5jfHulqZdIv5k5rQAUhwBW35WdCKWBBxpPa0mDWFxReQrSSGX
G3WTZCsGfIHkovI+UayGdSa3EnnDxpGMIPhkFtTivfbb1TKq8Mq4YxVooGCuwJnq
npAnrdg2c+ywrEhRUPcRwRS7VCXj9fakMO1eygvDRLAD0WcgSJJxuT7GC1LapL3F
UT/CMCVkSGqe5gOYsAeXmvJSeW5sCYZ6aL4wADeABNe/aJWv21rNmqh3q7/DW1ri
vXkE9zZvOcAyUfFhgt8MEzuut8ZB+QiL5EtVHGLNFGrqEHS1olRssmWQDpBfhFEb
RbPVqehjUAzwvikSEZPjZTX0eByBu+s4JQcn1TjuGIJ5WfsR+7fhOThU0kPDlgg2
YfQSYOy9THoD9Z8QEIBFuhXh0XlVmVAamyqOz1tpw56C418tmD9u5hjv3Pj3+1uU
JsRNVvJfxRWYnb+p7o/c0xx0Uj986ts835pYic3vnhXdYVDc9utcMBsx44eOCAZd
76nlNrXM4G2uY9MRIvTsBGkPNnz2X/0uS1IgpU5pv09fzoGOs/BBKdenhEuQpccD
80pf/y+VcgLu5vySdAcsSO1I513mFlPmPQSuGGp8x/1U3FiZ4DeVwCPNhpCz3tii
A/ntXJXrBlsi9P5IhpA0ugeikqFPhlUMLPQrO8SNXNfu+0CtlSvD300DCkilGHNb
nR0ndQQt4bZbdfexYGJE/3MBiKEtPWs2wRfo30GirbWOKufB0vAP0pMGb9LWXH3O
khnJDtZHdmWMYiAcuAdPvWkKjwU7NkZXEVF02aBtO6GpWjRp2oDV82jpz8F8rwxp
mtCm0c033xghpWoaZtjnj3OmgLhzkfvhHaTD4/crf/0KpjJE1pFVM33K3eMEq0dZ
BqIdRlP3gNREDxXMlUsXcPs+Z/+uUVwnE/ut3Q2dmpcwdtZ+97DJuThosPo4c+Lg
7RgzNJZO/V+g2ici/aCblYiMDJkr0SOXPTlCtV/HExnm86TxCktip42Tiy1ev6xb
n709ps6VpHdVkW0x1cDw36OrFgwWBL1nGTTxXYvhbxkqglPEM1WjlTprRd6NYDEd
kkbFoMJlzb5DqBhumb1VzOSKmiNmK+L8X/QRamwcVtwAvzHQ6rooBHfb0kIo9hr0
cHvC4y8gZ1yVpIYMw1a7ESQqtAwnlFPZv+BpnXOLRmhQr863WdJdVp5gck/i9lSy
Y0Au3fNUaSbg5oJRnPaS0mV9BThenAUoTPHfChEKAMYZZHYPmszkWxz023l9SgZm
Ir9gUJ42yAAU8X05HdPipl01dXBhPUT4QpEKAayCtRmFuQqly0cnpsneeCMSsKQg
4pdBmjqMrtGFcMEFJ3dpNcADOQlKu4A9jMiMeyC96rboUkEffDB83j8vC2wlHeIu
b9GN2yqJGkgi1ezSfZQLmqE13le4LALoF8iTdR7h9mUPMkKwtyb+5mhNsotyOge9
R26KP0H5SDeheD0SOYziBZV7Y2tG4DbioZyr2KX8izqdnNl7gyHN2ekTldc7V2Rz
vFlBdTpkxd3zFcyT7jrAZlqumB3N9LSdWbVbAqWaDjligWKHjvhDYRSpHHj4CDTR
bPESOchJvdBl+kpEubu8xhii3KjVWxAq/PqXuYTfH1JzMOaRr+krveaRsBHlVkjN
DtNBYLusdN6Mo6zCy4bi53yiaz/VlLSmtNQKPlDp2EkGmgMrRjd3ffxzsdUhCAhV
zJxO+G9i9JDwLBmYBMWLEtCkAEhLzmLA6lTBnLyUolaCzn5NwO3ScKTbMw894Ft2
SxlNxhjcGcmu8f4Ty2aa1btpW/oc/E1rdGinrICrw+1Z2b+EHfENHXOmQTtIy1QZ
b8dI7IZCDUP9sFrUaUtk9FUULeBBrFTj4ammyMRaxhSLRWPXRTndmY/adR75yKij
ZvJjCuTxaE76LQ6RaidnrP4oKkOFuX1Fv+rfFgCUlJuWzbGdjF1D/W9dEI4aOHzQ
HReFcl8vewocEQe4wkBXd2sNwzaruD7512/s4kiwP0zW83ck0openZuKGw577/Vk
aXnwh1E3sL12xoIxOpau6D8wkH13QxEv0ad0+0z12uMdgzHaIkUU/QZKWdiidQrK
S+M4M3jmt8ym7cz+aeJGp4NBgRgSepN1t6CDO/ysBKn7PDBKIqQHbU+vONEQCk+Y
y9Sq0RyNRfbWXnKI2+w001mVVUqJjiUfzsu6120xz3aDv1aD/NqgKMJPiYNTDoyM
l0xVbHt7MDDTqiTKB/oRYHp5GAaD/5P9fjs+qAFnNPlUWWkgyqKGD5zdJtTjOOOA
S4IvH14LZR+bemRYVc3M+V44buu3oYyD2NJdZVL066EDzn39OnC8hsFdV96nrXxQ
88UWABvT5SeWODEB9XnwpcGbYaTYFvNOzBCl8jrZu8ow20NGtcfIH2h0o/W85HWs
jlNJrbyQfFt9lQBqEgVf4tWovj43IQIrIY/9GeB0gNf7nN9kUjX3zd7hYby/h82v
nPk07Sv/NKqB7ccNnpQiyTsk77AMB43hF0+gWNeTjS6kixCyawSZCtcxw89UxYMB
nQmTrmSk4lM6eq+NT8fcYsmpikHjeskSLuHpnbMNz4/cn9CqtPrO25MzvKXMFZCO
fwh6vmWwBhjGCCJc0NqIjE478YpNdcCddyQgdb8ibliiA4mnbuxHBJvK3PRQuFxv
+H2v7a9UtYColS+OFSzHo+VOfrCVJXjSS1Gtw1x4K1JkZpOqIC9jSb2T4aX1qGBK
ZCgEgius0yyvRitSAS70Q3jeTZEK/tv5LuE/WIKfX+X9QCpWdduFopvMtHAi+boV
nhHz22X9yQnXlo1IX8tE/hrXDb4axLNi87XrNkX5kdHvpBqqCdQaxRNV8KznzEpf
GWHS1aVJ1zim2GNAUjck2rGnj/iYeaya2NFdzup/b4B8zLQmdqrxMMK/ZrjG7OoC
HiRIJ2Mc9xKd2QKiUnETFUy3P6Wv4DppN5v4EsQsO8rIILuDfT9m4497iQch9962
JQD9J4Izpqq0/WzqluBWqyFiELTbJcO8E+kfU8Lcj/GGxcUCy6aacSQCAyPBlu84
rih3TqelgU4kibDJGUlyb/JX/cfVxdZZabm8jj0btTXMIk5dlxZ6/SNQ1WO45+M8
bQ96ARoP2f5Vz8wiB0O4lGmP9BgihQCiBuj8K1ffqZ/PJzA5aBnnoaO04qV191tZ
NSdFNk79OGD5pK7lF53ZpH7WUinFJDz8bqEu9dffF9KixMzNdQMvJQEgBm0/T7eh
cIrDy+f8FFRkbfpX8H2DBXY0jCwE2kTb5yFICe7R0tulabKxKd0cKatfY1CENVDn
jMA9WOPGBbKw2rX73XtGFSbcqlF+rS5/AShdS1x6zlsdwdovgqGs/0+RmodNvY/Q
in9p9l5Km5NSt7Kn8ty6l0RK3mh/RFNwEhtZB8pVwTJynfLFA42JvmGRRxuDEXQ4
6q4RDJENJr40uoyTSuGWCrQbMjts9T8hCadI9nIkpwLZcOjMQkftxL66Fq9v2QSQ
cZmo9VOXlZD+37vbsB7/GvvRP61IL0yEUH51abCa0laNMNFdaE4RqUvaIBMnHnIn
gJK4yOQtOli4+YsQ8M/hVvOrkKngeO936UyPbtOhGw80K/NtTFq7ji+MM5dCjVZL
KwGG/GfzXp3A2RhHo3wmte+zDHC1ways2GGm8uJL44zl8RRpcAaeyvZuOHKkfBcO
e/oCPLCzjzlOR2ji2WXTgDUC1+McgoSdy5g10jdBtcrttllwvC6rBUbJg1scj+iX
78kCadMHfTmBqgGEN1W3PJ7Nygv2J+E2cutN7tX7fCosi4iSXhqQ7wbrzzJY+cwf
biXCtiyk30dkUOdyJuWp24dEq8k1ESW0aDiEElzP7Lb57AbpF6pG37g423q9h1L0
IotUj4qOQhunCHLTp3bpi/38BrNgG7Mcl9EaUFNcpagS4IB+T9ov+bR7kkUU70Qf
1w54mJTjLkLwMQK23fiqEh+Y75MUVGPNib1zDN1PMZEvJESviaeKj9tMCmfSmM9t
QOLrQ1YMR6oS7U6Vni0vZZuNkcFWjddKPiq8Yff6zibVzKte5n5vRqvQ/CF2xSgR
8Dxs0YAP6m1UpwSxU32EwKJuWKSoV0W011D0KghfqMUjoPM6DvkdQ8gXH2QuJ4os
Z31q6Y2Yx7T/BvP+WzSVVBZEpVAuoippL2swYwy1xzkflKzs6EKANNPq9NU/PpWn
jQ5CovSiqmU3WTs6SBIvCdWW2d+GUXYToMwlmcJ7suzn92be1aWE3puwwnI8Vm5X
A1xOnwCTocgT+nWbLIDk2etlDG4BPNZsGJBxnR78qNLTNqZFXAGokJ1n4HD4KkE6
8Or3QT6CfM2jlEijVgONnVQKeNWsLLYGamBLrj7VwrYJzuIUBW+/ssHXWFS04tSs
72i7Yodj+eR6dVnUXsn9jHN71B0clLW8ySeNN+rZQk5pl7O80772tKgZIYgmW48f
5l+UfjjiYwqytouHUhU+i1lTBuS0U6RuTpKr7mQy14Aj/1jh0fx4I0TYZxlppPxo
+/3MNwPJJLpbEQT0ecYCyMjMeQCkefPWaiKeluMnNu8t+hMLHLpz2STE8eDFZD9k
bgGeIbWmQ485iIeK8JHYe39ARRr/Osun8ZryZo3Xwmdkt+aUrUeA5ahCSXA3nb1/
Cye/NOSNzmwJ3Tdm7Yx4xHe0yL4t7nqIft2lLxvhkno6ALoOmt3gPO4tMOwFpTmS
bRre5H5Zok7CAeqZ6VHIxZulgXdmePq9qg8aiCzzTmosAH2EeAWyb6XEZqhJ07Rw
1TqjTSIyQNA6WdMrWvzBYqFoK6/JpL9PNyX6g2dZnVuvYsc6wP/TVoUyTZbBvKHA
xzlAFIGPTiImVTqXyfHOLJ/OLNL1HKJTy8iLt4DsGUG6g1ghnFhz1uDJzqvyzSOE
MfkSH+IZhv9fG0zD8tPMywft5oQr+Uyi5KD7hOrAIiTwza14nAZUOhgdftc4wIsb
qrfe5Bf8/Ha7yCg8xGgnN8BroO0F2hDll/GVu1Yn8zEimuzv5GKxfp5LqFZv3EUR
fid2klwTnmW8s/ILGx1D2KX6CHYA1l6s3LGpOQUD5EkA6myoluCrMw9w2zz62x8x
dYq7lexOQPFn8cvgYzThuT/1rywLZ8T2VHWBuqc+3KIK38/NK738QkcI7uWCGZNA
30xFs1IZ7p0IEgRIx1gAOrdaAaH/fZFGltWk3Fbq3jAN9U4W6Nsb53HpcKlkqjSe
JUip7KdM3F2sPsJg95HBNtnKN6j0nBoxIwXQgaCbnvUuOqgBq2byUZyT2fGqseN0
D2H1bliUN5s9algmWTZlql2cfTBhv85JaH6YyAFg2NzBtFr3F9KQTohbRSTsHsbc
yyIHBcOh9/HALRKtNVICd2N2MdNiFw3V+DygwIrCTpD4L9inIe4o1D2H0lgdSZw9
fJ/yBx/neptv761BQCCc+OM6cy/YWOayPV2JZfbT3rP9Ai9IAAuzG3CCNMM1ya6e
4KccLl8xJ94xOC+Z0UxE5jbELSeFPGTVff3CMCGcWTBfX7zwud7v9iNv+gr+H6BJ
PCjP/ow/fJd+CoNiCBUV0irnVyghzd6vpMtFH7dE0Uu3WieXi7swSWKLi4Rg8wCo
mHC8sZP9chV+rSMkPIJH+MR62lOkGtxhHYlUKDCVXo9h6QVCNaKMNej/BUWyxmmj
ajr+fVubLxVSFaHaO4FUascKI6/8PEaXi/ElOxzidquV5Qoc5kcG1lhpErbi5KOK
jeLL+pqTV9cliJBTWzSr15zJftb4MWJZuKg/yaNHBRwvlw0f40h7DJolK41QHScH
9JSoRSAtevr6udgfmV11Sq+1Yg1bFZe4lYNlge5PeSLdKW0rGRUlbY/Q9mTi4Iav
QjnbaR+O3ItGvs+s9xGxDbZ1iaXWpJl2fTlhD+PCT0q4PRkvghKl59TkzAssXJza
UFolobalMDkHP/WmZgNeEWiGnL4AnD20oQEwxWZltBd3T21eIr2d50tuOd7p06/V
5B0uxVYRwyWy2j+85qyf4hdyn3Rvac8SNun6FOLsvcUFbx9UhEP6VD8QBwtmQoqm
LJIfzvsVzVU9491+DE07hjjC1eXPEM0v/++6W1oDPby5MN8iKXV+Q85ibUiQ6rb7
ZKvIgl9aToBSYlh40inj4+N+kGLPdLBcW8Esaw5TAMGsiyrrXQKhKjA3BfGkv2Cv
8DRYBcT1UHqxO879RF7xmWLpy59pYrH46ADHxJaPENZE1mK6ttCx8JXrhs3NOcq+
6CeUK+F2b6VV6ov1h9zMGsZfu6aH834XECVwWlZGAaPeXiNds4ToUgc4HC4Oilk6
KfophZzyMoT4Lz31qBQAZsqZbaIIFN+9LcW6bdKvoU2rBW6PQW9w8LzInoKBLztD
+cHGBlGKKIJDR6kIHma4kqa4Pc3+5RWvqZ+yowuNon3NcSjU0/80y3nlaFuPSdnd
Doh9nlTqAYblfWJ1eL2PTADfHnXgKQtFJrpXbiKCzkJmnorm+1TxKvnc+M01IpQN
bhBjyp5s7rUNLbwxaA+BlGVfqcAZv6ZgQhrvPXaFQFBcH+IE+BwULTCXkb4rx6XQ
/soQsQrZf8vF2zrKx61q8jaYZGoJVT215d1yCie1rhYQ3O4w6r2FuT59NUMELiRv
oVWry1eJTYSvsiwYo8+FnUlmTFLThlT6TSk5E/nHHQcJBztto8ZlBVBdHLFxXJXr
Ka8ZEYZkiaQ8G05mXa9TTg8mQ06fsl/JIkajOJwVYCJaiZQPG44N/dqpKpuYADJf
WSGq/MKIAtWsf/QZ+g6VrxBeCDR5AgcJ309Y1+18syGOiMMu2W4q41mQh1SWcegc
2XjczfThVB8STuyVuQypfOcadNs2e0a9AjKK/RY7Sm+Mg6IxJ7Zrr0glBaLINQ7M
AO+iDzBVbdtS4yqWQ3cT9QCc1+YQRrW64PVw+zK6uVUgaSv01UcCrzrSKiVybhgh
j2z9rCPuKehzjUBKNS7sU5YwNUdssfD2B9x8D4tFfS9WC2WyAVd9Vk4A8XekYil9
4oUSsMqgx4l9bG5EJvVjB7ewPvA60Kh+gbqPjadekllfxnApaInAVIk13yX0LMXI
QUfFBvXYHpNnOzKO7nqKSyx0Q/TzHdPNVCuUQiIFYrNjEo079pkLLpMf7VjCZVCM
HqQFdm8Yaj/JC2RYbkQD2tN7jxa8cAOgMyLuqykFfMB9AKv0AXallb0dLZjQWwW+
7gLFY3036ZsQYLDBOY//MUjaLezAsnSYOXJXxmi/Rr+MOxzpgxT579uuz4jJNuDy
AigCE54cSQLHdDlCtWvKz8D2XmDIV/Fjtvd9njquPIqZVZObfwlIF5CZSvySDQi0
/J1dlH7TWyDx+ViicI+DvsguOL5SrCWKR1W/DL5/DlckkFRj3JycR3eYMcZ9ERfO
M3upu1kwN8DimQxx4H9JpOrev3Sc/oXNjKAf4/pQHQ5V+uNbF/gwNugwTQD7srak
sexQJ9oMFtdYgTJlwjz74F5OhrPNvJq5iZq7jxUgjVFAtpR646Yntr8gPpm/+XZ5
wJOpIJ1iUukmG6W2BtUWHd+I4ewXcRSUvikD128BlgUbZTeyI7C6NbNQouI060fV
/ROpYW1ATIp7OtBZWmMGoWODPedZg1OWPoGMFDLtGnpQIG5gOPh/oNNPZrfx205Y
89jiknzPaKRa64HLjWgrO8PuUY3ykskpzcpDoizfTpyodOkd1yyzKsePZnYuOL+r
JDG3Djmx7l1+cHax97Ns4tZ5RWuvO7sqG/gl3sYBs5BKRygtyPL5y84XkYYMXtSV
jWkm8ccTEHDmekULH+L13owKH9okGbs+cFRr/4VFIJclMpO+649GxaE3R4t7UXsd
ETQuWUraFjPO3LWM1ZO4bJAlvnlN23cjxlKxQjcRXj6T2xhGhuBIT28oGJh8r5mK
sCkTVijgbVqRzK7IzZ0krLDP6V64mA3iojNKEUIQSifsdixbISCkNn1QXlKTYtFe
O7Afl+oJTh5FQv1aoywOi4/8ZCVCrLAWcbXXHlMOYwFgqrnT7z+5bt9JvdXFUaZU
a9+qTgTomO2jEOGk2PH3KhNwOE18d7SfkzcpvZ/+drYJSKiH8DPipW4uaH0Ra+f3
3yrwdlkAFASBK+hlDtx1hv2XxROjL1l+mKRYdhbWkprTW0m3BPDLx/cmgBWZS6xY
rwVFB0hnCRNpxM5HV7CeC5oydHcPeWp1y68iN2Cc/zGtIXIm7yKETeyJc16WzANV
kCBIrqu15vDKwtBHOmw2sKyX+nq0XpwMujZNfihlIjb223g0nG6YemHqZSLdO8JX
mcWPzOJBx3+XOi5NSg06p+vamrhYJpJDE9q27YXasf0AYZwO03hZsZ4z17/GWeO7
Np5/h5M7tdfsYKsS60BbcFV9xQ9EWRPmaVJCYzlYybb7cljdq9RKIMYz0GVKFN1f
8OPO9zXmIrKXvuJaI/DgK8ckySi6jnKm/wCfCsk+SqLNAhLHKrWle5hs99VJBMo7
frfy1kPIdKw+9eb1XfmzeiKQ2WFUM3xp+Tme1JAkhI25HQYliAdwWolsdJBss0aV
A6lSvKRG77xAA6DOn6Cf0pCnm1iqJke38159AOWv9AxVSSPYFAeIVWok3/8VD1XP
pE/OQ54f6fMdQpT/gbE2qulywTOTlNFF+HkTKL0UGOligwVZHaiJxGD8lc1EfbqX
trYYnWh4Rrs/TzK/oROB40KpQXlFTJcBkHxEvm2SDw9LRdokK0HiQYS9A2tHFn7F
5rdeHCNy8l7s07CBvsxfhq8vBQLoD3yzags9ig/Dro09uBCHKFtbeo3xyk5MbhP6
Nv+sZRL/Fbv/JsSS5xpKzpOn+fs6fYQ8VyuwgONLTDPpSucktse/rqjpEshG17vZ
utN5JGX6W31XoL+xR17uKDsyKk+iuDg1JIvBWPiVIL2BEKwExnG9Fq1TS6Exqf/I
r8JWV0N/QNy2xy0x8y9H2go8DXVs4QqyBLPCPhBmbS6b3+aQy0JBJW5CBrufs856
/U7s6EeCq0RgR8Q+zp4HQEmn48o+P3/s79gQ0b+4jAkzv5hPsi8gKdcPVUul/XHK
R1X14bPxaZr5I26YLLNPNgBwDNrurX/LWL1CuH7+64HF61OdxuLX1QRebJTdmQcV
qZotNF8nGm13/POTADKb61LeVo7dYnfEdsInZ1p42Kb/H/VANn/wO3qnHRBGVTns
nKmjgSwdcaNqhQ8eU2uVlhZDof0nuabL9q11mqkqE/X3pE1ZZ1GjLqmsqxgCsvkY
peAss1YDNxxAZtRF1qDl8q3DnBWrnXV2CLXjQWAqFcVZzY2NyAjuQ/d0wqP9lwgp
QhObiCol+UvaWvw0ADxylruPu487vDLG867I8IkvEeSgtqas9KG4pGtqqH61eh3F
0gz8dnQqOIITMSQiZB99XlkarEYPwH2IfO0OibJEV7qme0Zb4J4zZ12Ii6sQfe1V
AWmhfAyYBrkWEk7bEq29wqHKzYQSsWyFBReNSR+zSr+VPBHkPmHibJon2BpUp0hc
WiJ0v3yFhbUHlOQJdlZ179pYDUClsHlkRhjud6l5lPLXnj5UU+HdWuwEyrBjWxp1
0/VjNRVNNTaJ1D6/67NJKZYUmnYmG0vtobi4h9yKuIxFbY4Occ6u6+5x40Ro7bug
7IPPLCXueAzvyXjgF4Kwh/00+hCu5zeRJq55YbH98tBB12Q6lOifTO7JzlDxBfMx
cuO2mIsu+iz61nzc77T2uCVQfPa5FKYg84TJ4xWKs1P0Vi7N/LV6pn3XNJLb/m4k
TRYLSCe8VkLTFSZJf+tQhKHI/2IBDqJaUj9/oDp6eRU3kmvphuhFQiIiySv5pvD7
umJn5z25jFXYRh0GdmPDUf0GrE/R+AV5/xunJbbSv6Wv+Uiu3fH7UAv47iYZPeZw
holArLMWWwm2NlUTmqds0HdFJKpgX3czFPlfAwf8j17ryuph4rO+sQp6ewzuaOjX
fOIaVmt7qVTZiqceupXyKXhSWfOWpXHr3RVgSgweTkp7oNxjM05xNBob0QnJCm1/
TpxDGMl0q/h5p43+X89eaqMGY2sH4atHi4f9OPFb3q5FKQ+07N2jVQ64pIck/epp
kJnrut4GlzBNo0OPrXQHK4xoPb6LgO8bHetE2NKyBdqvRZt+Eopjn1Ml4mHTitc8
8rWGRoMFxiT3jCg1jVFjwulpThOGui9nDlzAA8bu9500h4iNLjmoAgGAQgP2h4pj
zvPfYDZWbeJN9UQv6UjF650cyXarGpKbYRYwsT75arvc9KQhauFOOYQSWiYvnhx6
GzT4oqumG7vGNstky+khiYAoh7WRQBbZ/IzKdVOak+GVKMHfxT+hxHPNk+qOVTiX
f7ig0eUxw/A7K5yKTzljtCBQGNBqqSywB2AADHdR28PA+P1CnMp0Rwn8jby1WPo3
6Yoyu7lvZnQwqUX+eQaEiwc4eSlLtr2DfwFBmkprsMPzYz/PaoKvMkMK4ZRHYjvH
ZMgCWQILgtIEd52XB3WeO3peQ/fSW767E27Q2NIoh4A789nDxAbFFawzVsQQnO6W
A944c1ynABiJwRl6jl2yswZ+OhBq+M6PxcvXv30mLnh3N1Td1zYWWNXy7BrZoYU4
5QJRMx4NGjVLLBRMf5qvtyFr3J5MfoNw+Lm0dHiNTy///RMLbe01aqRvIEgwgYIl
JtEv1eZiH1fMnGEy2trlGZSY0/NmRn+Aa05+5teqbP/VTknVueOCgT/0hiUY8GKW
c64ma62gY8HKcLZV9LNNxEoBD8Hg5cfnHf0mWihEGDt/81gP50cbGUt6Xg+ZVZbt
/mF7JNLJjdXwThFERz3xO7rJDnnnq6yo16GSaxcn2DfFb70+tFDhaziuuL+lJu1s
SRtrkfvjqNclhUx2blfOW+cdfzEGAbCZBsEOrpL0O541P+t1Cl8sluEfNZ12Vj6L
6/7RRCSAXueFkpitp0qj0vYg1hd0l0KIZO/6fukiYgTXie+P5j2h3cTXantc9V+P
jSFBH5zQkYN3UAggTIFdlSW77Y0fi/pBn4lwpx9ERyRkY+8XoMygbwDDDg73UVNC
K5l8pKbdx3jKPW0ODV5PbebgHYP35UG83oriv2ZOLKIhlGjyzZbWar5hgTn0sF6c
GesRjfr9zqlANRdt1dP5fWXO9NA7sFgieJ6gInEGSsgoG5QEifUEAF4yh7GXbrX5
OG00J2qCxJy1asP2BlS1uAozsW9nJBIYYZfeptX1YibZeXGXXZ1zteA4lwGD12P2
72oImEtMn1/2vv37xd20tR62+EiyADpAT9jpXYozOVgZEHrka/G2ZaYScRAYJNVP
rOoIIa1s3CB4UEyRipn+cwF5rz0cjwqrTijPpBvjgFKd+rh7JqZT/x3SdFUM9jYS
rDlzIqn2P5P44HzE31h/Zm6p7Z/RB4tQb69GzjVGY1co+B32PoNLo3nzVjEJHeX7
ukGUyFc0q11G/GRNnfwR1mS63YwrmRWMNz4DC2bxSLyapldvQJpiNgo1hohLkH+O
meJ8ZHlDjwKOrRm82Nxp6u213bVTdgrJJpiUxpqo33HWe4vYmrfN/UhJ0fN8C06i
T7KfRlsIhI3Wo37DM61HuUKR6o7/ctavfefaLC06Ns9LY3lPkAOU+qGADB+xowjo
FxFWNKAqTAI7o3hyDPOPVQsIUSbGBKzSk8kmhEQlVdcn0+AAWaP2PtYQy8RdgT6t
pLzM78FLInkmBLfwPtHpCUzvWzftJ9yM+faypEjDmTVkgcDalJ0Bqv2YjNdL/CyF
h5fz1gYzxTFvgJDkgrHr/fM57KhF0FJLYpAjDVPf1EHtBWLFXnOIQs6oIdBgcWGC
zLyn2Rdml/5Guxoqza9wQ3vwF7flimC4bQ9cY4KPe/+sui1EV0+massD5yS2VWDj
Xu+KyubZ9Ac4EBY5dCRotfWsT3M7xHo537cupaNMUWFAyVy47Lhkg9gRBZW2qPEE
wQKhIocDXmHbwc5mPHMqgjB3y6SdKuCvGBf8kh+Jh7bXf/7YUDcUW5zqPMA48l+z
BxmnVDxHRmmNL0WziQxKcikgfX9It0ARoK9kKfltN2oV2i4b6Iss/eyorRJdvHne
bSI621DBCjIBuIDE3KtBpaO7rK2e+wv7fv1ViIs2iKPveN3SbxHYNaor1bwtdGhO
Q/uGXRIpVv4sSE3sz1bJXf0PYlYLO3Mmu4qQso5batIRYBfVwiYcLA8jmHqEz7Pg
7bBPf+cslP1IdgWjbKY5Qy4TIbWs3g0hxYuN3plnySR8X/N6+h9xKsWE72rx2ozw
9vcz7APMReURwMfaUpovEe0+PcNaEIsc2QbnmIKa4L56IbmlGhF8UKrqS7cON7R/
u8Q3cqYDU/Q+jY4YiTXBSsr1R0eWWhHH+wjYSKGPdCHn842KEuju31MWrhzT1dpZ
PwpaFlhh3OGIx5fHyGpyGYq+mmT6+gXO3LaEDk4iWobRKw7ibAA7h7D0H5pOJVA1
x5W8xfGxzdzeGfd47pPaZU25QExzZgEnbJjIsxDIDDa39myLEr8aLLChouLrj2Ez
nNr+Yor63+wzbVHoKTHRU/sDw+KE2IPSZlrJ/aHFnlfdAbti+hrX36Qb+rE3ybsS
LoyFbIxj5THDOjdxJqaRc4V5RqrV4kktfoQyvmOh7freJdDvSAFF9w/sk1YFSN1Q
38cOYneGeP4IcjyNPJYmpC7FYhmJEHdEv1qLUYCP8F8cR1Et1evcwPYezKRoOLQ3
Bj+ZEt/9dUFDvlpib/HJQMvePf2ujZs+IA+dw5V8XsTZ6O25+cTve/t5OwwtYBXF
XhF9h3qnNyjo+ixIcPVdP64HcYEzJbBdjGK1ZoX1IqjVgvh9IvT6NHXW+CJVvo1G
E0W9NLlHFLJAcRkcd+w+FVYrSk2XMaPDAwnXcAH5eiRKivntIVdf8/c0JSwxM2Mm
SaB+RhhpjhALO61KTeL0pbD5KXAdkaQkqKOijHnMeK5gjmhSlLyIQs8hc2HGf7+U
K1K8ij6eOCYlGx3pZrkydlHKUnSVx4ELRaWNXr5HgPPA/Hsmg8eX57qJnUdDiakN
XTAMt1d+EZmKLSZtO+Gfu5w8vLL7MSIfUyVsKu8Cjcw=
`protect END_PROTECTED
