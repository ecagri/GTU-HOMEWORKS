`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qn/930j75AI5Vct2os1PvL2xTuI6qoDBZVi4i9DEftW7ussJWZMzCLd2XqQZyS5c
TkmOcZD/mih0pvIK7KbHxtJauQ/bLerXPqWYwNOlU+SVkoHZ/xNmMcupsV7k8Pwp
KQ89XiQdDZ74QkFnM07RHdvAi0X0YzGeZX0pu60zlbo22eSkeptUvEt9Zu/Faq3e
7F7ULRncJWHcw0hEipTOHBgv236phVpEzSrprPAgPerQxf/tfbBTe6NPl+0d8NZ9
ylnUa9Um1k8B4Gj7avTfDjvbd/qZVX7nOzhO1i9kib9ViPPSlpnNnQfDFUOwbd+0
Fq5upnVn82fz7lJWHkyfKluqiE0AZ5j3LFzB8aomuGac8S935TNhKY06JUHrg2rV
gXvthuG73tOI5P97F23UW1mcUKhtY+agDu1ByvbLJ9MmrLb6JKwc9hxmD1fNSAOI
6fxscu7wAIUeQtUGUDmoCGQGkpyRw3K2TYr1h0NJK0b5Q37/paH96Mkz6bN2BrGc
2ODxRmfNfUsDeW2W5qmen7dXpBCHzLf+LjKy8s8jNkwuZXPxtfPv/Ki2Et2+G6TM
QV+3kY8yEXt4MYJsh3gF0WDrrnpSOVlNDtkeqPV1Xr6JHyuH5mbJF/WvYQXdw7HV
GVAmn6A0GCIReW918h7NFYs0ZDJwTppu2mywAD2i1HhYRk1M+dE9UZQPDgVAkLLt
yQlsyk23rVex+Ag00dUV1/mVXzDnqaNQBA0bqQuFkx0UK7Hf96nWY6VQG5bLK+Zt
JvmZoy5MyNbq29qejt5fpO0DnsTlhHPWeB7PiLWjjWXd4QqQZorQoxvKRB07PR6x
q9HOcRwBA2FOPogg2gQzWpEOVKLhyvgGDNuJJk2DHMwrLi5ALLKA79D1ic+cMqoO
iErQW2vHr6s1ukzvYPhG+VX/RE7pSjpDgJhjsWc+7wytE94fVMe+5fmksIMYujlP
PbDusqeCXvGn023Uk89EJJll6D+avWeK3hWnTlnkH9W9+mhZGvrTk7uXdts9K+lK
V+u7fu5gp/e7WGHwNKYD5MvWZMNnzkUjj7zz9707c0bVjPr63oe5B06POQoKlSTV
nLkLe4oKx0DzE8BJv+Cvkv+u2SNFwGZsejvBef17r+bJhsIfkUqcbe3tD8cX8M+1
OsBzzM9hlLKkMUnw2a1QBGEkmBxCFCqLsg737+uA1aaIzOxt8fXLZ6tHB1ZEckBC
kRwVzmlcTbBMf4SY0WMyLL/iwDLJgM3Gfbyi50dHM6DpQ3S3RfVSoIZvL2kzyeD8
S50XfIq77h8CeSGS8kXP7oKVKnf4+4KWUleushBigPsxFuCnQgFcvsiPTlZpE6Zt
xLLkJtKphcMVo3jxEvQJrnHxkR6IsnKDYfnxSiARIhITRpzYvjYB55aL5reWWnyl
wHABsjBxK8aM/3wfF+pLCGDB0l0DewG/4l2WM8hocYcjUIofagS4BR9Zq0sbyTt6
9Aybvqw9HvBnPjxBTEc3yXLo/DLN0beaDHkfxDNaf2HBkrSKht+OuwKMPGXCheGA
vmvwrXBrUoLWBld7a3H/R/kBTqKyjwyLKBurIhy86H0Os2BAQ3Ke8E1662WkX0FS
TjluOHPL6jEAwx/QPFNh1DRCeGvsRFItuENFhXgL0WWozzTrDe9d5JCkzhIyft4z
mp0skmaJQ/iGUT//gdYPxhRuIh8JCZEBljqNSFGMnvMjBH5/XtIX3HDzK4XiiUOn
Tk0OyEl9L1g83A0o6qs0B3Nj7c7vJtrSTHjjR8uosvRHg9OrTwWXchM0FI/7+Ok6
VQXjSEYpPjXJklvIJAXYUcqzvw2hP661gw0qwHGvFa8Hke7hBUP8iZ9rlNFXL3G3
N1bbHsaPLVw4oYGAK5X+NFm/aH2/KI4iytE+bMzrZTmjXKUGi57ZLh48OamYaAtk
JUbKrDrwiAfOFcDTknmSh3QAjoPpRJlYvXHFmxzixdAKjn2d1WjkQMXTOgjLp+ap
0Pf2OJauCe/QfbyzNMyVQZenzkt/gSE7GjXqyBjbzUZMk35VM/wxCWjcv76RyepH
TBUdsT8gGWYMZa97MfwL+WvhYyIqyRLEcs1uHR9k/cuCgP7C8IQHRzbmesxC7Gs8
P1y1GxDstBnVNSAkMFAGLES8QHwE+3U4yhHV3QMAWrUgQSF91qSWDZpo4/U9DHgB
SXnNhmSUJhl+qHb0f1h0l+ydt90j6XUZPVvA+WQnmgOk0lye/GS4lAHT+3oIFcav
ssyRq54LtNtIEh3ag8/HQYLmGYC/g3pDuiON81Zm1hw9ZMI/SNJ8mxKecoy1yD+E
lPLM9PSPqjc/i9tz7D3jgqcQqiiXBeJslz0FOUUvtKE2UF95bJ909MRvQgqbXwxk
9yzYtS/M8tDjpptqXq6s1LfAQ+BVfmO1qsc28/G9gs7VzKBfvVGFGmxXMGupUPK1
KP8I+3UbSeXKVNP7m3xdRUUKia6FiA8UHwPKUbE4DH6kpd9eckkjtr4agzQHo7Dn
EFFNv7t1PK67/DhfJcp6PbYQmmLeBKtjJhnREP3AP0hyGG/bxuysFJgmPabs+SqH
aUK96VcmzPDNrNGrGUkk7yaBgByc9gsKYqkGs8EjpMP4uQ+1j23fetkpBb7m5kmG
9968+v1Sf3WvcaMYCI6rEjITQP7K+jX0pdcTCCcA+Dowtdni7DChFC/P9muPu0j/
AzTot/Uf44rcYI0cIGkR96G/8SlXC7OtfgdiRACJHF1gRAJ5Gjkb9rbY8ZT72lZc
4hDb1AtArajE6TI+gPNV+ELL57sKPcqlQN4OqdSdAZp9gppwFewzmPweLC2jiO+V
lD+Upa8QE3CYfAK7PvaMzIZ70knRQthiQTLX/oRZiD0eVzUbpMfLIiJCggQKSXIx
pDSqGELb5x9byfMgrRWMnoaHFfyV1D1HeU9+QSQnOWj/44Y/FHXnveEXPr+yysW8
VSnNVbMvv3o68w6EDNVlwPgxDm0+A9jYcaYnMHedb43uoeLLhklqhj1XaPeVplnq
Y0aiXxCcTyWMN54hvEudAFH3dUpyPxvd3n4SR+EuEpQwi4lMAdI7JMcpT1EQQOnL
7eFmX+liOx7rgTYO7PbP1HiZGVCPPXUynrKQ250ZovYPwrPsjzYOeSCMeLeEDJF8
OxI/7zPs54dGNhaZ9zNSnARpE3h2c+DXKd9NdImDey0fQtlCBJ0VIZDHSA8SPKL0
uDWy8EKM65xWOHSbEc8i7dpceOatM7LfYgcFx9VmqenD2IsnlJ37kQUhAE2cu1/J
2so9IZDqQ3bciKlqe+LCQMief3sAW/hWfGmjWqY9CL+ybBrpyUl/PWpz8hzjjHmx
o85qnBWQvZNs37Qdo80kHDM3hyoo44lMZ0sThwWdl/SoxEFZrXn+qPK6XooH5R+s
0Rm5mM5Avlqta34JSD8SJb1cKqOggSC3bj7qVwZCa/dvzUCQc/I2cPUZtt7vMHyc
q4Nu4AGdeHwe6FeY0/q5vQZBR2zSvVLEDTlc1mHTdUIa/W3DNeLmbQ2UmcznUBml
Jw56P9KdXfsGZ9mH/jasP2Rd2wBU9eXivQi1LRNZuH5KRQNvYmqasVHhoRwRnYDj
k0g7JPBMVL2DrpHW1BBEIcrBJN2bSPyhgVcHbg1sVuhS7/NO7rrnwuoHPzV67H4m
yX6frh9R/6yR/SSCxdffI2iN2qyJHsynCv68xSCV6Or5i1+aWStGst0RPa/3BpL1
CvfV5yIKF/DAUdeBNBUaPnv4xYOZUFV5isxSGMEybAg918oToo89uqOZNh5cbPNW
wKR/DrscsSHEr2o5unr7C54aCOFlEqg+TtX3cVhjzA53yqhe0hxV03JQeBjmdwey
Nszeyo/AT5/w7TKpiIXKtTqEURhwQDWwtUxRqvdoz4S4LwZBqRcRdhjWKi0bV9Rw
Rm40lcfsChgelgLn7SxPbQWrZpkUEVy/srH0wz8BXaa97UpnryiH00r/tCA348vB
`protect END_PROTECTED
