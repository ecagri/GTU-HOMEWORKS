`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mpJzC/nknYJE4eNjeatpP8vNvEG/TqFcNnRiIMdIuJMNMe56tIhAiDvBTIh+ppBx
6b6mMfMSVck3yy6Ms/sLZQgMV11QVmqSDko3uy9PPS4rxXJmjXBiyuJyXeM6oFJM
Uf+9mJz8vu1VHS/VwB6zwMElG2kFQgL/BIPQoIjRn0Io6S01/VHbyJHxE988R4ls
yQBR/8Icn6wLfArzpseCoyMhWhp+y4mETinQXwTP110Xh57RHed6PHmGnyh8iooo
DEVeZTYs0Ytodomy+7Gcap01TBjfu81OGisYjamHnj+EFgA7UF035BVR+OgRjHFI
x6l0DoJorLf18DyQpuJWtyfWWdoJwKJXZVhumhuzN0yPxqk+NvldgNbTZUURweTK
fakJid234CbuVrtFB5MjUSV2rt1YodR4qba5SOFNNrMQPESXgxMxZ8WScjtFDNof
OGpdZ44j0d1n3noIEws8EGsa/sBdCLy87BVi7EuA8sAXc8+Nk0qRrLwbQi+FsgY6
vDiXpI3O6aVhbN0Mr4pqQxUXrfi4JkrpdMhPuYC6a+KCinwzs4uHXBkdmhU055MM
gfh5tCUBy8DcbLXqjOBNJu3gUyxopvSH7DhvljVZhHdIOWadJguvSHVZ8bUo2Sy/
tTF+u1urcV60lSD3ca5wbQBQ3xOGSV4iSAMhehfgoKApeiP7sy3FC/OM7uh4jDP6
QDMvyth+Fqznph7OrYXz6Mta/3gLRULGmnDffBaDG4D0EQqGhNddKcaXhtUTVsq/
KVYXENqVuhNT73p/dyKGK3XS+Y8rJ8/N5TA1ZxjKOR7G95fgORV1m+V7+EGWta7p
uhxDFmiyZrOrcj9/vIDL40qtEgzlmCWl8drHIFVjImISmk03zAnNwfFkcASjhIcA
l+MVm+zpdwkIuNEaWxCBymXh9P4jGdpskN7A9Ara4vNmWEf7H8k0GZj3TlF8Jxv0
YD6krRzep8G7FZCR1Gz2cpk84OTvbdjOBUUyO4yeeG7FHbRueEGsIFR46LC3PtoD
A6MxUeGagoL9PWMBwBxislEwmMvrvzeK8M1tkq9lEu6KqL/z7o+XOQtSmYjM4oQe
g9N10wSPxnuCBw6CIBvZ2zS6ESG4IOLUXVrUp8j1GzSGR9kpDgvzC/x17Hrbp2AX
g/h7emvlBjIaszePqIUEhXD+CeGfm9CLulFy+iH3Y2ZPQejPkwdnNUaen3yiAVs+
RnGDusf+6VCU/9bgfBIDDelNR2S993TEq/SPVdRtZgR0HtVr9iWwAZ0YN++B5Tkh
O9cTQTZVt09lKO7hXMcStwbHeI5gP+C3H+BeVBPdNyWo+pod9EFjziV5YQn4hOeX
w9vEam55Tud16E4RO0b33nG1G21UNW9p7GLqaMkGtPvFkYIzLtVl1hY8niImPHDU
Oc/8jaIJmLfCvEXjEDIPlgfeyXH8IYR/MEQEWqtQAG3/gdj8rFOwfryh3SH5/ifZ
yOe48GikpjNsCWOtNdgN4ULEp4sNDvAlk/GRiram0fMoNsDh7EQmTs0TS98wSGDy
P1wuaEEnTofDG+zgVlJN30lLhq4NEMzU9sZElfDNthn245HKDFOCZpBuCHuNnfhJ
HK7pq/aY1q2i7/gfygXEF6fOzu514xlktPyZmNqGwKX+KEVg5cfjf2I8pLEL9Wto
f1pJkHy9wKuqwp+7znHasJFDRuoCyVED/l81FiJz1DjebETifbDzw3SFjxo40SEP
4zKI+E0r5hpFnB5+eGwqVzaycUyQ+FlURjBG44/mamVN+djHtjpDm5ZAPEpiTZa8
elVIJBy4TFQy/p6kVR0CZ2uSNqvEHq/6XAMcajBEAfCX8OOYnyWPoYgYrZbdAb39
1gbwAzLn+S1tC34lOeo20/Nc8wYzQ+ePHhbRH3Du+DroQI15VxG+NZmtigXyLpgB
t2nY+4EHEbqSLwpZiGNgKxqCVYhUN+5todI5YDQ1feN9oVgvobnvnVd9+sXMyZok
V/Kp9EE94X+VF4mW7FSlDtOU/L15VW8zM5mwY9vuBUPeMuM7ZK3DuCJlQ7DwnUBd
TV5or7+i7xdCZZEuQnRHruEWwKg+VRqWQjSzAAlcxIj4q0c33CfCp6K/ZyL7O15Z
pqK2qIwnNUI4+ykPplxllirl9/RLckduHMNqXdg8kbrlfJ7rFgg8CSi4a2dYjHYE
eNpc5VTmZ5anF2m6HUAs5JC8HnsZ+uF73FViOlVMPD18Z2qU+spwIOJNys8Yix4h
t9AyQg8yLLkYGmjnwAtf18bQ81yWmAw4HXKDiJILPjaOhptpBjuk0Juja3P+42sE
PdKNSBlM008YKVknq9yT6JyibIUOAxUzm+Nt05C89U9FU1MAlFRTJYbxDa6Q8M2L
W+M1btqIk8mF74wcFdQOghQ+vwXQSCa866jirVy7Tm86jWr/J4xr6I70BjotLqHC
I5R6kSiEyxu27GPBNoeuFXcY/eEsvS5zlj3CDSkraNi4Y8uGC+FmTncJOqmdOaVm
WqXboZq7/WAHJkCXjOyCZgQrvqwkBACkutxyl/yZJmfb/ZKyzmNMSHz/7amLOH8f
8ruPdJ9hoPHz2e2pwbsfME/atmKTncrMF7LuzCYn9ikK+CrNq5dHZfl3Y2JjD8yL
1ZlRmFtlVGdDZ2NlWOSmR5fKDD2YZU/YHO7uBIkIh7YzcEekPAhFCi0fJL0MQGli
xzib5PEVvSLNdKev24itnd7WjJaYNp1xgrMAo+8Z78HbcUhlfCT2jEfmTY3gBchj
hnykZEvzJRKQRSR+YzYdv+/p1KkSKpwiJoc4jo3d4LlaUB7YkPxq5PSYkNj7+0XH
D5OJ0qvC1t/YxT60GQIhd5VS1AkaizWZjZsIWFCH15D7b2wJcKPZkcdtQxCw2yc7
dyZ5j8ZLTJhB2pWuM3og+fwBg9jpVxu+g8NPAqbGivkuA5Hn6f0BR6wHEfs7E30G
8h1yVneIEaOsnQdXXbq6AlaKQp2tnsj36pDisivdlC8=
`protect END_PROTECTED
