`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ePVeHcXUGEXef8g1yWz4aZvQnf0cvDhvFAkDlgoNcVNE1DXRkjyRByy0Iumwk73X
Odk7khJUUnsYSMuArzFH2ODSIIJvoyOSaSCFlHQOVr8/tPpPN7ovI5dxbKJaoIpW
gYNQSJvrabPzbv40CPAKWVuKsvUmDlKEeBt16ALKNJG3gX1F5fN8KFeizKQ6YG9x
ZU3Mqp0XbXogQ7P53PF5iIC/T9j9IZ8xRpvI24b304yeKEWPN6LuxYWld2FKrHIT
25feoA4Q0AWdJkNR/yrCf6X6ytIHZiWWulHq00AduG3yVOa5xk+4NQ5Jk+wzofKh
YRZ8mYeRdW2ypxySbgGKt5EWLcCx+6A/Gc686FwamKKk5k/5/JkNPRLprMFkCzZl
PbYNDQVnXDNwAllWwOzTxJYURBOGOobZRZp1pW5GZ4470uZv6HaEgfAVZydsYMs4
3pF1PDsFolk2v4PU5e9r1vHvTTzd5ug3K7dZfI/+dCxw5p24QClo7eBFdZmxqA87
Od6GbzfKLN4f0fMBcn8UG95r1FX96KOS2+z9+lPY51lWugr2YPjzHzYViRP0UJbv
0Vn4e3TGegOJgKhkhxQdphhiI0wDFLRnp+/V+GLXf+jXj7Gl0mF5UZoHABldy+Bs
`protect END_PROTECTED
