`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iBgcI7+E7TtPeURLHaRVY7v2i4Q/6tN22/Srm4PW7RKEHijXYTo6DazjfpBGarku
pqHdBRY/dES9AtN2frRGCUKWLIfHoHBlqgDjgDhFY8pJeP4HdaBWR+sojwTorG6j
bC5I4UuhRGeoQzvF5LxCsolb7jMkMoFFIrgzPHc5kZObWdX6ILvfy+0vt0prjd6+
zvsT3xTwEjH9sv+mhIcalfjJN581+VAb904QoHJQ0+kXaVdK5WAKOTAv+PYlGjDo
YF9fr1FTP8EYPid4hP6j7yCeKkNVEhpuPBhUlJVZgkOQ7ndq8KFepLUrcKN3gc6H
vpsZDkR/c0qHkHwLATyLmKv7dLuWSXWwbefMOM0iP9whRk03WebtQibI+MPhQP0W
mszqoPtdjiJ8WUQKvm4VnCllV/QJykw7abv+9IxM4iQRIupRfJdebtqLFdghonrx
s6cra1PZ973iMHeuCDGeSXoc9wFOj7AkH8m+9lN0LkGJP91+g01ZzubZsk1O2fEI
b3CCaZMsPy3Sn6AtBs+xjOXWaWPmN1Vhsv0umU8YAYgpi7hrPjxNAGxFfCkFa2pS
1NDglgn3noToz0cn4Or4tKA70pll2s4mGuAE4mixE3U=
`protect END_PROTECTED
