`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8aOrCLUA8WlE5dw4th8IADcyvrm03weY8kCXlHLTveV6fiohHtEF8EfckY8hCOmc
CaK6IUuldK5pVzKnCPiy34dqNxOZ0Vw4H4M7SfH4Dan708iCWYIxqlp4uWPHYrUG
rBzRIipaK0aO0vi9iDLLL+UI8pqym4O4+vF0Juq+8mj+2GUxTMYYl4kKlir6Sg1T
qqQmMezhXz1+jazbZz4QKd04Pf5oUQLM7j/dViHuSSOOuL9Q+8IwywkJFof9Xn5u
DM5zyqistRnBkiOwdb+KDAQaBRGduGFS3VbsKTVHbVCMcFL8+s2ECa7w8u9aPXje
6iY3MDYQlxhioqisYXXpNGHnuOMJBSP8UjwogodeVMSnS8jK+KGl4XR2GnHIe+rz
EmIUE/d1SG6Q2bx0GY7RJ+PZXzdHi89CK3192WkStXJ8yFhx3fUqEA00+5TqH4H4
PiwdLVd+MLuYWf9k1os80xRzzDfsI8r7N2cHU1/6eqwaqPPkjr76pVWEYDo3vyLV
3aKzwQl51Rspj4C59MDREGbfyh9hQzzNoMyd2c7cAX4X20+7+58Ne80D3gfYqe5F
Wz8wfAoxbzO5n3DzUfNFcn/RwJ3hw7dhUw0N+37WplduNiRsqEcUIvVLAd7COo6x
rVXlBsAokQbNXFKZ/P7u6KhRIAkV8Yxh59Nri5vdbCjeYi8bf6s/Q2Cs0/3v6LNB
n4cpgPJkFiwkoo1PxGHuSYvIcnscH8I5c2ST0EAVJ20k3dERJeNn1kuqt34MT6H0
OB9V8VjvYc4SFdYag/NWSQpbpfaiyIwZK6OkkhVFo826fmGyCQVZBGFf1lDb8hMr
2gwk2QlQvMKWdFdapuGNTo2WtwiwYy8u+6AoLohnuzEwxunbqA3UaPntX/c5mPb3
wO2wTcb1ROWuaDmlVrqOvakKABl8/7VbdQqf+1V6zZmHKukl/pWrA/1RboVFJH+h
ktBudhVDe6ow/AQfMXYq4ULPU43Lk9lbIOMpTDIoPTNV39ObElx923wcRRBICx4X
2jmz+/RtENFxnjg2/K01wUQci56jk5oTVQcjE6BxZZ1m4xs5OpB5Q7o+3SVUBxeL
0Btqj3GRw16pPrFQSZwK2ms+3hV7mnQW5FImUOzT8dBGKOK3h52mTI2fZ6yd4zO7
xr9a/B4vms3+crzTtUMc10AJ3uxHZ6HsaIIHA2QwfqDUbg812JFuQtvILn79e0Yv
vYmVFr7ypm+/TYtfTVme2NvjIp1oWxFuwED+cwU76SiaokM2RlsTgQ+2rHjoEOH2
T4LIwLmxASzmrWzHmLIere/mLUz1Ho5VrWwzJ1dz7svSQgVJaYrOyTa2CtNC7KMn
zgPsn47W1e07MovqJv6aZH1soWl2OiUf4eoc+yyQymNrXORkepIHxntYwfyc4tnu
1Kkjp//GFpOUA/0XBUym1IM6O9DO5fbcLBv8LUpqvsUMTOL4+bAVZy86YpITwWxz
`protect END_PROTECTED
