`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+ON+VdLmDYMlF+zJZWS9ysDoHpszFHwPepx/qrRx9FejJhYhslxnwpmtJoP6A0Bk
0GiFNaRfDnRNoeUBzsl8l2xDdtqx2CRn2dPq8oL8TNl025TK2BkLnjwugvzRdSTk
m1R52C1tmrCxxKlAwBN933ETeBbsSIYsMhnNuqbNGagYun6u88mYJwR7Oa+xjotE
drtxtXAHX1xTg+uhMTP9QfL53WLEzrqUve9GsMwqcO50HVoBcMDYUTuqECq+FMQk
zI91txQMMuaWNR6Wxa5dL7NWR6yh/6fB2MBSBxjES76NgKORoWrJwFi8HaVG5GIB
iJwCbIZxkzLr28KET6IvDfupIPNgWBA0TjDyxQhM49hI6xjjkWMNz/f6/481Jxtc
XLB8G2/1sIJWovpmLrwruFR9G9PfrSMDhGNWoovKIoNY4PtgWjKtFnhGfVenmE9v
Ad0/bqYVz0wF3wFfDOfLBVuRoVjC9ao74AcHSTjT6BDGnpnq5jkNmBE0qHHQzSPt
AFssOZ8FAN+F/pH3LB6vP9jPYgnzY671eqbDxTnKp0teH6KhsgfYM6LLOICAgZ7G
Wwn3YPD6aBCzDxnkD98q6qIib3ccnfp/le3zJt34CKmlAeljhhx+J/zx7DQ7rIt0
yx+XWiQlh28lZGmKpN8ZfA==
`protect END_PROTECTED
