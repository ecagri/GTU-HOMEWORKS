`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xcNXKnT/2TSTdNiuF0wucqzArxKpjaS57tGa2Z75zqD61wpEOqHJ9EJey2qxW5L9
0uP/nlng+O1N3bGpPmXcXXNuz48pS1JtTnGW5+4uuNDzhAiMS9TLIvYVYE4f8QeZ
JZVvJ1TH8yLIj6GaaaHtqt0biHgWDeLV3lIOir/NPwc/nd6xoY38jZbsZL5vigBd
yIyQG2zH8mLyDRnn3Pejg5+j85NGJbkjedlBKoUZ18ydkpx/yYm/Rc3vtC0BXKCa
qY0wui7IMjV/jx+22233MHAACsgcwypyINUolUp6SEGZ5lyVd7jb9i7yp5H4/Nz9
iR98/KrULOda80jISzCViBPDD1TKrdt4sBLCyYsy48PzncpInUXpaR4wyYU3Z7bp
uqyrWPjAED4pTJHmtWv1M+T/PSNiaY1yz0CtZtWNCM+B/7PhturHgUshieLjFzJN
Kq80B7WkWtH3eNM1Cm669X9xMasCXxv7cDdwXx00dbdlXhvy0ubjcsPg+jT/G07V
jydaxRCd12cN1hBLHVEwhz/mwvTeSi2swRcSy/IooQV1Pt43szN01HaLcuNbHtb+
QmiyX3vhCj/RNWs9kImahv1rZXnbpALg5+sjee6qlOpxF5b/B/xtD2BaP0DdPNfz
nKuaYWFamzEGVYDdRB//Hxl/F4CFttE0JU3QhQXG+k82hf9osMVKrVF7jOSXjlVJ
3VSsW2dHS0in1UUihBwGdNaPT5d9xHZ1bJwRprRg1pIFbiGO8b88xbE8zh5MJBnk
5MhWh0k7VnR8bO1EPSXqz230wRetXb1Hu7HBrxysC6JIEvnvzps/xwxAwBF6S3x/
ZOH6IlZtYpEyJiOIngxoFYlxkxG120qI7Obx/3oQ3FxACKCjPzBaOw+BGkveGPy5
9A9QqnOBWwqvvgikph2VLkz2scpgbWrEF9Wt93hGMsBMwmQtuSXuIYDIRk6lW699
HNgYRNYgfluRCzldA8ed5KuhWkH9q9UFzo1P+bwn1YO6vSh4uqbT02FZoqapuPzn
S2oHESFJSNeFHMuTRPiY4jfQkQ01cBwjZZPew5LWVDVKv07fKcf3xqC69hsRGAKP
RSpy5JpH9ub6TnXVVS/hHMyP0MqOP0OcoEbPRUDASI+fWQi0/CD+lMCB+O9LtNsE
9dicltzpEBW73K2KnxL+OSnvJk9/0lAMCxbCLXzeUauzHfFW5otvUazqo+rSqQr6
1yDQ+b7CLM9QZHvz1MPnynCCgxGAd5aMk4K1vogd15Nksw141waOx0InQ7qeKj+6
XVJMcsumxUU0+BB70mEvppr6AT5GdPIMTXFflHlcOnSghB9gzxDGUGrxHEBoEe5i
ngcQsv0HArwSBLZlEPiwQS59hm5wbiG9JeLT1e8yyaLgKafVNLNGhy+R/2CMyyOY
zvp9f8RiQ8SDAeJbJrBbuCMuqAq6jMr8Z1SYZlcAoFIoeFpsDkT9fOn9uFdWjwU9
6c+y4srmsUXkgbFlYWUMPRcJmBI4522LoLVCoMXBxfH48gRlXhjrD1+8JgYymA1c
B6lkefaR3uN4j7rZu7C/lys9DvwFTj/torY2kgUqd6a2anovkOOd5Ndq8NFxIlLj
iL3766+0iyxqukovICc7VmqutNlkuKw54XDYGP84FtRZqTqswyCH0OFjsui/gQzY
bChTwolyJjVvhdx9Fn0Dj+FO9KMMcPfiUp9FNOdAE5cYaahGYafqog/AHLXFc0KJ
uTBpScYc4d+nw4O47nJFJsX8uSYmkceC4VO0vuHE6lQUXc2Jtvyvt7HvqolBQCPb
LAedB+On1LULbMO4bHSd1HuRlynayoSCHtJGhp17E+ddqodymhBPF+i/pgwUTLqI
PrYbUvcD9qbBwusVqirgKOoAAjzdi29edro3IJhgxMzu0zYlBKwJDYek2Bg+TuUF
/a3jISXNmUZhaie2GZdltKNLqijeZiebmJNdg1p29Tr7+gUM3rB5k081iDPeQ3l1
08b7vGdCwFoh4SEhsMosrqOR/Z/S0syV/Sb2vc+5tFG+H4qILAGKJ7AHEI3xQpiz
bwIxcTfv6ppUNbcUPca9GJ6kAv/udVt8H7UIxexeZAC4d8p/LTdPSqtCBC/mM7p+
RFpFwi2CTnB3r9TR0FGmBM16/qh2Na1PWTWR7BSBV0pUTMJQpRlpEj31Onazd0P9
8iyiOu4bdTHpfF0UQ2lrLhK9JOYJRHOZ6Ht8W3dl99Kt2UXUhsLPB0qdRnb7NgcN
Ew0xuyR6Wvtt5zW3edigW3hXQJ1G8OVLrimw1e0iR6ueFTekc870fcULHlj1rZcx
deV0ydQcIajM4Rb46C3NT4H6l2kclE2aOEz3EOc7SzFulJ/ruasaaMsZW4ju84G6
9kNj1nhPAxUC+brwCOhk2X6PVGvEhbKJep0au0cBhf0po/o4CHTtn7mvmJBoi3Ko
WpJm+MkDXs+mxR9hmFmZhw+TdhPS7uSmW1ziVwXqZsa3lNHS0jY+/TCuCrOPtwDl
optYJHp9NXTFtL6V0jPtSY2NTTtp3IEg0yq7Vh2HcJfmuOm32gjaisk7m7kI8meV
dS3WJ+DbhIPajXeAsn14wRY4Eyf0eVjN23LjeYc+6ZYyvQduuDXSTDkK43chwu74
c9GqKo2mXz9uyJrG4V38RcJzAeT2FQp02KKR6xWzMTT6vCWjYqD2lyTgSR44QmhG
YmGl5pIs3w9CvCU5Po9NSi2aFH8hyUKovJKK7r5rSN5aO2zsHNNpxW3aIddHdjPT
0fMgIRfVAc0s/rALM39zNYOysNMKTv0fGfgK8h2bT/YWZ+JNevgQFfCnBSw7+LBu
8xA819dIkL5NncKlomE2c3ScNzccv3S6VAO7teJ5Q3YjBCMrVAKvdWXgb6lWCOj6
78I6l0KONScyDtjZUcboCjaihsHPsx140tINV6lNHHv6R5PJanmVJUacVcQulbow
KK6lnBV9pbRNnk2cNnEt5e4ts3y1W/Z5h34V+5QYVkeToGVNDyHYPECqV3iNpMFg
98oP1hBjRqnfwkjJ6pRDy3dOKfm9kcCDKL4s29EHa4mpTpcEok8f5yU/ytaiKvCd
xdRFbksD0Fd1Vv7BPm0Y+1ZkVwrP84j1mK+exBiHoRgIgoAFk1QNphONDNaqE1Rd
AHpivUlG79MIwDhLtv6IJ7gdihg7PiWGdceNkbVNOuJHWs7jx+ZFqx0zUzhkeE/e
jv8t4EUFXH6TftHUcAdgoR4na5fOmlkucHIsLNrTh6vBkyk7lU0Y8/AplRiJZFnD
1N7MWimf5E7Tgd1Aal+4NMPybu2QnOOmoR6L/rdvaozvA8ao+WM7pqKnoO8ffDFM
7WEtcGia9QvDZ6NEumqasiaUvdIcZLySKqMg+AjqOOqaqRKQKwEqP2fRIyvGLC2G
udswdmq3df9AKlc9E+BsnrpDHneeKMMKMgVau9XwpCkF/nLXDgtzOHwx1YSgYsns
ew8wu5XyjYaroHkaiGWaR4hGcaMcTs1J0UqeiatpXTbZEObQhnT5NS2z73Ui8XN1
eIdQcAvVGzkENpLQ0Jj42CEZVOlKrBLdmcl8q8RHI47zvKjAWGQf9/ypbQsh/ek5
Xu6Zw/eplvv/CY9SvTwzhbIF6DFLE9FFavdMAJmbSFwx8jNKvt1sNvskldMHHqbN
I9ZODMqw7FxIMZO/tKXSAt5I9L8lYKEdNbNNWcsSXW3iG1mj1kR17qHp936DU3M8
2fEzom86V3rqcgaSJksZ2SDa7lBDhzV7TeodkQmOSnplGpuMMzzOg/1nlGdKo+jc
S7IOoS4x9DEWrHJ2vVBy4yvVyS9aBw/uoRdJw999A0Y3EOKsCJilza9Dr0PvKhWc
4la95RhV2QSq+5haGJKQRk19MzS1eRi7B9dfDetfDacg5XHkXhtlD/41cZGCt0on
EACJuORStqRo7wYt+ikueaXWd7xBlaft0dc3XDe0J03moM9wUqULBMfcyDg9yB4Y
KZPFRzdhXKF/GZiJT+WSrUFHucM18l2cXD5AhxUILvDXOJAiRjIelhwJFPxWic1n
6Z7PAJqXY9aRioFjZlWt37LNSvkxHwFonZF3UpeGvPbil2rsbBMIzcKFSN/Ch/HZ
`protect END_PROTECTED
