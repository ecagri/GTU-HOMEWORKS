`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KNWybdOaBrnYT9GIw1OyE6jjYfFqnuygoonAPeb5YYrItyLGm3FkcAmwFJ4L2xLl
Vl+4Prv+8MkBjTr8AkDyBrJA3gvUyX4+PouD2rZIRb6c0bYo6sVEWkyBb88Qe+r7
baVuJW1L8NHhjuEcgwEh1sKKCGRL9lbWl5zUdnaUucPaqGFtJtQ4yab+03JE/veB
04VriqzwkOd5ee2+KfEd0ymsVXScY7KSmF8WsKfhJ1WnvLK7yiIZCsTPytjtvXw+
Ai1OcdEGYnDjOTvwLS4FR3mmPuK9LGI0KoISXGNPD8EgNse/mnbIN4JBW4s85uJO
lMhacHnEQlrlxP7bKteZ8XieYdc0M85xkzfDvE7YZvGcyutLdHezjoSMl+lzS6XU
atlMRRDySw15VkjDJeTRdGtAPmDV3GVIF5B3+GLTdYNwcEpxq+Rg9jglLtKpxuuT
BrYg99c4b3HJylOYssTgzquKTdOpwoZbzmVuxgxXAYJaYJuT9Ny08ciDpsVeVm0i
V660c/yXEawWCr/q2mXXCkKLIReoMpUwBRTYtWe1/TwomLBRz6Eyceb2EvWYjIfH
5c1dLVSG7WXs1c7x+OZMFBmJQw/CLZsAW460hM2NRfXMeS5PvQ12He94GniJgHl/
X8BpCnpwB3R7rtAsC1NKZOv1346kh7zYON8lB3sQ73GktNZ2zsL8syk2esqeK0dS
lwt/ecidQBlm+n3P0F/Gv6OgyOVW+0k4Yqnz/taNeeQ3XtHnd+wj+7+EXMJThOJb
YvCaGXCWHt+gSIw7/6HtxDQdpWeLmrOZQ0QURYkbyAp/C0TetzDl0hZWl/rjXtY9
2I2UrTfTQ747CecxnISCC2E4aZMcPlt7SrilCf10REqIPjpmyaPVG1bVwvTnNLNg
5yGJfwvbSJxHq2uODwhItoq/+izsfJBSG7528HTfZpmpdsX0L2fmBJspW4Io9Tc3
gj+I3cXJAGkzCCJRpYZhvX/LPMBvzfK9bfo8Y6nCmiHarlBDDyspZflif9O46o0v
N/olRrE0UFZZUN2D1f+GTENaZK0VZKcW6B+rDfPAxZKjdKtA+CNKn4q7WdgbpIC6
VqKrpqgPTMlBUaUBncEAALGrJ+98vXFokPtzTT7DYcH8OAsaQzvmK7fyPHsq9d06
ugYMJg1dL2Fj9tN+QSIKPRqopSNcS8uJrNoD4IyftbCrdmY0p0vyaRN05lAxPCbQ
A1gJ3swjMRQ7An29pjSwSiqbInjrObbOQbCIX2w6I1tq3zdZYO6XcSDNId5qGV8l
dplImQm9DJiIwIBTmRl80yjDklB7PkDTAKr5JERD/vkYVPtKGVNInagO+ItBYyXU
WHoTFdJYMNyOJwSDLrVF+kvJJKo0Vr8goEl9+HZJ3EAmB2pzdhsUCLJix0j8ocJO
nT2PwwDbMZU6pcUgUgw4A8Z8C/CdjHWQCiDStT/d4RNHvCA+4VNNRCsQXPi93euc
WHWWnMS+6mTH7FnEZEgRqGa2SBxhsl2KMAg/I6Ba+VnBLXJYcElk0P1rJb1781t2
XUwZPhNhm20ShURr8YTBOQ2zvzPUKL1U+wDoeizXO07yyyTJY6eC4qzHGI2AMvle
24tgE7WD2HjdDxPye5WpyFqCh4jeh3LzvbO19bBXfeQRKzWHA8iYs09/mbnWcGbI
EesmwfcuxwI5yddAE3qx0Reea+hQCdyGoizBPG8e2h6vY2t6CjeO6Iu5NkbC4NrQ
xlYYvRBKPZOvAFYcwxwiAmrazBklOGy/ygEMGm2DIO7QpbAzZQkeOUs2eLeMtAtZ
tsIQa3PLq9p76DhEoMmbkZdtV9U4KDjBtGNDVWyBc7UuWwI+vQ+6wUgVl83ZGR96
o2MoadO8hEmwJCjXj8ZoqDT/6VgIO6ORSSEAHPInWnNZ09GAkVWUE6CJlXvofPl4
MAz/2vY6XTtKqMF4aWAdY3cS3+ALLfumZUaofzRWfXvyiq/3NJdZ51LjnzKy1ip8
3UZkIOR5X0nQbWqeENCZhZuh0sZXu4o7nKvdggjHVYFD3MkaSwWNbF9u7t0r+cAd
Qf0Iz3z4dgUGfVwtMbxFnaJ3HotwDPYdy9+pBmpijrk4F8Qr91SOLm1b9erIrEv3
vMhjuqI9lesTvBmJeyQqfV11ZzN7fTJdYkklQIu3cFbAL7wZt/Os+yRaPcNtYzdI
Orvfoh+kJ0pYJC+5KNy++dn0Pl8E2jNBDEnG9FvBe/FtS/RrM8PXF1lp7IfqKasB
nuM+zHtmHEXWStaKfrJVJLWReuy7ylSXO5Ywpd6/hq4wfRQk+/GDWzFBx1Raa9JK
WosdcXs3m4uokcKOyu9xXDqPdyZU/iOlPHN73lLKxDh1WHtJlhcPO3aveP7I8lZ6
8SK7pxNgEgKh187mj3AwohnVFxu9JlHPePViQrUvRXL0e/F3wrsuqfCgGm0a/Jzm
6oYPQGLyD+oLJSsujz6VL88N8az1xge2v5GYuUyxdFWWOBnL+5XJ+TcJSa9PPhxo
qJUiErNASFPLVH+MC/SfDMDnLrO2PpasMnxDS5eah3k8i1edvKocP9B/aw8CQYxC
EU0+gkrl9KRwIEUiKN3GQeaCL6LEIeF7FWqUozgl8eEWw0r3ns3AqDXY/GPOLusP
yXwWFitfydWlG1L7OOxSqOwJsy2QPAULheRDefZ8jZw=
`protect END_PROTECTED
