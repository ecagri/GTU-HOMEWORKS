`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uQplNHkDwACF1TTRgMvVrRrFnFDAsTYhg5oaFE4o01jCxPFqgwo9wsS4oOL8qTZV
gcWn6RcrxvKO/zIFvK6bCfMHAN6YEOIJL68oOTEOM1LZ8WpDP6LDy4GPTsqG3RSv
eoUQuJKOgV/5ug0+3Rn24GguMkK/YKR4nsOR9ksqyq1IMC5fM/irkFKlEo6wNtER
Xo22Z7iumh0HWCqIzyWu+y187IL8CVENBNvfTlCM7WuN8pqcMZxXDUEZnc0ETEWY
74J2K+I9BerWPZbyUQPBQWAUJ5PrI76+QeC/4tKtIb80XdvuwQkfQif8/d9R0ywX
B5KpHA/vwj4QS5wZa5p4rw00QcUP/1fOwHNfrZaSPXSMgcj5Tb1obdz9px68ovgN
QrXm072PNBrhtaPVivUiBreDJHjLqr3OnWl84Sn7stuFnBZgvWdH3R9TTwTLWm6x
p65TGwd3O7Hv61WHOazPgikoRM2xYo+GRsmDa7u1XY5hg0JjOoPMFpXAxBX+DjcC
34l6RYy+DCJvHVeDn9WfsAtNNa0Ym12ks94baJlM+onRyMQ5mANmtZlkSmdm4LWR
aDWBo5fSL80Ky3qKa+dfyMfmhJS9cO9tVCpBjyqevjiwybDf5Pd718Inh1wX+VfX
EFi5itz4NBF2KIW8++cht0asXa/ijyamb160toPLk2ReudZu6xR8UUpigwrdMtfv
3Z3lZnv2VXEGyrGwYMoxSIeDUVlvdfyFbJkvgVXQw6HzgDELs07OEqzwOK8aSlfI
vxfbRVUElQ5fhRKFwHjVpAxseScLqR3tYPLfrAdzEDEVIUPes3xT61frpTdvXTBZ
u4crhTH0VqDYOfMsGGFRdNAGmrqKBMGzF/G0mbZ8KrYBsxukehmA9XdCBKDlHJBL
njGREVbwWtPBbdKngyoR/AKpZAFrXBWf4PkkezK/SmbzJ0KmhgoYcbWrKE7p54+O
IY2Hr334feb2hE7cu2fHLQ//2sLIDblhktvGq8BkMz1ZkIdi3YKZSHqTqNKCuVDx
SY56bESYVafbMvGOJvXuH9jBsSA3VxRuSHf4e0/MXTEP0YPvQyai4n7ybPg0MiZs
drnLr+tjjDzTOVps8YG4DXIWZIM8Uzv3WHUTuYCi8dFpRlbrtaO8ejp92QHulhi4
YOhHbYhWDcD5ScWOLP7JdEdpYYWhT7przBnekq7utIvfv7ydN4H/aPf6ZxrpI6Ii
cqhvhjbM58TTNml58x4VJgjuAzK0iUBb+CY2ur1HwcEPpJNSMZrej7qi/09n7UmC
TvdoK5WlCb2g+JHR/lfPkl/8Id5UR8AalVDZOwZe+nbDKQMcZygJwBLhvzSOaCJt
jk8zNrBo07+dCvWneMqDJc6ycosBAt+I7DcWEisPQAQPmOIBIn6e0bbXvtUJ5uxf
JI/hPHI5p3L8LPQAXQmPPVDLv9LYerBcJnFEileNa4NsxpqFolvXt3SYX6YE0FN/
ex1gVXUg5q7FMppI+o9H1CFfICRNbd5JBe/bgSumB3s7rpcsPTIlHutfy5dYQdI3
1HwseEcu7a8dfFPHrn4MO5TiGLN7i6iaevLchM4BUjZBFrZk0CFbzGH28fq7dqtS
U2CxQLEluN6Iplz9QuHbSZsYz3EAtWzxrV8jkkJ9zPBOFTk4L+7b1A17g7trVAVZ
ecibeeBmjQp3OtTXA8AY57RaBJacnSTB9SjeHSQceXTwq5uS+UCTd+f0Su5GODRW
S+a6rJX2r2aVWegVmhNNg1CStppjyyx/Z56P+MDXx+eBOgP5vaowBJ0nDWbnTtir
yAtGRYCJdQZ+ciEOPwzjJQziPZacX8H/TY+9dbbqf5h4G7eu+5pkpm+O4ODpLTH+
1qHmPavEJR530mappqV8Jg0UY8bfLDi31xzKRPLhdgoh2vKTzLYS4y+l2YCf1/j3
sQrqLy6XFVy6KySCya3oTyusOMc1Shr2svZy8tyiMXH4ITxNb86JM/V3JJU7ZYEW
X3gQJLf/WtxsSljTIn+fLhSjUNyGd2VHeyfGwAYDm7POvm674MVwgGbq94RXMHH4
dDzZS37IoX71Ua9wsqQm8zvYK5JPi4EtBEmSY/0xtqP4O7N8cB2lU3/SebRzim1B
TaKyLealT76iRzhAI/wVAewMfnZX+Rgm/H3disisBo6uDB7oYZW5crWXlT3sGgzj
ocYG4MtltAzReLZ6Y5hVcw6x1T/L5qsEyAdLa45WHJQTuHTNXhAzrkOLza7+w+BC
qgeLf6y8FsP0yzdOAfx80Gtuy+c0ZNJvnk179gJ/+Lkk4CYrifL2lLXlZtcFazv4
mpXo6xRBPCSoGpHyxVb7cdP9ZVLYdaVRngw/LbpXY7GANf9+ROiNV5TMSL/t2yHY
a/xGF4YIrq9oK7nJ9SvyCZfPxRkcF0+jbfNJfHPAbYf9rzNOq4biVMyt4eXnaEQb
BabG3ESkherM3uDMfOh+zmIcWe1+64hVZcgqxHEE1coqCdyU+GQ75U3BpWUQ522b
axO7ukWuXUa1HcmogYV/RZRXQ4XsKz37Gb3ORSB44I1K27pf5dmBWf0x85C2RiF2
FGAvI1esKPx9SG1nhFe0/pRHYYHnflhU5L9d71hFOY/gALOQ2EXNhP7t/Yba2wxh
9W9PaMhBVhjCe+lrU6zXBJyuHaYHPxd74cfPlChD5vSHTcPwoDmnXf//kRSBC1FP
wxYrr2X4/oyFOQXJbbH6P2edaT5fTNehYBFTWrBgnxvSuk+/KDXqsdmlddQQZeHx
0k+294MGL7uNbW8sEktE3kH8yi0Nr4mNi7DaOFu7mngNgwC2ZaqoQVxiYZTVbpzQ
i9RO0hPlg29TLuDPaNT0VS1J1m30koGMGetc4t8yqHfF2CcKuFnqNZsnSIQKf+pA
dl7Y7syrbk/Q7TsVZvZyHyWYN3CV9lB0GkQGsHqa0n77q5YW7Rg03hvJ4nCor80C
8u7wfDR5sBnAFZ+7s2ZLzv5qT1PEfkmWqABsGur3rbvhXs8j/T16k6n3E2ociXnY
WGaogiW6nbfl6F8/SyR9Jat27NjncZ1ru64ufP6oTXb19FKp80pMh+HBCzvgBdKV
/jG3SIKekF3i4ka01nrxQsbBJSjQIVE6WmSI02590fLQG96DS8AoE2ZGhCp8Q1wB
JVBrGzlvg7YZ4Qs8AP0Wl3Wfxd/fm0eoeeTvTDz6zito+md8RzOIXWa+AW5GB+fr
az8M9UeYGoFY6BNdyy5ESApXpx2cG+BkJF45WKwiSgajPn0qG8ar0jU7orIl5Yon
naQaNiEu/2LCD2Q7f51i/fc6UTYouPvfuoET78DUsItCv0H/aFOQ0xNOCFguCT1f
ys/Ks4Z1tg48kLKF3jQ2wYp8hhH7sSYBJqqXNJAk7W9UU1TNI4zDFFacI93NznFc
TsMuk+LDWuI8QWPEQ27tCAbdiAlBkAfmnpsq//XSEBrZviOEcoX4w3zvaNXFAxd9
xyNop5F9n0MtWiEuoPQIn4dzW4pvJaahxPQMmEao9TCS/1VJp2rZd2y3MVy9h9FT
rw5X/oummPswn24MkALo6YRCIuw4FuS5TQRjHXoxVAS2i4IEOz7pVF6dgfgODWKz
S/kBPRCPFM/aWa6xvpCYTBInijoUfHiZRfGys2YhXqV376jy6zdnGjOFzUNDOxyF
1a4aaKoYOkdfY5mwbfWll+B5xSmkp0UCIvdxv3erT4jMFS5eU2/uvfhgkkvFsloq
7hH94p2t0Ze4YWb8gknd5pgr9xbhU3pw484n842POYaej3YizW/plqwENLP6e2Xk
sKmqqyASAoMmscPvC+xVY0NOxxywK9MyX+WIHuDtznisbxsavl3VvUkaQH6Zpimn
M/fQ6TLBoeh8CWz7nyFHjbhfqjq0cIobkGoWwVIw8WowBVdbVrjP9NlO7sz08nv0
c/AFKgZpZE1H7F+wjNGjxmuWrdrb4979vS8okKGcMSVSrQuiAfAKUQ9yzbs0yXMZ
JOi2aDa73qYWI+195qwklSc42jD5lermErB1kOtbl+iD1cKElvteMKgHV/CBrfXt
pgjkUcwgxifXzO+yzdaBsSVng+5b7rJKXwCYppxpMoFpHNvqlIeqkd9b8P19g8Ta
hdOG8OJTv/mb+KnOMKD73T/oCIkiiNyEzQb/f4UDjGg25RPkqDkHMbrxoPCrODD+
3dKjH5EdH20Ks5ndxd9vsSjQMKplYsS6UlLSha7TtEUxhl1Ad+LmS99269cSoeFz
/S32QLMWz15kKFhHCwgGgVoGd9wupzETvfcTEtkP0vBZr7lSbWfjJnCEvVJ8S9sw
Wb1m5ZSEWNaGYvcgZsW3pCl8IpPhCINgeoy/6y7HRJBQezEKZhPKvBctfdFUZD/b
Ej3jGFtmcWgAuIttmIcbSR/aARDTpuYp03LlmBpZT+D4oyEXS4Q1zYz4UWL077tS
PzuCv7TFOMbz2G/mTAd475N44vcslkkEFEPK2t3MjUQnrKhbKA4cnO4P713lMaMI
tLChtvEFloBILXieSCD55u6aauKGs1nimlykM2OxbtZdZY07pkysglppLynTm50U
dL9hllpsT5/DYbwmUiCqsSquUUni6xcZQS/NTKZkTUBjqLzeK7KVoQUau7GSGRXG
DyIg3/5CT/2Ja65IUmgFy7sCJp0nc10K/z3sMgB7dfDy5KNqrUXKShcORd1T6Bi5
2AQIu3mVa/XL4V9llcioJQOYvIrpYxkDkxmi+cKn/IfO9jKqv3XBG1R6gfM89PdH
6Q3o1IchKutAUFAt4x2uc1H1mqqoM9oyClvMLCXVpayj/0itp2LOO9pmxr7+HESe
TwhuwruY2yKqMDtNGlm398U/PGFCymO1beiETcTAIIhsRgT23dBd598vg9pL5Dr3
w8bvGr8Is6tgcjw3yU0zXIs3m+gVZwDcwEBVJB5fd2+j0Qb/3t3gqY/gQMZL56IO
SBq0RvHAtoqJJSA8ilLjmto0yvZhNolfX0Nz+ApMvtQfjFGfPAFZrR6/c9RvZo3T
YiOQHfeTqd7NWuQyeerPuFs3b2NvSWBve5cQtRWDI3krwbsPUDcn6AkHho+r4MCy
FpXMojF4NlEID3aZrVdF/LcU9YT1hvM7c6oCSR8LNIJC/5/AqUX9XIvuQOfiEH7g
WhhG4ge5uhj4dxwCuUyIbjeci8AN+7I0XoJIRulq+17ChmAkPCxDClpjiIZdOPj7
Vf9DAzIe5AgyUeQG5PVK9VxLucnlDi/fl7VnjxcJtNGGk2ezvEeXIL+WIIBnmcTr
lN9yjWeWVZaMD6axOiw60+BbX2LyEQj0HLBn720C/dJZJA3OcrMEcxW+tDhByXMj
OiI0NvjtOFButQh1DFQlDRYlGuUoo8j7HJlERBcHO0/prPxeP0UcLFPLe38+CKFe
FNxPWr3iCGW32DA4+jVgg6TmqU3fphy05JY9fsdRoggIa4OI0P8pfRkoLfzw1VC1
ln0wChuBOU92UStpycpjLVAzE7pSnL/4RljkU4w/MoQVvAd9hsWYGhaeIhxfSYK0
ZUmQqSfx6S6iKxX+Gckoh65R8CQFqS0oLKPhoFwai465MJKIUJMVF8ZhsJ6WnXgT
UdbDHtNC6v3uG4ppVMvNxRSTetClDNotRlZU5E4ryfpdH5Df+M0wBeoNo3rYEpDf
KNfcYDGuYUeASoHX1UIQs4hu5yb6DNauoWestrkDA5l/Oi4B/5Ed/UrBBz3w48as
jH2ynG/HiHkPxINo9C5R1dGsLCw4SxvgyzbB69cWuhBUnOpGD58VIEdZ/E+u5fMh
PLnjM13EiHXt6Pov3hX2gh6DM8+G4yFFFEk39UKquIJWIpT0HR5DMfTyoz6b2Qql
pBdZCsMmg9X3PWT6906YXXJmnEYgOpEUqSw8jU0qKMjJACFOnSxniSSE57TsRy5H
YK4D7VTcj3FiJaNKtwfev8Icu+sZCQnLGvQ6OMw8bMPDkwdEOrD+wcrX++R1aluj
6g/jvJKbzRJa1fx4oZI6XvWqXUc6DecOUdPT8D0e5Shgc135zsIvZx9YaG0Cbl30
0yJKYi0Z/hJHmaxe0tsdkk0tX19+sKsv478SLpmxpg6YYb4FOFwOm1fHXtqI3+c8
GpOIVxR/wRw4jFhPn2ghqWSatpXVPM0cxGdywY5kYmrN3kL60HwcyXVosl73/5mQ
X9smk+etOnRmSAg5AEBECTWNmW/Tei0cNes2zGW+tqED0DSbNI/m0LSRJE+deAwY
HeZC5UItfJMQF8SSOz1gyCjbOf6zRGNnRYPcLCxBatb32b5Kh9X1SgxvnIAVJZOi
e/YdOV3aXBiW6RRU8LaJ8ApkBDY/FyoZeu3wQw5X7Ntz9Ua0SJidCi6HNprzgX8T
mxqiWPP9WTEpqbaJJJE2AlJpci3gxGkBGSJFP5InhT12puKExtYhxMGInq4PI0cH
wJfs6KSnt5D7Da5b2ri6wEtJHvMpl/2VfWFbIrAm92s7Hg2vm2YU/qP8LLpY6/5c
nzpNN8CgSTQLoIXZyqFRxBJTN7qdlrOhrFOxa3q/bdm4NpYYnK4QVrqXaXbKxoVv
kRngt8Yw/cU0xzpUHA6bHB0A2XIGYVY6yPoj+WBL8nxAHhragyR2dQ/sRDgkxaAG
zJGR6pSMd5qQDeXPCbJ3UB7lgJ35XpPD5VTtcwP4AV1bZJ6MJm+hmEyr8astAX3J
VpRXwDnagpEkUqXXThPbMHCH74hEls5Lz7qbkJ5KlszHYz9GhOaqiW/t9ta15VpV
wriWlFQH1/NlHwmGrNP9WMxDPGTQNFzkpOiyFZo5M0Rr4EO/bB+Hpc/Jtrs5fv6u
C7ZexcEvdt+RqBBS2bFQ7rw00oqVW4y15CjAXd2k1UynsdlIZg4tbLiLnaDkCY5T
GyoTB/N2t0v4NuZwYInXXqMlvxhAqwPIW5EWMr/iFO6DDEmE487coYGGLIRNcw8n
Hnt+URepVo4tJPPLgrILB6v5jxomkZ5tHtGlKh2dHdofbU4wT1UPYK8oqgtN1frW
GiOGyeKk6rbbD0knQsiLWjp6cRpfNa6o5MT6sSyhLm4m7OGweFXy1Tu2qo2Ksx0B
yzSgcbKZvKsDmTBzLHbxTgzCeExaI96XtIZrA2lrCbFW5GKTIdK/iTokWDe2Q1xQ
S1RbtzmWoEl/3qAh9H9Y4ZGcKONHuvuKU5hYP7qWioE6/Y3oy5RHXi9Dbl1qLTv5
OUEuQk5TheS4HXtYUJUHty/k7nu7N7Y62rA8Yo0hqgyy0OZz0L02DgWwiT5KOsOM
fzxMHniQIt5YXIUK8qh7juvVRsRgnIoT5iOj1ss2/R5r00r4hknekTv6hJCWUMJw
HH/rhrJ9S/x7AFx+EYdYACknorvjqWvITP8DeZKWtRXhXyRQWOZtMuesobWSB2Kx
IoHgA3SWdeBT7SgPWVHLqM1noWCnvnYjdIGlEP/ye29Wp9Xk+oIToRTqvja+aZo9
DeV8PQqzoaW94SDFqEBOaAHygxrfI1P5i0UkeAQzztfBIybcZJEEchVlUGIJe6eC
gaxj2ZGIqzbiNY8mxU/+dW20llW2zxT1GxtFZ8JpB88SWVvRU3+IhYAc5SfPE/ju
LQvJ2RZJJQpRncjhWbUBXpmEgzoz2ghCqGlwb5GwyhDiKVlVCL7vEf6niGdOlST9
vBV7brRtrHzeA2Y/i83fiMbml/8Xs/5rNIXexXJsP3jzkocNad6qCR0bivFRcCCP
cQ11WweLsaCocDx46PGM6d6CSlAhMkrkk0JOPFwBQJdM9H6NvV5ODgZn3u7icUSM
KdGzCTUyO+zHVbbVvfe1nJELqjDizX5s+bC62r5L0NM=
`protect END_PROTECTED
