`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CpWmSCS1Tg6GTIK/Y1EjdhjDUGMJQDfHs5iI7Df3Ob57STiTAk+HZ1/ie7jhDudI
z53INdku+Kkn49WEyxvOED72Mx7jNRcLI+unZQnFplyAM7pQYSq4+TPFK4/usJZ7
cPpEBLs8k9qdO6WVLMIzZhXUh++Yv5kHBbiV5lUr2C9bHM4qMMf8aFaP20TGaExO
IrJlXNHGFro7Y5j/eKIg7Le8bcsp+x9xPRYTCwqrE5enC2Alobh7RhrF5vXFRA5a
qJM6L2TGd30YeZr4mBpId28QvlWcXIsj57A6IagAdG37tWdJuTWmmQRz4P3rUH2q
5kwWvOFW+xNzOsEvoBhw6dpvYniPuwp3A8dEY6GSKs1UgcHtSlhOrS2kF90m/VUO
g93Z+AbcICslcVI64mjlnzi/sKQW34Kwl181I4jdBSjer587q2wpVFsHZLftl7yt
zWgROrMRN3oxky+5/fH4SGzw7WhqE1yBabh52xkKbp5V0rzgfr4Qim75zzP7YG7G
UO1TDIZwKtUyPs/VImIURf8ord9xgl9tFKlFrl5CdOhsZxv/SHlpyXQ8k5WMrjXz
j7LshDgsZEXo6xOMvnZdZQ5+H/3UQVzHtcpVdgfK39zgHfKNzYb90UrBE/1mYfuv
iiRS7HbeSlnGdLVVLOS6KJ/ZMpFz5s354wdTK1E63M50ig/s2RAOO1BbZxkA5lJh
bU25h13pmkVEgjaRWZt5xbwkwn+1ERnfowbWA8ZEoM4zZHCBMCkZKEuhVCTzpP0W
ot+1RQ72GPPHPoAXjqV0U9jkidB3T1uHL/aKwIP25mlNnhLgDI5qnA4Hn5+b1rPY
GA3EHXMo/WrXw+LHetdH9PnebQEewAuJiwDE5z7S8LKIVKLfEIbgeGeDK/cB1R9a
cIvKToFe56zf7it4caktEymNMls/rAhln6eff+Fk9HDajW3vZRANU7mEggfR40vI
Y3XrB00MJcnBhgusUOD/pazKYGxRtXbaaYS6jia1Kr34LejWauEGfEZhv3iJwpH/
c85U/EvtQGp/WfApWCUbyr3LiOWgyebygJmRZ3rJkDJWRGr9n8tFsv5Zq34DBqkI
bkKR5sCqXp3j9O3jMscAF4HpACMzAsJo0ygr7BOvuoIVrcRXf72Y8TaYnyOl35vw
VIClbUlccoQcQtN0UyoZvHmsOPQq/M7p1McrRiq2lsbep4mwFlMOabRPL5ItFCh6
aafcSo9NJ1e6R2lvU7IRY+cC6j62u4txI0ciP1ZJz1vmw/Q9qr4f7WFNiZo1lDey
3YRDIGSNUBm8MnI07+s7yY1DpouzZdkO+H4q3oGzTrhms5eA/qDVIN+n6ZusDg4n
1EJh7hHAU4xR3vI7JYwReuAsGGytD9va7u8jdtS0bJkrTPrG6yFI0GvXd91BryFm
Ay52bfgoMFqYZ3d9qS2TLn7qSmczaZudkPPYVmMJsYMJFgFB/WU4XkOXuYaIctFd
tfODnLgXuGXoamGZQqX7rSBP6oGC10BdBw1o76KmrT3hU5PfQt3GOnsomW6dCxgu
LN+k+jTYAd6EEPrfraXIThwyPHhlXhQP0tZlUbLCMOX6xdHV2epLiu98vPjTWtEY
fMHMbihWCDXJW48kJOxRE2snHIssvUXLTTKX2M+hdBzCcueuSv9mtpyiGTVq6Qfs
DdBZCczJWCSGc2HQ4a5skWTVwQFQrl5MioHnmfpXv/CDWLQx+E2LtCyPHsQmdr7N
N9UEgpOMbHlmWu5kQCbGZdsKEmja3pQZg6yxAj79If4+JyjPLPxPaPYaSI5vNSCA
qGU5mibqRU2yt+do7jgZVFAXw6BRu4ZTGuj2Zrv8q9GE1fK6mqDEd7If6bVTZSIh
Nth1RdeWflsRp9Qrom/3xu+aiU/s5QRlAJhqZNaOcGQwArUpCW1xYD8IH99HkDuc
+LgrRILVAo5Z2zCC2Ku2kAWWMj9YN6VdVCj/7RBZNlqCUIY2UbdgGuDM1bgZ0PUX
HTr43IQ5TFxSTcttnfHMWRjFy5pLA+JlFwu5IovH148sr85mo1yq8zYMU3eLCHzY
7glSLGRh38rAaVdVYuP1E+tgwY2xzXXk53uE/XO+UMA9HKJ7pBoID8/G202X2Fni
fWhawN4Bdujs4H7IyB0PV80fv/rH2xQ0WD/BirrUsqz8yS6faE7oy6y2TLqVAAe5
lH9xZCBiLSoep9ZGgl+Lmn7pwAYpaie/JliPcBm42w2ppG3zJ5mtpDz23HzmKmuN
4QB54uNPt/VC4GP/jxcsDyDoFSAjmm78KgPxCKudRdjmYaQ1hygNSr84aDBPANPh
UVmfEUBmjjEFJlZ9IyvdPcgk37KJ/FYrEjrW1xZnbq0FgmNAiLd/NVdkDgHuqxEg
8WR15AB1Dd9ta8NAZSURx8DtZ9AUtUY42mTy+Gbc/le5lLJS/HeqAd9HSblVvS00
Fm2IuVgxqX2hF9cyBpkWad6A4Tm+36oT9JBm+Jl9tO+AOtQb/tYb9q9pk4zqqn1N
dtVoqncmU2wmdMgk7FPkFpM3mcGBATgcMaALDC8/s+ThBM8M7m31ActE1lZsNxac
OZexdCAYYt923FXdhwuO7tzqosvwhoiIlxp7xPi7PIC3B52SGPZvNewlMVRLH+nR
2+zdWBdYxgLBhoiZXXSNiatK67F2Bw0d/KebmZGzEQ8UE/lrHfzEjPLAoOsb/gXP
YVXMz5f/oiXFOTEdt82bDTtd5KvRFcYfojhnRr/nz1TUq09L0kKDFZUdbP94Z8Jv
a779uayvDCG4qd4kxLEsqyX2Wd0jaGPWtEI8kkURs5kSaue7YiVZ537W8E7TRkoI
nxf+zWN2iAQvS3+rvS20Ifn48lzjsoeQpregRyQMCdJzzxRClipgi0U/wgDsG0Kh
eVwWs3CQhi1B5ONYy1sqHANigxIWF2Nko+w7SBrkjReoEmuiWNXxRfiRC+o+f7xE
1GBmHG/xV11tvXXsZvpVVkmICcKsaUZqrjUDyrddLMgatq8LgArJIB9ExQ9lS5GB
JYziTr0fXKxK7cXEFVyxp7AgWTYTDXCx5Rfx0vNDk4NKDIfu0N2FeneFUfYxSsEK
hBVW7p3APgmpC9uzvvt+B6U1NHM3upz5ryHvkNMBgbA4iHPBw+sCY1tYHs92ATL4
QwhPUCKD4VV/t90Ez6ndNALkxt3CWkTfCPPTJhGSUaYMULhi7cuEACazuIphBwpC
eVtqa9G/wXckxvDbPVY3LpUE1CFGXRbRFRqwJ23izLwvrj8TaD633jnC7IPVQZvw
RSZjBw7vkd+9170YWXdcgn6hHgzE1e7F5X4YkqEzuf1bT83GltbLPDAY3ogMRb85
NP09kRMPEsDxsSXvcUv3Czys5T1nos7I3FLmEXYKCEVeo7OkmfBCswQ6YrRaXe08
qmOVhqfU+ApX18UdJ2OHru57mLxx17ojpGLTU8ANM4MMiGHhhPf3uYt/5r8yTfHC
pQP8351GkGEAB8JjjHu93MqnMVhIOYBL3gtlY620OR3ED8wM+0z++yUxFzz/bWsE
n6iO3jXeBcoW3nrHck9diSN6QsCzjw88q/VWFCny3/eWlgCSiO4WhCPfnM8VNn2k
nXK2UuTYtp3Ag8njJ6XRpdcPiaqfGsMRLX8/So0PJJ92v2A9gK2BkFdhiaehGwnG
SAjI7HXr7Ku/JsA/OOudR+WBfB7MtlV+UC8OaqhW6iQhehE5/zEIqvr+4hcVjFma
G4FuBxaWkH2RxNAzZIOAADbX1jaHbQc+hzrhTw4PVfDuBK1E4IvAfe9OKkS4NkKo
8Ft9ajfnoPTEswAhkzQ/VtbCCIBsh9IPKDcdfSMIJkkAJd39XBYRZntfpkzEgonw
QwABabqfrB4xgdagGReeD1Rz+Pnk0dJMmVGDbDC3j26EjFifV+XyPkafAy9Jv+L1
t2hCSs2LIPAUqt1gMTY00St/nTi5Nkun1deZZ68Lt/MGtZB5ExVuSeDPdnH4q4JJ
GqB06L3XTW32UWaaPolAtiwwDFOSZ66hDWvEGGingoeDcp5rivCre4mp3dmRlYtD
tcyY4lvbWi4HJnI0oJX6HM2G1z6Q8IQTA1hMnqBOIlIeNjK+dkGtDaUxNo8hy1Pa
uCxBOZEk+o02E3+ZrypMUNPS1+mfNFDzmMzDaYO3aJRQ4KB/OKwE9NV6b9WK/K30
nuw3Y8YVQK55dN5ffwVHTahkySm5bXuI4lWGsPpAllTiXu3G5qiV0LZOHjiBUVRP
5HO/ef+fiq6+Y8tXlk7UTw+GXEqlZdOfHPPj5imdpDPJUSc/yPtq5vnQGcX7gBFy
HFlZ8U5ya7+WDkHmyMBqAmdzFyJsMI2fjNLJlrys2rfAvwJ0Ej0GpWB9wMCgK8mA
u43B8wi87RW4uY7/YXG5pFicJWqgEbwpno+W6wiqN4+xrfOmBIJfVUweRf12KUcj
VdXqClJfjNYOBlxe48PoVgPmsq8p16vlJY1eHOL6XdYvIZHzrLZI8yjsmMRc7UUo
7UIfOvXmSWyy6gIBp/V0LTcAMYNAV3+/4Qb7kMj33aXtLeXZCoix08WjsTaeF49x
aD8fM4qOnNg+BpX4+NtldvhCxn5Dmc2EYGag79Nu5OlVyz1YJ3dN+frGTvr5mDXH
/LSNNtlwQaAFvl9Y0gHwgeV9JkvmP0RcpIyKNz9cyzJL1hawEqAKHD7ffiN9sQ5r
8GD+bA+BcCLa30e9tczy3gNvtTf+9rziFJLbuI6eLdF0dE87yfbzF+lOVuYvVT14
YC1Wy/mHq8lBuZ9CukpakEnBxwkcb4dv+roSN49b/JSBZtKx2ck0+x4Ly5nNauA8
t0VKCgEJNbCyDuPTDTMRLZI6hNSvH9+m1wDVvtlVYmqIQRlqa7fxPy9FWIn1QpmY
OrvDVEfzZ4OMUZxN8mSp3vVMt0E1QG/Nn6asigcG5ammHiMPT4sRM91SAiZtoa/1
ZsNeveGjqPfZfRIh7R+RQ81PliHR7c+/cDqBlg3JwU9H4zbmxiNZdYUP2AbD/VRr
0OgXUTdhOd1RyJoVUSXsOksiOBM/G8c+wbbvgjJ4cMGCVPvyYCL95Mt0J0bZyqx0
FGjB59dzU19SUutXxXJ5gCG+UHvipvZdDzsXK8wwbeWR2A3ZSv6M9YS2u9myOXr0
2Ikz1FHmlfP9I4Rd5TxX2KNy6BufQ+yyhDMSXgJs7iBWy40tkU1Adb3nlp70fxAt
AsqdxlaA8aARjha3/2j2/43ogRBfD80ekT+y9TG3WU2SrnOPz5xtHIa4WExQO9h1
PHz0mLjlrxM4HK7o6Y5ho9H6Wp0sg7/FTVcjN3R/LmpcbQVXNPErfeEW/sxZRaLe
LpgqxjRV2y1wf70awSVx4eOMBtuR0BX50M2rTYIEP3Rip4FYjt6XWAgBsxK+2PP8
DTDW/QHqwSAT37hl+IBN8FMJSg2ILTQKib+IRPDH2v4YUt/PjhfoCuZnOvl72Ffq
YO3+EgaE4TlnRU8PYJQESVRehNKkgnBz3W6aZ+G2KVNEi94pa/AudssQ5JIVOFwf
hiZwjxpvXhsZwNul5UYvVS+d+CVbTOD4S08pd9r0vIY5VimPHOMd2EFyZx99OP3J
IGkuDOBwdsysKF1UN9NzzPYs+bLRvGhshkfH2IUpnq7yg9N8mNrS389mrhUeppKh
MRwTyqMMrJa2D7fIw0MRegZ9yRXaR2riBAWR1znQZfFYRFwzw0J8Fyz203OZvG+O
Cq2ERTExyo7I18i2R0aw4dDN8sPZ6+pfF6rH2IyrqZxRuMnu6qLaiCjcnY87sx8j
8KF7pFzmkxynBFJ26Q3XGXnMl50GKt/fzlKttqPhABxYU7wmex+Ujn+y8GYtN5lz
JQe31Fk5SLZ2BgTvuEe9/SKpS6jt3OjMPY1kWTr2DFtnUqPeFupjsIhTf+J5xgLQ
wejwDiubwN0IQkZGx3tGdcn0WE2ydnaK51r1HlM1eRgB2oIVG0eN3x+4Zpw6cta1
UWu7TSWAO0cnpyoFFmNX2K+SvakOiwiuvPHfkNXHRYATl0oyMIL8UTFJBFvxugm/
2eLupk0jn+k1ElLm1QZ0osAiNUv3urBIqQFz6WH8wplAqzM97IWtB5u39iTtXzM9
JGx/bPuJmVz2bCglGjcg6yLjVDuhJOf7xMby57wx49AAHw1l5zlu6gOLDTSuABgL
HWR2m5LXsTeQ1NC9Ca/cHE7qzkfnsYQfK3y6m92kqBiNUCda+jxIWWLnX17dHZgv
CmPzx29yTlPUk+XB7rIVJW0gvR5/fkcA2IzZXm4P7obZY+KcxCAtRgj1cFa9txRC
yEukjJP8AUA3C3gz7Ouw2dzDB3mSxzpuyQK+6+8izpDcRik+TINNT1h5ICssZ+QW
xuYyMQgSc5lzX7aUmarjUcsQw/fYskNE/6H6auVOja/s/DOWWYbTi70R6PIO5ahs
ZjNMCMEZUpJbOaJADnm6RexlmUo0jg/IqVBFzV3s25WDaBO46vfFr37QanGmyhWj
5zCCrib0UH6xmyRfTIdxHGYuD4/eh9KZPBFXKmDTFMRgaVevlEYhqHD9DX3imIiO
WUoLCmDlOYWHpNO+JdmLRxVN9r2RCQ6iFVN1qNpRLQes0NB4DwVU63uctn6FQDmh
EbJnngdcnPIAhqP5DBU10vi/w0QKwjEE/c25EUjrMPnZnLZtTQgDNm7tiJzMDj0G
Mmc2vYhxpOH7cbZ7KY95gPrBOsQhmfiVqDB6nBaMYx7ak7hDT6HJzi45PuBKvwF5
j3lO58qM2JYl7+hgOX5p/wIBPY736XU2DrEB+2+fZNE5idbhC0WuvrTrRm/wwPJP
CtPTXIy9C/CjV85ASM5zTZXQca8t3ne3nTXzNipnlPfv+p8W6EESpDwp2VlBXFkw
TvH4mBvq9lJLMKHcSwyfCEt+urwPWVf4DdlpMdIYdEo66C+CyAHW6WalgDjgO7Yg
SOrP8YmIhZAo0dgDaLlUEadKNFKHva/ux5XUsZBHc/bHQynD0vQ6umfnlI6UnFGF
6icVFGu2t5RP/K3ISGNNsMiQ/mKjL7FdGZE3UxnG/aAL2r1hRbCG827DYjRqOeVx
Iu8xE9KVz+C9Du1Ci7slwRazcKlC6DEPczPvGzihiFHyWMHw5LJ/HuwKzfHNeMJ/
rMh/xjdkAn6zb+BYIph74ZtY0OO8xzzjp6NTWTjNb9OjKViZxqZIwnBxqZXHtPV9
no4jHMsqW6NmWZsll91FxRumVlbgU4YLvTsXjsVSqUwBtUc8C6gylIqkDE+WNczs
WUMhz3T2B2wznpVmgHXWCinooWQOQq6Ajxt2RICVGqhDrEF0PfpeZn1yoShUbIRC
/IOZHP56xFwOxQ6WRCck5M1+Mc4+K8EuE0knNVuPcdf4KYIiWkWii/fMtph73Ok1
d/WLFYpXJvrvJHoqVXZvMmVV9BuFEaE+wNYZGUYJCgJ8TTkcR0e7yDKNujRhHHql
9KVmt6F9kziub9GHZq6jKdN0R3Ag6nzUqJ5L/VLYC1D8TMazALYMT3vGJkbTEm1J
6yW9DfsTB522kFwMy8yZdQnEQDKay3xJS6SPw9OvftkNHfyonLydzs/0X5/qOIZf
c8y/HKh7mYULVrUpPIRV+stJChoS5Ow4un0iKf4VncZsouXgw+R7Dgc466KWAHjS
ppETtSTqfsIaBGMSMkgTlW9VHa97eRFJsfBUM8ZhbpYUUamXkf1Zfu7CtbCGjWrq
UyHvrmwYsXZmmY2GlUp+y5dC9DAqZkX6z4U65l7nAZw3zIx/m/AyNUzOR7BoXBB5
uOpAa8k9Zgtx21DUV4l492nFnm0Fha2YgNX+Bz/ygJvFTJdzbT2o1IoSTYtg1gvm
iVBvlyeCNLOnwWVoyOEStGQf4/BECZxF4lrziLX9ik/0fnPpgdX1SVHX1eP578hs
GZAfAb8o8djYcw8xoeyMzCeTN/85KO2nU5CS7zNYhCw4DrRTWmrUCR0EDj223iJc
eoebQ+4QPuouRj6Aj8vb0CcBNFkzkuL41ug0eztev9yb/5g5p84hp6t83RsfRHWN
HY/9VojGCp6cdn0ZgIvTsPGRuLw+mn8QzRRKrMmkAOMW48KcYfjCcZwGbQutMQZE
P9BCljGILUWDg0VE/etTIYyaCSTOL7x8+xcNK8BtGYOjrGfhK/0wticTRR9kZxzl
SSwvbAOvtw7uGczEk1nNfI9cGKFcOejeo+7YdRsB90QztX1KVr1KcOlMrw7m5Jpc
dpIvRADoFD8hmbLIcK8XwW22lgA/Fztzknd5r0r2+u3XtWcECuwZuOMPu1rmupIE
dvytzMxZw7uTfn2g5YZ24x8EvF0TtQBTO+U1XL9h2n+X4HHmrRTMiqbIIlopj0W9
Eoli/AWqLiVtni8NewNHrUUSyWvWFVDZfvggmD/opH9EAfi9XQ5BE5dB7ojdA8xQ
V8nS/RaQZPglDruTI4Nw3uLKRqIn0igO89kHk0A6HkJD2VCXdmh8Ql7miHYPY6+6
uSfquco0iMrHi035TuuDg03YMQvF1fvLVVTkZ/con4yZ0c22zwFUeqGgoUXD32Rn
2Xx0hp00uJRMUWhGMy64I4161Q+0GzfAhF9dk4/pJmimG+5DF6jWZbWBYfajSSfi
Nl9ucBNelHUSCWsWRLlFXsM2RgMCMOePY0Q0YuRduQlv2hO2Zu0au9Fl61RuiJSl
zJRIie/yJabF9vTV++ObXYYjzAsnQOq4dmiGiNRcnnuH6tpamP63CaUWbbpqqnjp
VaHf4VBXqf5Kw7XLNDVbihHN5GuR0gKoySM38r4NzjOWm87lpcUKVvDvaROFX1eW
hnNPjhK/OB/s/t+x8R0bqoPQb44dogySpXC4H/Z/jm18mU9Y5DqE4S5zXV63S7n1
9zG9n9UpsgfucJP76KRWjfbbZ9ouCoA9PImdsttFIs60F5D6xot7xYfijUVpGawI
0rSFknjsDNQOQVWJVffZ97TzVvu959kZHr0FV6GtAYFP2RZkr+Rk6HcJcWnf4XRs
ezMhzBPGnKyWG5mRTS+eGoc8mZPuC9/nsPaGPn0Y3c6PPvWIONG89OxcD+vsW3AG
+y4IzPSTfSMHhzh88abVKah7bqLTVUQ/PxmUNavQBJhisSQUyFqTNZQvX5XWQocN
VwxQ6Sj8z4SL4i3b6P9jA1Jsx0OiC+Ug4rXjw2KDnBY4i9Pu4t3CbKr9LctmjptI
3euo9uQEMqEs1Rsg5+0cLxnrpaA8RWBqCQZ4oJF8yWxAZ9jKrcWKrudXJkQjxY+7
iHFY9caid9SOdT7ZFR+ugo8ih9Y+YcI1SMrj87bnbAchSCZsEjir984Bc6RFXOgz
rb4uFiKUe4WCcw7PGShYCFtyA7t3h0hNWUjEULeCZ0aJtZE0rLYUpx3dv2c3iu9D
UYKaSQeT1mSJ7U6ProNtMRvioLFAThr6+3ww3bsH+GVeQBpjmlhRyX2u9rtT8vg/
PoWvKNd/45r6vDFWsZX6/TxUBWsmkfJHDrdtvn7Yz2PUPoxnj71yDjb5z4Ppu7yU
JSTSyDXcbNSDCPqhf0ktx8COAwyaA4pxdqNLMMAuuAsavGrrmYMqkLAhoK35iWka
ovILxJeoAYghfRdp9trFO7uo4MYmPjTxqOftMtkVloVj+KPtCknbl94SWHwE08pe
Ii5Zui6mn3R4oYOQ5h/T7OyJ1JkugTkM1bD3cMTzXjAbaGKxlT/YKVFhC2QVsICO
OEIjvckM+Fxf4nP97y1WXc3EcUucg8rZ7Y8Jsk36Rx3146AO1LBL4NDJVPQ5+Xyt
bzvvDRTfcCp0QzflFiuF0kcLngae4vSHdjBfR7px78hJWx4FPc3Hkzv3KEhmL6nO
G+bfZt813xFvHFVMEg1PKmwwQ/P0j7rEit+1+bunFkj4xSZEyZlSrB/XtWIwStGR
Tilq8N7yIkr/oYhGXWYCRoCAa0e99xQy9sjzzQ6yPF2MYD+96V2KnlKN0awObs2i
X5wz9mbgDeDGuZgST2QvblQFNOrhUQ3NxvxRI0u+k0poGKsqTw4oarWnb4x2F7p+
iFeFz2zx6UJonEd3tXlmRCoqKJGjbMjZoyaWyXrLVVCmi2vBonh2k188OdqbEn4i
Aeysh64yD+ojUHChFSNv1GpLEyvio6BMEBbaaU+4Odqun+04+U5FA1NC8VksPgvJ
uiBhQUj4nwNrXLDFvj2M2nQu/MYM9qPrs6vHShxNZD1e9Xx4u647JJWTpJ+8MgK5
cOEwDh3LflYG2v0I59rzv8k33rkQUmIZYNuP9hVQ6JmL4AfdxHcwqg2kcNRIPvk9
+V8mpmvYd7Hr4Ba9N081JSMiKQMhNOv3QTflaLzM+wfz1ZB5ZNBAxgz59E12vRt0
UTJYKAphUoRn+iJPy9JeOi3ks2NCMsW5jJ7t6lLFgheF7x7Z+VzK3U2RSAdDjqLD
/5ESp6gVOTqewkgqegYvT68NxFOLpVqjbwKtedGbWbxigxhWRXnITGNRMC4qhAuM
YrseUl5tqxNuxWYKZxo5jNBII5Y7Y7eyfupzLODIOHw1ZJoEE9MicylBripCtODf
JUKQU7bbOgDQ1aSySLJ8wImMgQSOsz2kh4aRqiMWQkYQIweIH7ZxVdYNotdaXU3A
CCJL0OVhBdZ/thfE/qCTT57W8fhFMP+yRD7XOfAzMh4BknJDgAmrAIGvTfrP7Xkv
j5b9Pk0l9YklXeowpdxQJeIO93WucCA+6fSIto2hOPqQfcq84GYx2VUeilvGzFRc
aZhgwDtBIXF1WDjp6WvEtTXg+kOvs9ccWiMmiY71UtWZxuDmxlbLPG/RmxLAk4I1
9mm3ycIgkKmSzuYNVeWm2XjwNlptQtnc0wR4cZVhvmPPdNpCAFJvwB1MX0x9gOCR
qMr/XGxuQSIsW0EPigOX0whEVnPbZ6bcWrqnTCXGVWIycofiyABKRs0caOYXDp6r
bTaTsI+kZJqrnm5MjS0P2WtRCBHXnAW14/i+MV54LFfy4Cu1m/yovMJNnqZjQi+N
5HajlyWzFPZYp8fLkdGoO8lyArQuQVe+c9gA7BaGoRW/xw387hnuIQfTnYUHj+ig
p441oNisKI8wuEqtXK1yx+iAKGqyRYrQsQcEYTc9hRXoGlKOYtJoT+E0cWNxC8T8
ZqyEH5Au+obhliFGLFCKgsHh6CADGl8oX4fu4BnXkiD78ocht3rlzfpREDLxOSsx
+SCsAfx4ROnkCuY5BGLW+9V7HfpvBi8IA76rFKILkwY+6yQN/JziZvEnt0akkIfF
Q8qnNWDLmEtIcIJr8RPf1AAu+xWKGB0qJa7KjYLqoudtGp7VPeCcpCTdjRsnp2k5
vDkiJOy2+MolyfGbJFMgzl189G7x8Z+xNYi0PhRL1Vq8VSukWUjf9u7VFPaZcTVK
aWmglQLMv1b+qxWiAqBSLqxegcF89mOGKENL3topDqSCHqqMCAB8CZJShhSkc9gb
9HC4TyCX1j5Bscc0BEMkfdwV0DSn0bnb4xfV/PruQLQfUEFAcAvXctFAMSlqWROl
S2cCk6Qecknv/zgy6gJyXbXkBDDlGskwkK4WY9Y8i7O4F3ZprZa65wq+47PecmeU
9AdmyR2DvIbfejUwhwVPXfIZh2hmfFZC7HMjVQGwLXhzl3nzqN7VFFLpGxH+v8Ly
a7FPBbn6P3LGDm3Z9GSoMuHTrGqt0Ll9labD8Hc6rQTNqN6SQO9VnljZycgbgH/Q
UaiNaM50rs2aoLG15yUPuq8qBVX9fsI9bk84DNusn1ieIOKw/zwhynzQ8IqqoN9f
1m/MblJQl3TJczJUpQ8bU5cG5Jk7v7brKYTKZIAjxbAZizHH9p4UsfLIzKXoULnL
0Qz8sFxeHPrMZVa2W/Rwzak0wr0SS8x51h6kM6wFQYgp2sM75ogzFJsyvhZf/yTh
2w1jUNcU+xb0353dsNl9XKE37p7ZItdFtTb6a8oiLK9h/iEFWMx/+2vrYDlpAFhl
9nKzxUa8X+M5mealxvAnXEPRcqB0TxnBD2cCamak3L+j9rryojzmTQPLuQ1Z+Aam
db+T81TzxU8YX7zZMTBxZH6WkFy/aIHZyzVZZy8GO8HGf87BprI24axFKXi+trhT
5QvGfXmY8Tv5370WT7s0CAJapLNk4u4glWVs98KUDodsm+xhiXTKxmy7xvZ2ri3C
3BgUGSeDSR1s443CLqJiv7UZ3RopbUpez0Z8IvwSzwq7N5TGkaIL3mxQQG6BNIZo
wcMtntJaI+93lJbS2d9mBTLODbMBV1eJxwpAc19zGTEVwhcDw9itx8QSI6jQi2lP
6PsRY/ykGBtoukG0X/xO8SueIuSTuBR+tooBsCXhoKReEqwkPkTeCQkfc7t0REI7
eKIa52ixMhBnoPaSGALwmU1fvPQduni3rHV0Bh6knz5j3eLLi+8752livecW2lkJ
cS+rlmnUnzj0cXjm2ZmpobEiTgEe86ZSm8mdLoYrhy87eXRbRFZuBh2Tu7vtu0FD
F97jRLvJnmwUTXjjY/i4TAJrjtx/jJm3lDnajHxROIqmv1ql1R0zqQn8ebzD5Yhe
znF/mIGqhil8ot5NTw2lh0krN55d2TDgjqmpHle+SC3W6USUhIeshkNJJBh2ZTiE
G599T8JXTILjhKHKI6JY9wimfi+0X2I9UjYPH0kI5oe9UJZdlLOaVd6FX5x0PSRN
Cz83/JrMYdcyJF0zVzuu3NUZanMjtnHfx7iL1jMAJveJdScmxB8ZpU8cpQEXY3Ji
UEM0epHMxfgZ5IBjsH3ET5NiY6lkLBEivO7YgMAq3wDxTmEvEvRefI0d5OSqNd+j
Q5YFNuamjELVMrhJYrc+7sILO2HW8xlueMPbMAUlFglQTPojQeNN7ItQ59oTki1K
SxGaj/fB3UUjlIV5oTR82S7s8SMIm5zzf0YWGBXn1Lb4LcMr0rM8GpJnfTZoOCGX
z2putGCZDsz3Yk+EWIiPp4ns2uWe7s0IG9rb4mnTK1MYl7JvZfGLGV6uvNZCLNUb
gH9JErMZMliJQUQ7Dgo5Hw1AAz23DxPz1qBa/8tVEvi5Ig7zenO81vjF/YWx+7DG
Cb6uWKGPjzJbFlp9esBtfEsBA7grQgm2dybHmCoFIhHUIX4wdKeIRngZ8KYYV0gO
+zT0AqonXh80HlNV/RdS1K+abcjpwrwRprLhjBCateU8pCDtVXYpiYxrkVZBc4G2
h512uO8JCIU5012k/PonhKrl9yZe8DnvNVqw4BCAik07O8EoELXrJse5fxHx8Ea0
8DMiXf50guYyduXC3KPVz5e6D23Tl5N2LDPDDkEsA7TM5LcDFi2EpSGICgtQJoCo
+ShXdvakpySscSMvX+u1PsKoBm3xgircAMPV7nFrz6zDbKSwusPKk9K71Rkhe7LJ
Kv2g1paSnPQPsygjl2Zv1u3/AgF2g8ZBALPL0JuBQUZNDOXu6M5hUocdRU/XyQnd
gQYWi5QG96dBR0mdRfwmASl3B9mbQu+IyTE+VUMtoaa4IIB1CCq6FggJzYkfCAZK
P0aEjemExWZa5aKK1ueCzx5qzmrfI5T8RbFJlGBxGreMwG4b05exfSZ5H1uz5Wzt
hiaFG0EAu0PtfdSJ/8CxHzIw5/3YdyrPjyibnKO3HykMy6eA5M6AVsp2h4rzZce2
iOVsRRKWIoEpP9iGRZKVVbZzraBclVvEO2/30cVrVrTkat22n+kdZFCs8pcRBmIb
nt2flctb+sTQmvl2y1oNMCQ7NbdX5BLoMSRxaNR+U7IcX6SNtExsC9d1Dnoo7rhP
Qup+pKomUAsrm65XNPvfT6K1vCtHD3lU4f0B6pGB2LP6mrm8sc0hGgtAe1Q7PWAk
3IzrqDdDDr0qF0A8pC+iDP6jZPgRxZ4O2bhzdb04phnABtYXjgQtc1LOXwymbkhs
lu9ExO64IN9bIQ4+BrVaxj8U0MbuPpxPbX0NRKdc7dv5OAiSexkTBnUo1JkwV/SB
VfaNeh8xEOcfepsJ5G3vbzPLHroHh1GzjFW5VG15pTvrGtMUUJtk4lV8FjTprwhX
DxJdpRwekmO4XB7+LuPQDTkMJETANfcA2PR1KWINRneSx0l6zO4SdMd3COfVScVb
pStahMtXMLcJbuDAaWhqtsP7C0KxWlG8cdJnK6DXEmEQgdQsGmXzQVn5+pT5EU0E
B+q5aoTrODQrf6d3erMVFv3+l027MlieOaEdBhm5SLjzbGxyrDvG+P8aqxlQnwEs
5SNP0umln/YPO09zkRN6o9+PTzAcIgUFTj3qkmepTpugRjUwKyXuxOch5WTwePNG
Xu6YuUK8xZFvqQT0SIrzSvLo0DYLwMIeqRaBaQYOqyTApecEpjSs3D01FV6U+b1n
u5VWMzSo0Th/7HhCLTNv8o0y6k8SItZdHSY2acOHh+i24fmZCFPqyI+jkhVG75lG
cbxQHOVyDFpTPod/TpDs5RjNp9YtsEI+0MBPzJNrAFgpYvJ+chIqcqaXc3+STg+m
fMhflclBhkam5LhO/Bdhj02ei6j5qMkBRZ91zYPftNnsVJaKR4BqJRewxNRSuxHN
IkzAb46AlAEaRx98j809u0Kskylg+Qic+jg6Lp0GAi0mAaCD9nl/SiYXgY4+lDEE
GbUInVhtXPrLohKtw3Taf5mJCqP9anvi3hu86+Yh4BXRGeObk0J2CSH1r8+dgSbG
N5MZiaMMxdAkbR0ZteQ4C2QYeiIBKmeCCI3Oyl9zleBvBctdarMWjwACIcfZg/DS
yU+Ku186a/L9BCQfubQw52K9cBqIVMvIncOJWAuqRWpLaE4Ah2GYDktD5LKMqkvt
vCDcZlTKRofF0JyPGBnHc9Wk+DAf/sZFkSFhnR6LKUV5qTcOmJZfKL7pnIys9N9o
Wf8wprwWI5vq2oyLusrA4AwGuPRwGhqo8n/4inNjRAYiiG6jl1/gzm8FuLb0LYe4
hY7S9zBHd22wCbJMDJ6MNe1uCjliD0dxhXS9z6b2I8nko5LVAzPK6/5p2uKwbmDP
UlnSx1WnylQAfmsYq6clB61pxMpTwv9EwsaxuLJBAu7mEtToXf/br4sdEryhSFbL
kGJOTEigW7VAxp4Q+GxOQM3sy4jhQtAicJsZNg3zOKjn2E/xS/wzJAuB9zyiZ+qN
fPzz+UdpLwOM4h+edUdXakzkwFlkw+fMpYh5blaxyM6SVBIMmaO9dr3DdFJZkjBZ
XTbiHCBz/LrzUzWeOAPVS3TrOWlmMO88CRxOTMh/8tLS7S3YCMaSsgQ5u5WNrA8m
xlLVmp7WBCRq2HiEU1y7Db9+3YDll71lhrmRhYE6UqQ+8BaqTc2MvBQfiv8gjPTp
Xlug8p0mLxZuwN0yuC1wA79QkJ7z3xOkX05jpj4DPSYLCcfS7uAGzhFvSwdpyGFM
QoSE0zCwNPgoAjMPa7j9HB8u94mJCL1yJBqRExQPCN8yAnC6xFf62J5rTLFdFEBu
70K3vNtRyjW69jVsmNgIAS0q8GKfpzrdeOe7obLpx1MJqhCGZanBXQNLsX8jwE4R
+lhSwrWoatTLsgiC+QfuXfY5OWoUAFe7jE7s+9XyFzGezoZDr/c6jjgyqAHjsiBK
0TNmtRlU4hFjLxSjdZ2GX7LIQJ7g/eID25+tP1fe6ccN3Z6feAHpQ+NMOTvNBtXe
l7k/GgWf+Ct1s779i+6bEi1uBtv9C5rXMuTyKrlSXTDix5OrHt5sic0A4PvkMyH/
R3x7v8TvrLcemNcxud2NoxRXsLMgjs9mT7nCZFJJy4TYEmgpYQWyVHh/9nfjCQTg
flH4sVoXY5gNOIGnhsldK1wZQXKTa3hWHLauDbAXnsfdt30lPBZwH/zSigv7smqx
8QuK5N+G8KAkwBYdNqx9d6lp3Slfw6ox1XrZVedo1INOxVPKGcsFEBOeQnelzsK7
OewpXB0M1saOXn/HJAB/4Oe84MqLawlB6WV+VNMmaxr4OKV27f4rbSXZzt/1kWaM
661VVlv32NOXXkV2P1e2YJhVfM7PRMHAGWZWqsXOgA7V+Fh/4Ns9dZTOesJ2SvLU
PMZSDl7eA4XvcSB4Mp31ue5PVpgsHxLCJCYdkRFHulblbSdD20vgOGIcg6xRzqZa
3i7KphyeSaJjOgjwZ+b8NSsnmnZMEYnc13iCcfHOqKRuhb6lPAMbwGM8XhFDbjkM
kP+NjvtpWRLC+V2AVaNnELcQgUccpiUvjhcFPtrSCw10v0HS/Q3QD1uFAlDMI/da
BJasPPdKanS3V8VSmdmRNT/GvGhbZT+8SJiITQAxcPfMsKgYVWyhBlljkOCFtUQp
uLK4vv+KsP7DFlQgdemQ2tYH9TUCpxjTphi1946CZyETGZhxgl5sQc246xiQSqCK
QaagsjnpvLoPLYeb13j8xRIXnDiiUBvBq2V/OeCOrdwQuF9Jzuo2KZFUsloUqEQU
Fs7CW9e9zVyCEYNv5iXGPl1j0I8jcJ586E1E1vid+G8TLNyNpoPVg/lECsaW2OYu
d93AT+nAN5kbMf13hLYZ77r6rI/a/KRM1/7JwiKcSXKKqRcNpa7mkr3FP6GJmJTn
xaAEyr7Hpa/Yh+IPZO/FyG9lWC0y0qLv8SZaaYejXco4+Bj3xhAjZ9TRJQr4Wn1H
xCXNmx9nHyM2rKQ656diRk1hT9U9iK42EGbCckljTy1f91ORaovIX+Uaqko4qaiN
pVZmbbqbe9MvXCraNc/B1uaEtsfqvLEolfKsbkdvuXhLAx295eeRj5yr/jKd9ONu
Bf9ytn7+u3VLpVlknfjupd0JBbeh/5pFgO73mXIpNv4mWC2wrnYsUjOv81+56yr6
w9pOOdv9d7FKFRmkUaH9Bw7j4XyIsVMgzv+KfL/mdbtpkdHs4/Lgt/rVwq7fLvxI
Opk8L4KTp4j08U8nORt8x7az0TdsjQPbFG96wm6sK/G2G203642SE5rolWbic3VH
1Vff4VF7AxJa1kOdsdamkRvaVMaCcvuHtJpvok8Cbvsl399TOiQ7QbfnBW/iawE0
yU5oswEd/ggq800Z+xHexbdvFQXZJedNI7EOMK3JAn/euQWiMtpV+z7cO/5j+Em9
mnTiKGcJ0iSmI//A7iez3TmXBRNVkh+KRW8MM3T96IS9RmEid7kpzq2yBsBOS11Y
z7NOJ37Vtt1HbdEO4YkHNicXSwagqzxbhpfd2szNOve3rjhirJTxylqxKzKcTohw
6DNQ0Ezz3faYw6RX+EbLXCTcFcVAf0FDnKxbh7cBMWPFX/0AqzOP4qg6Zzo7ePiC
Umy9J0mO29wKCaq65Ob7XXG66A0c+0nRMAFX9oPkkuB+dyf+Rr1tjVa9AovxJeqR
UEY/XgFBoss/edFMKO3NXHpwJkakNgWwSf2KbMRdtFU4yuBytSIOa5V+feYQt8q2
rE5RWn+zP97eJ7vYPVCJhYRvyxO/ZfOFbNamd1oW9asTF370QVOeJEylwSSLN7UC
gqmL3fUldICdmEt32jtOpmHNLZA3UC+orfwBSm6U+GIVcxy3t1xeCbJ9fV36CZZ6
qDMfawUssoN1M+a+R/cuyJ2CWb574cd6lxPcjavCUmJMEv51dqLBS82Qy9/F6FKC
J7IpqGUKUkjl+64g4HaoGjlHbbz0YbkFFgJDPy9sn7ZLLaobvpm41i7lb2ceKmFs
iyJO+Ay/+ib0E2h3G5HBWkvn9HpJOKIowh5y+RGRCsVlSpx2+x/D7+lYQaofcrFb
JNyhDAOCWFoKl+m9cz9A0uW8M3uBovDQG8VYj+bprKGwfqTpuTUkkiqM1D6Xq90K
+8zj4CTDRb7tkFnbnz3fuP2zNoROa34sPB7XoaKJigLqs2KRFv9rKS5yKAlPLb7n
c/wzBnUMdGwQY0krzbVI6tXeqK3ukRs+/1IO1LyX/g+Vg8n4zMXtee3xAvRHig7V
3ybzRIwKaU5E1UzW6Z+x1o+J6nBVNGnRrs9YNPZoX6J1a1HE2RhvFmWrqs6IA1Zc
OCcctPXYOkmNsg3O7LDz1syqi/bnaoF49TnLpTux6kWrlmIdnQsf6nQ+9Bx1LtDy
05JTXSfbriX/M2QkyXpHHLFztbrgvIhKrSccyNBHk30HP9sC8k4faKOaSueGm4dP
mTRPJi0eAFCkJeMiy4JKPQq4S324jCs16IBY7bioSNONj2+680Izkpsl1ThE0BRy
luzu4W0fEmU/ex97+4FTO4kNzhNRGihFhupze/rfdTJcc6CB7YgQW/XU5DjBjo+c
2KfmqdNMF4bCbTddwxALkaj5BWgwqDCPyVcQYOhb8S46vXh09pUStSltZFNfsAN/
dsxZwGGiO6xApq9lu9kBFBJ2CN9G3Rf1rTL/pUKQUWyu7k8h/6DlWzS3X3jqnDNI
yrZUMJNtsebVzJGpS24+kHp47oICXFDNEdJhvrZcBrMzZBMOCQDxAvgNvp50TCHs
HZ5KltO/dG+d4/7FHyNEtvE6b/Fd+8p8hTH2VoDefVqiTaKnY+Y8J8Ab2VdszGfR
y2flMETZ4O36O0FGUnlK4a6ZTGF6WQf1KVyJlNc5cjTwHk1EcfGeB87om/LUM7No
4pa+7Bm3xsybkFZlAgPF8+vlN9E2xTVit3IdPqpqy24zcyJyy/gTgC9hnuL316/q
zuE66Rpbmi935w2XdA1a3mARYM3hcBm0pssyCND35sAuzKGenEb6jkAy2OK7YTWV
9j9hIAOQ4lXkMszt4i7wRsL9H426YcEgHiSw9M+mU3Z1Chptp3wcrSgx4Hou9pQp
zZ881PAq8ramH4PUUxBL+2f4tVWuLS3Mb26WWUE0ryPob8VhPjPLWrdx/GRwvaqU
bvZZv8XNhcomaTrvbZZhh//ZdarTIXV0qmLTxjn3UhjP978tWUHLi6zNCWm2K0mx
pcapf5MlSFqsbGfYgoyNFTMapjrIN1a3AXZ9gZkefJbvM1Fc7KT5F33ckGdGNfL4
4kaSSpM5TIUV3WB9TJqH8aGTw1nLRyKsw9k3d6ubBJBkoBy1xnNrWnV0o7DWph8G
pCAk73Zjir1Rb/S5V6ymvDRcphIHRao4D3eHv1iM6TItQgyVvDpLnkSxxSac+VB7
79Q1Zv+ccUHeSRII9eTh7wq+6vLRAUh7a+qKYAyo/iSoSzW9H0JKG64rWCqTK9MH
Xvg+EwnyyVa/mj58IslbF1eoxvYFNvncpCxFbHAChEnO9moT9VPIpEUadbu5SUfQ
ZvIGOS+O3MqxUezR12qt2m98jGiqaVYvi4dJc/k5w+27n61UT/FQ8dYn4cfZ9PyM
u6AZ6wxd2vni4vxNatR2b3a0HantPmGVLkpslmZl+x60wnVT4408bDRx+5KPpsrI
Om303xXF0vDuE7k8grAST5Bhev1qPOoYCF7SyXfX478aOsOImxExEwCh6K/9GpfP
YjqAkccsNirNaxkfHVgAbwCvWSa7Bq4CNp3WxZnLNzO/MiMJhxXmHKz+OXOmsx77
1dGpv+K/ZggZX5MXZz9Em8wjiMJkW1dmCHzAeEohXviKOrgigEMeLqL9avS1JpTv
jH1x09JnbtE6vjNa+MkIuWC4aTssLdwTsj/EdRA+6mRultkeIuMphs4CRke3XpdI
r3j5eU7QJGTU0VwV2MPD1EZQwS3Bp6a/tnziWv4+5levXkYLGnwBrOgpZEC9Uvnm
ZaPa9naDdCIyBKifUftwZYKjjTBWj+dh0lfv/f6jNWafivoruC0ah7Ws4OLWLjFz
WcBNifcn7I9KGZVKiDnu++Ot/TFStrDFkcMvx8WygLd1duM5nIDd7hKxJFJZiV/G
wu/ggYL+Q3CYN+GdCJRL1uABZyh8eJ8TWmLDjCm3Zg06tVXNuwAH0E9eHQfbQFlf
K7o6XoNe4RJYpmSnbJGy8R8SyDVkjy0/LR6X0X9/jOfbn1wqa9yx800i1xN7gMBT
GlQplGULzflgHMbO+l1K7Ynawr7Y7H8YsveEFMTi99Uwt9Z6PyMlbMwhX/s7i44r
3UiZwhSF+6c99GCRutskTDJXsyM7p7dNwhsRudBfAlWrdP+e1z/XoW6xa965HRiE
iCLB2x+JeD5B1glnkmByzb4wp4S40WLzSTIBiWo0kBCg6sZEYq6JNE7Hk7qQula5
2wrj88yUYGu6ffkzY7HDiSQYGjzg7bvlOWl8czYNaNFQ6GH8CYI58lmsGXqPsU6a
pLw3QY63ipoqM5C9qfg+5f3MVNLrfhZ8ZFqOKCbhwhXlSmJLrwgVMUNptturYqFG
U9WddXcX2IQyn1+9aQfxG3zFwmqIJVb6DG97dzlnqxNnHcF5lEiDeECfN7EbP5aX
FbDRUOyYOk0OSEwAQkUDlqHKfCCpqJ0z7S5mhVZU6AYgmEaFXaKJHA+f8RG5BDt4
wyB3RhO3hlTHpw9Hklm2PFlyf0DACQn5PIzEMT7/CIrm317dDqPfR5O33NgbFaZ3
GlgMQxQQG5+tyDkQZI2h0SBD+Dz94N2hho+EWOKlHgliEQ/FpxBDkNwVn61i971B
MKoz9r3joaIPRQIrsTPLRb194RxELNklMA4J6ZyaQwBUwNoWTmuhbHlOGPahFvNq
gcXtlXwxxe/xA5ER/cDRrqFmj6DuSYtY6LefJ9TvqoHOIr0U47QN9Bksb3Wpcszy
7zfjns7PHxy6ONZ+1tnqq5s4KX4avO6rKI3U2NGjIe4U5UhuGfSoYiQJ7HNGISc+
6NV/WFNwsvkFN+l/+sUm8K9JMEgiTFdUnTA48wRhlhw6bIlpcLO47yB0n3r1cisS
02guuemxbh5b++LZh8s0q/d5G1uAlH/XAT4sXfKW/8nw/K926Bt1/UZ2Z1abvgv8
VyBgbuT548f/rZlVsjlVZXE4bW0pyhzuDQVae1QkybbR3k9K6MLgB/Oe+FVfkzoJ
aZCttKkySwjDTln/xUPvTr251xbQXDEj+ZzUOtE1ujSlIHYyNBoKDY/sjukID5Ko
QDYs6VlDi8ibHpNpZCZ7gAMcUiC+8xRfb0UndHRrxhVYHgSDmsnvqnvs16UI3Emz
IEWMHtlQwCHQGzLdNsJUfnjWFVqDyz6ZYrql7OCzqHxNQd7vqvJdnvbvftREagas
V+migIxc5tQ/zDFUyyHAkrxS/sZEm8WQk8+oa3qOfIQ/v5y6Hc9eyzzY5G8HsgU6
rP10+zBQqJhTIxMMetTg/q6npevV1Pi3lfLhjpl9TycI7NGvmDxP4BBCcpSIUdxD
SLr69VlltfcAAqy9vPS6bRFNu/00piG7IAIxZZHfCLMnMkAJTjEE2r+FWkp6QmsJ
C2/aD4fYqHeNp9ejQFBNFn5iiFx8p50/3LL5vi1tK5CZPVuxk9w13mHCpEbtHGdD
qzcIHkqc1RNeKsHoKEB8B+5DVGrhaUFCXh/pYG8zG+sp2y2XM4f6Nw6JlmN7OpB6
wTfuA6USvZJyKtMkuRGz/JrYB6V8CN82ONccd1VCn99rYDKSBmdij7wQLZTcVUJt
h47R70gOvt025TXa0X/i8gHOykiOPSC43U2VhGAc7wzUlH4m5OQ6xWg+pbtY7U6X
g3MDlySNV561tGP4UZRMKT/lXoBltimv40IB4RnZbsFkka2sLaAUh+bDFDivpvUs
6dzd85kDPUSEmBgjsvDHtohHKAoQiN+UpoaAf0hexv9nhfKt78jc4K8v2+IEJ3WT
5HsIFWFkUnwVzRBP37Vo01d7pS0jTFiSjKdyP/4o0lCitNjlrw4eGpfsoiNmBh/w
crXlSXvcZk3KREgGghRvadP6fZ5hAdloezbr+g9OaH6VN6ZOUdqxwHZYg5cOwukb
aghlmACego6v7cqpMtGz4co2C2vXYYdqhY5R1XNZ0qz/kKfey5NtWt6k1+Zh9DEN
MO8cEnU2ZI4QNi9fIMEUXODHqSFkRDyU6pwdHRzlySku0IcP5S5D4G1etD3kTC3+
5Qa7lDuv+oRXNCjsyUfSzoDkZUge+KyYIwHnG7qIFYdlksHjW9TpVpGC/rADobqr
KVrtpROF3chVvgzM6S/fCnsai8AAhOCxNI8iuAQMiwGZlN/VnZKMyWTHPqmfTnDj
lz88CP8WUkaXCOFVhpT7+kYYdG18MgbWGuQ7a2aYZtdGLgaKfc8t8fh+n0aHgHJP
d/+33KdiASxoZUxiLZIHNXrJhHTO1jHNigAd2ZxsvtwsmEyq2+PHZPGnoIEU4MQo
kO54XMYcpGYi2vklAY2FUXDvI7pX9hXPNyMx2H0ZyWLKeRz6oHuY0UO+uWyqh68B
/WW+bd2IZTUEua6xm1Q8oZlvxZM24Xx1VH+ilxLnsG4Q5uI50dZndUgB97lExsyq
ZoMQUt38A9XkvWNgLfXc0bqVvCB5Y3BX8mM+HKsKiAw6piJIrsnGunzU8869sM/v
1D4zojx8J0cqZB6brBVU9+4vsqqrRW8YY4ujobSYxC8xg8Eb2T5DdKdqmGvRnhzc
SYG/N13uvGSpUrZAbEyif12zR+s+2mwxAkfzPCl7UOAc40MAoRVD1cPwbnSvAhcM
c13ux6Zzic2PfXrCmZbS/WsFIjhRvItbcQBTvM9lIYkOo50jyIYRKyv0zsHBw5eI
fcPCckGgAH8Z5s5keZYiR8Z1F7qIV1aqtSmpsSfdcY8Qvm3wAlkpcCzxtSEZzvhd
WwAo100hgdcr0fUSRm5oc2bDSflZ0pxnmGZq04TL52CmcQb7Vm9xxmrE7ljXNh1s
r9vZfCMzyLYJcKm1VajEVwElVcdwfl5FG+af/ZjN+r9IcCpNKyyEm5LZg+zKRH3Z
C2RSFk5F8Zk+9BjBZmeXGb1SVuSvQF9xMArrlqHjrXyiQojOp7RRE/MU9fg3MDgp
SCLNKBCzOaKasxY6FMoAuQIw8Sp9B8quIRU2M1iLW7WpQJmclDb9Ikp/gP8DAhZD
g02ZxxxgLQeqgBLRKvfA8RI23owxs2yVpe1HVfWvCOXRXmc2rrixCkcG0Yc0b4CM
nDOMPRNfpFoclmtJIflBl10F36T1cBu2WlSQkZ44h9qK+QRjSY1HyDLlTXSgXui5
5itBtCKEF7imrA/l0m/11PcYHPhiPMaMulhGKQRQ7lL55Y1pKlNM4tBRNpevIhkN
zANdvC3SMHUG6yOKx2UqOY0LM2WrRkMsbAHb59LJY60r7QqlpVXblJ/ZHZkcxwrZ
coYVPv2nfmJ5bkbGrrsFg55vQ4julIC8wl4cGRYccm7A+lo50v+7fnLZe5LN973n
QuTYiwV/FCp5/vUAm48NVDc+8xe7KcDzaNr2xU0giMVGeLLc4RTQS3zji/UBlnOq
iiJumDPyyRqSIxOr45btzN2I7/A5ZieJ/46prUdoMYPtMZGFa3+I+FAfAMWvaZ30
/lxBHTfHn0Jv2AMsCAS15pAzujTCOxtkY2uZELqfEvd6AWjUfQTexJ1VdzjaBRrO
xG4lmCPGpO3a64zveOyyQqQCwwtePwl7/+h1MdIQe91Ca5k3OwviPTVM7SyrTLeD
d9Zx1bS1EzoX0pCauIicTQqb0a0rn0sSzCKCDnWqcNPFWthb7OlKZyBqYWnbBJdC
HPxsT9aBPd3vxQ7HmEX+Q8b0G2/dAIZnE/LnUewQ6agfhLjXiN+KtrKM2oMLVq0l
6pv8Al/XswWW+ThvlmpVHvulaYv5Oa7xHL9Fz9Qtpo4S2IZpO7K0itce+5xdeKql
pisaWAYRy0hhXBVCmz60U3XONX4Hubtk/usCZ/EPvnLJUh/wbmU9X1fGnkiifkBh
ZzQAShuGbAhBBkroUSXIQC1RMBr2h8mp1oYYXzGXJe7IJn0mNL0PohgHVQWhmWF9
H8/SHZMbpGZQtTAFktkur4m3ySYmwHq+VYqv2PVvxAEU+8KvIqRuqDkN1A+iTAKp
+KOHTsAZWYdANr9F/wib5QibPY83LSJpzz4tueymS/J5BWwhmKx2W6tHE0to6R8s
N4npYfArJBcQppO7PBfrRIx65aBD56udbQSH9BccUZgzEyby96ruBjJqqBMnIaGe
vl1uTl+hIe1OgHxTBQ5cWSsGr0BhOL4Xx0GGoWNUfCjP0wE0M5WGFKdddCc74bd4
WGrKs2FtB3rZp606tWyGhyr+nDQG+5Zq/Z5gdbFIAjo04+AheiG1xi4M11FYwfTt
6W+qpfLPPUcoP940eZLZzs2b+hd25XwyRuDOqCk4Jx9Gc5gjBPY3j1k9a8Vr9buY
8YBB0ThZTnzWgYDSc83wXCIjh5QfxsHkfui0YgH2QYNKPHp3UguHGK63bHdZt+iJ
PW3/MlaUdsCtv7PMvpRfX7zxKlnFZhn4Ia+bnRnjJz7B/wViquSSZHMr/wshlAPy
HEtqKRq/t19xCX3olc8PUtBGwDARBXhPi8NDJsqtAWSPPbleps0jRgxCpMQ1hPyu
JPJ/vWpKVoyYMKsL/q/9TazeRAJleFA9GHTWiXfAycbn/5dUiLF85vEgNOwoZ+E0
MQvZ48/+DV8r6LVgJady9jNK6qdwAO0SHTkCdpE6cGsZyX++eg6xQZIjFMk+SZCL
8oRzRRusRMugGYHax+HeXTXRh6VFE5exl4xVdl/xoZKpB3Pp91Lmc8ODuHvBuQUa
+N649lFOwH/Q4gNFnWh1Jht42PkqIBOmZ7oDDXiiAXIIvyWea8B2x58wPa4/JfXl
lDFTRuDcSSypfMXnNJKzr6HlCzkJKaxPkGRuPW9lY5e/X0ca5957Ec1fhfr2Is9D
taOsAtH93iMp3q2SFkgEbjf0DikoSZd0qGDFIc7yolgTbsdvgF+crAo8XZIxfdlF
qzSZAyph0tVXBMXieUSJF1deZdncQxMgWeBVBTtMjihdsjpY5xd1IcqwqlEC79QP
Fa3Pybf/CMu2uiodb4TCboe/bbAVDdS6Q+5oQjF2smdieUMf6gUXC66RjsCKjAgR
5Ixh7vNiso6tXzFzF0hRHszlzyi2h9kEeMR1lTXyTaoCUL2Fg0HW6RkhWdlZ/ErO
cGHn1jHLeJSWbMw2/cgp1L4tnW1s7j9fFIgyJ8tWwgFK9Agy/sH4/VYCkD4CzVHg
HA6ON47xGQQdXEMqw7yflRTPozVsCQMLGQujjwWnT/oU9Dx/ZQPD5HVE/ovuQTpn
sn00K0eYuOLjHmYBBjtTZ3wHglbXgEgV3GEx0I5pPSDdIjtMtDQbmiGN94fDbdK5
NoYWFo1Vnaz3XmrgcTpGiyda8STGBYTiONPhfhNW4H1hHyh0LcyrwikppHLFFvS5
pv33S726z+U4qSoEdhLT1pbpDgDauBCMGzK/GBABWsdsjscxZppNyBns4HgrQg9b
x2irg8Bk6hBGpbX8mLIic/17YTObZHmS4ro+W5jKj0XYtB7CQJzIRgyb/n7Y5BKX
JPLZeE6JVeTiFbbejfW+yZM4cCbZmqb9QyVNBHed8FkX7O9xDJomX4v6eIOLrDAK
uecACqYCxelRt1q5NoytG0eMIeWdwdqsU+FILGrHxtdIrZrl3RYxq2LA3ev3oRK/
jkt6sf+mAAusZY4x6sqd1sRWySZ+f3VsFwkyORQo8BPI6oHkkNybYRb1k2QAVuvT
JQkH7Vo4wZk0P8pzhVODCoU4XOI5590rEdoJ9HHuTKEWacm5JmR7EcpSFnvVOXnl
kXudpeHmQ29xDYV5zxddxUNZ6Zgx5yMjci1H5BYwxGErKgttsZW3D9WoJ/uzcJOv
Go/zvz7JcMREn4VFI+ZXJem08ngc/3KsdJ21eXw2cOJgDQHD3ji4XpppF4Fe1/7w
lnV5YHxu/C3FYtL76enu2gk26UC5V7i3UgcwJsnLZOsGvcapJhUzTEz3+HyleeyQ
bwhsxEEX5n/oQG7LPZN0i5/9w3DzYB+7zkdVR9TafBfYuowzcw0fbf8xdcMdaLIR
IeQgzSZpDNm8+Z0gpdSyu/ASWX/zgXQ/QWVAMhbBavc7pUZErfMdY/sJa9CxZupf
OzW33Bdw/9c8NoLc1/7N/ShADGd1AYCxhWtZkL7abb3nmP7FXCd1UWJ3vCJYT2eA
qQRYdwFKboLe01jcU/3IGJfXowTDPejHr46zDAqzEe6/XARF3K87E+p+dd/qYMHL
znnZjpyA8zb7L5hGfKiXJNELnoWgIzBqV1OriKFWoWZ+19eyMAoo4ePTBV4msJEl
mL1Y3P68ryGYTaLnLIwGCTjv8MghIBtFXnH2LtnPlXjnByHMmEDV5ESidlmvSdjg
L5GZ+MG8RMbWbagpUmcCukHZXReR1F7Hfd8T1opOHp+Q934W+pOyNEmRkwnmliS2
skDVlcWzooqdzRKoheErJcT03HvKuFeS9sveIAGQUjdtroNrFy/+VSvuNu25csVo
y7ptzekVT3fPD9HPFAcRekUo6yXU/4sTlU4mhVLLV4sgDYkCM7+COG6kUSMrhRJq
24ohxCpwoB7bxLv4uMWMNX24RnXa6wrzi3z/XRVScu36iynUGtoINUnllLi17o3m
vAss5qGvPMjz1jJBRMYWf80r88QG5JpbWDq4l1bBmLbDvluYw4fGdxJtiB9/CMLw
UTtKM7nxTKMtcXazc26a/8s+X5++yO5bwXxdOFzk5AgCwoHlycxZgNbsRQUgQjfX
CDIqcMV5uhYEVf9BX4Yvmh9tsa8HDZXfS2drtX7EpgEkp9TgppUimfTjc972cT8g
VZzKLrAozaUGRP1WxkmwT26zRTSw/ntuRFl1hQHYAVgc+CDGFgp4eUgePAqrOzAO
h4S78Z4PQ5gllyjKy8Te0v09dGH0H9y5ry4RoqdJ203BhNrXrVSJwa4Yr21bIKYr
+ylUCLfDJ7a/0Jn4sJi6nPLqyjP5bQX+v835FcVre1Ov4ve87TZNW3DR6x7dEEW3
bowttOV/fPiYpr0e6C8HZZEFAWo0lqHUNSV8MNB1HPftFXbbhsNLCcc4bD0NkYzx
DVEzaNiDBtpkz8lxc3Ocal3S+pWWVosnfhTzOe2qO0PXcMT8/CmJ5c8wBR6DX4FQ
3Gz1XtAN809aGP7ErV6NlpuccX+PEoUCZXU/W+0/XxqhAQriwU9HqvUkayJcmXW2
D1qiZ8NJiqH61jWgPl0k0xza5PaIdqdQFVWdC3K2CdsY9x143x0UPs7XiFRy18Qv
I6tY1jWzeaiw3hOWvar+N9vouY8o53HCbb9K0jB/6mdINLkRPQqvY8QenVoDG+k7
+AcQpUj5vyDxpz85COZX+LRQgwsem921X4SKHhog0Zo+g8nYFuh38Unc9kJYSLiI
+tfua/3leqkePpxemSKdd/SHb7BE1c7zHuGoZ+6AXCyA52GJdqJJ8KyT0HA+mIk/
28TkclkU3TXg3QrqXgHhE1rWKzZFtHU+CuDsuS150gYMNBbP6u2lqWNhDrxTOP6I
yYYBybChFWTuFqhj2IZJ0nBQKwIqkAKhz0h3cy5T/SF6X2523puOW2Z636nMMkZ9
GfEUtdaHV6HH/wyXT6x7/P7vnzyjij6O580CZW5PiKpWYuuNNyRCxRzXai8bAXdT
BRndg0RvXKDEMlAP9Fa2513YdEmGKK7ND/jJn77mEGIVZqWRKNMDGWMHkWpO1HDU
Y9gZYz+VBWO4kvQaEFJ7QidP+OkGhFT23pjxjw1yjg9VFag9M9WrHrYX8cpCZNqn
GdPl4/V0nX4ZHwMt1/dgJYuV7RmOe7CQrgYEI2p5ASj44k4kpOsItlZTch3z3+3h
+8lA8uJ9p2zuctLpepSTpTwStEkGjSs+1WJZl7rA55W2kb89SXczJyvr2syKSei0
ANX78HRpo4XIOIQyU4IbWMDBEMi7NFBkz43wrFCpgjTEItSEmDl5IWERRM/TBCEw
0C2+jCkWiJ/jrd+9b3Zt2rJRoQEFoEQuKdI7Pmk/rXSU/peqcAHAvehDEub2xDht
QOs0ckv/7Jo7qH0c6un/ODrvcmHS3suGLEf7Qi4EzqowuKuqi0Eo6kewyLphrbm8
7NNulvrQ+APCzd3Z+zlvA1jZfZQOwKqIAxC8yqJX56P/hIdm72Z3tMDklD4P5HYe
Xq1FfVFmycuI/lAUxF1R4aIuwE8fnLuSzaT5l/9nPeiEKEO5f8G+NXEXQNfUd88T
z+2Ibz2tXe7p11e+036iNxq+SSt+kQ8aoUC9aMcWDG1Uln6UT5Plw32ypUK+MtUH
o8KMNCsIi/CHSucwqeTiUq8cwXQuz0qHc8Z/8MHEQd+wg1pyTmrQwu0fGoguBkyL
+X+Gud5GRmTtY282ls1nHlKiTavwULV/QO71AO3zS669dZp+jem/Xg2fSMj+SpYG
6U6Gy+HdYNdIyIEsPGt2GyD1PIhAf/Gi4GMDmUPlZfAhkiAuZm0nv72WWfpHCN9i
cfscON1XhE8U97J2TdUSmiRSuPYSfG3o2WoXvJFQ/20bVWbt4oIBBYlz3T0nYa7K
8ux7OlCsFKjCN2QI4LG7XzNKV21KeeyHoAZcVHxJYd0YvirlibHW3M4In6xq09oB
JErS6Pc9mfPZ79UxMWcm6Wk35/ffufLHayTy277y8niGoXph7X2iKK0JUzDKJ4RE
16JlCi2pLUO7mc0xN8gedIp12uXgmRX93TDO1aY41ijhXBVu1GdKqRhIl/mlp+Pv
RnQjycaDCB28klsmC7i7Y3WseNebfkbHHToWsQ2U+dmzq0MWj4eSfXsYad42Po4G
WkQrk9Shjot3rrut7TvQLu56dNtJILffkgsfa0ot0gMpbwHHkoshZLhlBpe9lrcd
9KYN1beZqnoG+nSMn0jo+JNpmnIkAZg+vd06Ph2piHA7UtDS1O+ddIaAY9MwaLJ0
DeDBKCW5xTvHp81EWlQFpwMetKQpVUpwLoAEExAxAWHgDVRiW0QriC0RJGSt4Y5W
8FgNyxl4OaHtWygcdgG0u9nsg3YqsYTj2B/wZLMemopdBIbiiVdGk9mrdNtP/KBo
tya1IbbMxKjAlX8T+vfkYL/kjZIhvLvlj2j1VqtNafU0xq4l2Hq9z52sXbnkKfvc
FCz1OuMcqdK0kvAfdRhxwUQuGiHaRdvxiOTTdSl31L6JblRxdaAQIRxoYFyoSRsM
1CV/uKmflNK2sSdiZY30UJwyilKBe3cQwKTKc+cTYf3sPBDFY9vwGOXY+uAgPvV8
CcBBXWnLBqyxK0TTkWE7ofJMwpK9hmdlVU4roEMHaCpQNCxsH6KtGJcERWihnWlM
Ic3EIRhrf1TYyFNy/+Hjnd0yVXEKK431J+ChMSA5/aJX1xt/5hZHZIiOQ5Fd1glR
gWv/x//I6dX9JSQYlRLDz5Ssg9bqweR4Rlsfc9EeHecMlSlDZuY5tDNKMwBOsW1J
hYqdgP9D3S8RhDITodR5FLelH4oYBhq7hAvxjDhSGZ8yu1zB1wct19MC3BJM4PlC
24Hb98KCT3rA1XOlCXZHDJMU28ww9OywJ7CfrSIa6IISK9ji7JAKjwPUT1L4SIRP
DYColAUmAOmK2C+mItNWyySOe+EbfYVxfjlzNZWpVp43h73jksD09HRw0OeB8pLh
yr8xZytOUyBQcO69hFzYvs7E837fMUBkB7KxKmrTOozyuPea/9+2YiRIPw10VD9G
Hytu52rbzV3gVUI8ZxKW8mmEFfWVv7jyOfujWmfkxS5wYcZFTI7fJxOhIv6OAH2R
k5X009bhBnVhW9Eed2Vzx99LptlVfOSu4KeAf1G6QudkQwslk4bQSXtB+RMT/yZP
R+h6dhN+rRtNIBwNMyXMM8+ZQIYVOsekozAKbcK+HCxVPIwbEo71zABUrFGTmHUK
+vcdbwLHxQPMZf1YyvD0P9Hvw1bYpxU31ZnX9ksvxWO+JGSYcxjn4YW9GW4aF2ty
9AX+9axcTDWp3IKcBj2C7CGkmzzyUNL3jgAIzK2yvSL29+eZos+yl/IiTiPSVeOL
+u1uc+eeQ8AUGo70OMJ3WH4QCUC/EZUDShqJzNqIVPyPgwXvzPrySDGPgKYRxYHc
8WmGM0FWtjDBOTF8415z0gL6FN58z0A0gBz/6WVj3zuq345BbnsKmwJzFXq8psSq
YUr2EW2l8D8sUAH3a3UTLtz7D1fTW9bfW2ZOe4kXYkAPTW0G4VfZy3KI90R3nwdQ
41fTIH9hIH0pRF0WE0y6MOxRXqeN50yL7Lbz8oaTlggbYbTXR8APPBY4cmIXDM20
DXSEJ/QDsQzxXxL4zW/A8EYkN9mdE1CR6v/b3I4cUahIeR+hPZe8llZvlZLBByQZ
SGRcVuuo5f2xW+Bi5zWItf9Y5cYNLJ5/s93tR56nzPR7icx01Vyj5XCp+f4CPfaG
lPL/cKaE71zatMJo2AdesmliIkBcBCO+o1CxX9tQV/vcAnXCbNCVLdI6c0mxWZSj
Oc5Xl6/rkmiM48ZrJiIGrcRwADWmkLKbvggNtpNUZLjZqnO8kX7suVKAYF4Mt3rA
CJ9wZjZh8d7tXaHXdGvzMyirduJjB4/cmwhG5edk7aXzxT5t8mU78UYoPF8sk02g
SdzWcqPL3V6xXIkCvsB0EUsi3AhfWJ06Qo9cHFaBGQ2/nkiN192I2UMj6d0ZpefB
QIah2z+AwXLl1yS4v2cdUKsmSDWeF6jWsL1yi/on3bMu+lNuCJDB+y7DqtucCjez
BUZhXWNatbYaVyMyOAVRgE1xU8JsSfHeXrkj+yWKorOPagq+AbgQFmDiC0wdj3wX
pp/3/3qnFNsTe3I1I5ZjbsZJP7RqxA5rAS/conCs8xI6ym3j8ehidOIf8klyqige
xqVHxSxaLKxp1tZYRlZvPeLtq5/ewp9YStsoGB9h+lCk5NstbOsYYC0AzfoaLGH5
fdJQkEvYfU1h3L7G3SNP0ZYwC1F9ZD9C1vTM4izSRQFoiM9k+SwVbz9cAEIUQsjc
8r+nNogarS/4BnKaSqb2+hd1Pb0EttWr7HFjVUmZc6nqrbPxsYMZmuxE53ef1Yxs
VL+aranSzZQ10MhHQSk/AvuC8HtmD2NfFkRUIqFUVZM1rjd69E6ySKJhIuCkgrY7
D2Dlv4rmjwGrncMUf/U0+gEO2gTeV0pVvq4qfoWoqG961rh32co40u3FABpU8ccV
y3VY0Ki12cZew0gaYBrHV1wxpPC+ua1qTAg56Vcdx548biXfZ5GyS3T6Nklsu/So
G9bIg/YN9/AKAmNe/EnO0+rbqtGjEhmCMA2xfdtH0puWS3Wb7QWirx6JsVro/Htj
gPuzP+CsVDqXvJGA4ujfJ9HddQ1CLTCzMG+j87xvb5pkHZoOKOuKBJBA0iPqabXx
pgfP2ThxnOCs0D9eDTNck4Vy0crrtrQxnuOmncFCOilLcyQkU/vq+8coVc6GuEyt
EzJEmfP0T9oZpfxtKu7c3mq7X0YmJGarHFkPYjQIocc92o/e/QjFUdwGEVO2QHHj
T1f4d2r6YHvssVmf2JSvBPvo0rWpAH5LacS/Y9aSJOgU91MS1A97RMME4/fSQO7C
+e/FgLHruIkmW2tGjPRiAMZYUob6MFL8CuOYQzQGNidPbvblRT/ZfllFO9oeIC33
Nml8N56UOPyJqzhXkFE0k9d8uYLBBAawshAw0kn0i7o3uCXKRdhqrUXRsjtjvdff
ZgmuHADbMoW1Ldwb/Hgr0VpcjewZiJOf1z+cMenGz2BMiAW8mJY3/B9AwHktTvz4
frMrGpdxpRDWInr44gRbQ8FdliWzMhAGQu0xi3KpfDERlh96bCTfpdexKA/b57Jn
C9yvXarE9vpjpCKBhRbIaSsOKQRUSeumdaV+VfPKJs6TtorNKslcDDx3Ro4Gmh9g
vYMwD5BQmGQh4AEK7F3jMi53SKAC417bIvCrXliSvvhQn4aby9twcLiT7fIesENz
ulNkc34ZjJFOtCZ645OQqNji1acnvRecMq7TVR2pdk97g/NVy5dUF4G0aowlxPdb
77qQmXWbn4j8Omgry3n5hgj1mCv3Ac1ezIVrtun2a0B5KIMNtIL+yo73qpH0ckv8
iRQFPTmx+54HyLPhqbk5MkfPmzCowosQ+EXFNqFGoCHmG/Zp1mdggFfl8dj7MszE
yHS5ZzhM8nepCnpHBObIxSpsOczt6LkbWDgCpjfsz7+2v/HJBCs+YAGaby5nAuRZ
2FHZ3TFSeCjvWNDHUSz/TpeDSghCKJUZAkRHirbrV3GunRkADjV23+SCMD1Jm9of
AkHg8yErIDAMr/ttOpknxvt2RoSyhCvcjKhKQdZUe37/EiGpa907JozJWm/1Hes/
GpTYywtPUEu4f2vkAWpfag2uZSDD4bIzCpm+nS7oQTbX5QxTIAd+i+M3qS/YZLgY
0gGfC5bg3Rm2+5GWIyg/qiENaO+AtwRx9Shfb0Yx2iIf64rxOtCutk4yWUQDM+6O
Cb2DkBxRx8KYqKJlCGFPvGuokQAEyjLUWvJn1/s/OYxouEar7rHoxeR2u1sVBB8+
vVppdC4U/zfW5VVuN8S5KY2ggpLzdrJCt9uxRwSxfLMeHJc7ICo5l2XMIoi7uB5k
trfBHQ4WcKiB0tQlAMGoFwJ3Oi5Wd9YSNU9Y7jnn0+8=
`protect END_PROTECTED
