`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4+KBQPwuDEo+XTWDu2tCLYyeJF/NqQu9Bv1B289FxHr6Nbs9TkkYax6+7xAKBpZi
YHua0aprxaFJ3V6OSwF5IPDCYMn9m+1BLqvQXDiYid7AA3w143i6tSIJoOvCZWdq
0JeYQPNFq2YgQXF4hCnGOdqZToaHXmN0kARHD43RTegx1fQGRv6cVYcBgp7d1ded
X7JGRWiHM414UGswW6FDFsd2fiiiStZOk9ae+1dj433CgMWwVYEMdou0e4CdSN62
DV/0DGokGlZXSfwTYFIOZiTgQmgQgc70843LXjKL+kcO6MO2avPRihl9109oXH5R
umPy/7RN/3QJ8M7UVcUk6VOHOpOk758fVQsuVU6yXbmROWXfvKlUxBNQZRKQjYj5
cMach7bA8gXV/wPFis6zegvAcBcRL1V5+wA2PTO2d6oiEqsmN2jEooypbimMgghw
JmKyPVJ61LpDz2Pmw8vDpciMRvvXFiesu0k4PwZ1H1RqqwNuAXFd9ysMtUGOK6cH
0hjZcEq2F2CdnH0XVazVtRbDoYG1dUlyXh/u0XyCBEjrjpcuif2bUktno8x8q0Ze
kFBWNtk/Pyn8eOIPxzvMnOy39q0bgI9bEIzy/E4h/lnk+aOXZLYBb0pnc7E6COId
G2od8DpQ14+wQjjRcrkqbk1RYjXTj6/rJaN5zUgYBFoui0UN/Tj5T6OFiwwhtXAI
9g2jHUdT50znwvfc8FasFq5pk0OWX+D1/gdL875QBDSeU0NowiqfkuCH8VbxI2gl
dJ+mHq304BEUZTVk5+xJPmDewQdjCrM+qEbabmpSSGsbX2T74ZCGW1/44qaF1aoO
lVPng38KNY9e/vcPeZ7U9RZLOIC8SFbAa90lbTQ5MWtMF7daDn0T1ePk6T4T54KB
mV9DfzPnux9JMSCOBrke0QglKMsQILkpCExVq9Y2gpdlGqzoBSck19exsLcDo7/m
Dt1qk/JNLuRwoAuUpeD/UlRQpf4Ojr2dByQp5vn2/B4hL4I5fxKtsIwUby174R02
vbn/ZTolNLJZz9f7PddQ3viZzv5MB5ggwEbv16OTxJYp9TiNdxNRYZ5Ev2B+rfaA
fA5uPRgP2iq43Ca41bEgHCjibXvM0AwCwoOuABq7ukmEHbEjArP9jQDvpNkODG98
+/Narhrd8I4gZ5mvJupAHOgGw3FH/TALGf+jgz0sKCMAm+j3y/NeCZ8E1YklyszH
GxcHCFO/1P8FLWQP5yMEDpd/LMaTfM+5Ceb72ILzKGhadKMpOSgsb1D1/sYBbWWT
OPcVhej8rTa3tBnGncBJNz+d0SMyrEzroET6Zacz+Hlvq2b78h71WF92pT6e6Oqo
Mx+s5RARrvOW+ztx/QCr0LvOM+9vKABgPJjR/7M5QnPUnkPXJsNiUWNobQTVBBz4
yKKlFn695ei8P9PHpXUzIB7LkG5xW11gUpyTl/VM/JNBC7XvzR5yut2InZAD7EwC
opsE31rRzxPOP0+sbPZQW6Q1JUE//vIH5tU4D6hReP/7dpCydqNcEd1ugGI4XstZ
/EplcFCAWJkayU7/S9VQ34//G/gqtyupFS7gd7y5dYlyxENlB4XuqoJiVSWsSHhY
2hlKde8/WTRn6+8UNRpPD5jgIU5yDZm9Xs1Mc3uleSpICPA2FrE/oSIRSW3LwPrO
WdyKbLt/XYvKmcmdiCM6o9rUX5gMgKAug6MXH0+d9c0k7fxk0qUfXgfjsX0gonmJ
DbZMV/EUJJhgSAtXzr+dtj4H6hiRcfMe25R2enURPtgfxQA1Wirv635JogoKdIBM
pX+W5keNez9Fqd1S38SKWPf7x6SNoxea3bwHZC4FQ4wphZgUE6Vwm7BLRulw6lGn
TPgYa6okcSfdhvvljI+XHa8NaF9051wtK9wKrWlgcma6KVwrK/Lq+zhjPegKs/Wj
8wqn0j3BECRiX3b9OnsgduszI2PogoeyKfAnR6USMzN6DWWTe5ABiodQzF5vQuE/
efB+LBx+ZBxrW/wTE6xASgpfZ7UmruVGqelbb5+t53TfxppQQ4CQepAJHQidWh3h
aPkO2l3qwhF3lagVjNtAp5+aMN3u8HABYqX9gSdlcVu29mHSoOVFqLQlt6wOgT03
AvWW3q+BwgVVEtF03gPfsOex9mxdpL/MP36k6tyaO6m8PL9BUIXSspY1on5Yrdup
Uxsn5hDWIkRYtt8792dOvNrfmW9kvcbiMOVtgBn8oP9KQLqSnyK6MQHjOjzfxcE/
dwyYf7LJrvSON6MefOiTS8a0ZmD0Dc+qgg/iDU8KmHUUkDyDawQK3f6yD6CceZUz
VJ5Qqg9y5PySTdkbbg7wg6PcvRMDt4G3qrTgEdbyDXkoQuE4WyTRp7bipaz1OxNy
wE/iRu75k6oo0yLwUBn8AQgLBimaAf++p2ovYkjafFDDD/aDcTXA0ELhhGRlX6RE
48RH3n3jRuzjmNtj3wWSNb8J7y5ib7wMF/VD/AcGuDlF66u/AcD0RNZT7BoEirSG
GPMvYwFgdegrirbvAuvhV6PejBH+N6MLblHpxPzSObEBXw1QawTM1KH9FSIBqQbH
lotV9PQc8VX1atFjjJqYZGUUyGIEgDUWExqxhl+cikgrDRS14LAaBJqXFL2sIIaa
00J7WCLna6a8AGkfjhqkbo9obL9v+Dge0V7f1E5mt4DMqbTw2F4Oi3IYsFxnsUTa
DDZd74mPd8dzdfVKsRDSS+CWnbPi7pycwfS0LEUsmJi71f2/pZL+s6IhLh69/1df
q/MCQD6MVkhKWfPtaOYd0HaZjtMZW7bB8ZVraC8LRNLAr19kLvfofYqCtN0JD04O
yvKRmClXiaVGAAiE1f5M1D6fzYYXEysp58e6N/PzGXWufm73Caqxjf/KbnlBEw4i
7Au4v0Rn1ss3x2nn92oRCBkZfNxwZNUNyjRvoV8KAWZ44WrRt9U1n3m5Bwh4dS8M
1Pa/LyTSrXO+HNmfpQYPR9MltWo0OuLoC+dNCFn0+F0slfbW3ZrEeDD2lHGXtCf0
j7iI9lQiZZIcNxKqXYQ41d9MpuJHYAtfoYJw0FUQJkkW+6OcrgRXaYFMBogSxmTA
VEMMyhPMedMprT9lKScTm8pBLDKza2LCmN27YeEUFn4iEBxmHY2lngS6J87r0Z9t
GelSHzE7GNLUnbb4EcbJ+0YH+VZ3xERIhKg3y083Xb83XQDt3YXvYSFSvHJdaYdW
jKVaSAw+aDNrIaNHw4cj8wb+xL7ygvdgjOrr89XQF1+7l61AFm9UE3kJb2xT0qbq
grYbq9dV0hv+dJnxeRDR9TyRQDEQerPjmEazJXmNfPNR7ydmAH3LAOcKk90vcSbu
`protect END_PROTECTED
