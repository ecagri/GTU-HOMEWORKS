`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QlcuiuhJjc1KZjW0sqhlxZDKAtOlE8ag9Pr+QK6a8NzrBuV/X5exlqA9IZqEAh8I
Ffo0yDGfWYum1upqF636TERVu78kJPl8ADMpmuLmvuIDB6/MwD6MlyPM3U2BIr3D
NU3N8JL5eWfr+p3jYU4TCWWs8fsHDFgFn1T8GUo6xcSrRZHRYRNU80uv9BR5u93k
Dxb3I6nsioatmcvwYoNvva+gF9ZOsuFMHBUQdYXTGkkBJbI1E0zVijWU9h0+4gTO
1F2KD3TFEWTjzQvKewP17ZE9zhbsSg3Q66cI5MfdyLqYMCtW5az7TRmjdOGSPghY
Dlka3ybB4an4n99gyuPmEP2JwyYoFxhF6bOZbRYci0oUjl9XBfb6Tb/kFC+SXWrb
CtFGTLdKoGkAQgJ8P5rw2MlYZJq+/gZDp3ZN8iaTuO/sINWT0lG7IZc2mIQMaB8w
umwSqxJxiioyhJQNUrYXVT3JfJx0EoPJ7LA8AkoVPDMkcbVnNa64yxMmwr79u4XU
sItchXYBDT8cYbPTr8tkKYWCgfq45x3jPVhFNddf3uxELt4l0R9LiJGSf3M6L5vn
xZx3WEXu6ES2r6MVYGJnlnkLJTmKTO9NvvBYEPRXb6soWLgMjXC0eO/tAEG86CyW
ZA//IMWSkM+KBcM/T/YPimMjpXNndHkjl5FjY+yIIdMFdl5gfGrNZ203g+cZskm2
8/LJJzMFTzPfay9I06eR+H9judD1vGbJI0e9y8Z+UZt1OoVMjt6W+IDQ1vHgvOAg
UtADbQyrgyCVORjxU9SNHmrT4RI1OE1BCOpe8Cey4e1uePXY1zXzD9TNGR1A/RsE
jizopuYsNBBbTf1sQy7Q3EnNf8svKwRfxPmxkwQav5eWtJDl6s+ghtHEufe18oMh
otHv261LicKnJFziHej9J5avh0PH1zl03Opjg8bPc7IdnbltHHuiexFBBysztNp5
lEH1w0TfgsowTRhXfKq6JlgU7MKsm8wdWgaku4sr2Hdsqvudb7+ZS2vk5Hywlls2
DmKWeATFmN7VLfZioi5Vd4n23Yt4ajgUVt8+y+lc2I7uGTJ6cZJK59+/C++lo/GK
FQ5QCFJm/8X72zINFT+N+XhFx/rClsZgqEeuOu0TaU3KYetSRQ65NDisFE3no+hL
QdhvwLeYAyJ220RdM5Puve2H9UHONV1abzReKP6703nPWNvjZza0DB08/trE0Aj5
0dNilXXpDNE+BSRBuz77uw/oACfALiuLnSiAhmGB4A/IdzJjRmHn8Oe4vy7pqaJC
SdJZuUJkhPMiIfJYNERYzGcdbqvIYZfivJWRdC7n54EbM33L7QDBZxnDKUhAyH4/
fTqiaeGQpZ0+63OqY+Hmvinu5md1xpJLdivpthfxDNgaeZQRMI+MwFWY+tP+ija+
B7SVPmq5PbG+hiTR0Sm6ZVrL6AgvYrhVn0zUpNLp6lv2pY2n5NbHOoOYVidM9VRS
uUCv3urxQpDe/GyJS4+cZ8wKPnYZP58gPNdc5UrIfK+ToegP3hKRx9Ucw6bUvOeq
dWXp6fk/R+TOioD3flqHAH1FW4e2kFb4ri8Wou4L31lolpzgeqfVsoqmszTME8lm
r3flQ3qfBc52zeg0Af4BhnvvJZRzpH1rqeiMOjIsl/PmJBzKRqGRfdj0E5UyuCj/
pRDsJMpzEeU6VhFOoFD56+HOm/NkUWao6piGfadxl5rk3ItKELctryv30aF7ZD3C
pnNaFkXVNhXVQ18KQ6PmNKJQvuktn7pirZgjG6xjuUjJJaey2sSX/1FIbUu0bKqf
XTQ/raT3M11lCX6yORKe/OtwfBA0nDe4vwjqzzr5pTzDzs7nRCK3Uo8AyFQV6puK
1/bHr2LSZyrtvlctkvex8JRMv6jlgGRFFVP3juDNreYkhtwrmo/FJsPklo3wBn5p
8IwOcSK1QaNE7JdWlc2NAIgO++dNUhQxBEi2MDL7Ok0EV7yvGuJTtGbq60WqJKtC
BxjhYIMUvdZxE+rjsXIPqslIS1vm/ZThbn5EtgFCtF77220/Ta9RbAdtm8dpArcH
`protect END_PROTECTED
