`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rJu5duIcQfB9K0OQwhk8oLmikcUbOcUpdVmJC67gfnIaiQkN6BNL7V0dqOMIxZgq
xZc+rbR8aNhhMYQwexoXD7oOhe15wP5PMNBfLhQKTiY3jeqJfuU+KF+8lu08P+pk
9dxvkQ3jjerqJcB7l2V3973Y9go170oxeOdh/hD4cAkXjLMA6aR1r42YdP4tl7pE
RvD8ytda0Zz2Wur05n2yoG/xx+K3/aYmB5DLC8RdSyZtJKPHhZz0EYWb5aYVx1uy
bEc5G13Q3TB9evGIuEUslVTwmlBhXrWpuofwR5FHb2tuLLOLbWqOylQ40c0fKgJu
Y3v658ArO822V5UOBn0m5qOYllJ+6/I6r691jwLXKXjzlmMhKxth0JQIBH06vwEO
3OfJ43AtKXXp8rieLFDyL1VLT3G2nI2bsZ22us3C8fC8Cj75ZtC++aLMrT00IqrW
+LPJpLF9La3G4Bs1Z9N1iNM2K6F2FWJ6+++C1L/4PnmLObcxfYNP83vi7UnelBDe
7Djsl1U4n72m0aVKm2nxseFqV3jJfKbKnjE+M0cjQxXV+6QcclZUVo9olkK+Kpgs
7Qt2OTZZkKq4VtdtBa6C8jFPHI8TdwMezPkv1FGOjaxyxdwuVFK69IWh/7rHZgfp
QNmU1ujgz/l1qGZQNGk5ZqmNqc2ntsp6Macg4Q6V09zyPthPNkzyzVutOH/jFIsL
VeyQdjzF6Sy1d/OjrFI7I7GCeSF59gzpOCoX5l/fEIvPdgNcnujbOw8f9eqYdmcI
3vkEYg25A/Vai9t6E5w3OaK9OsWouNm9XSTlCbI36HhOlBloCdjnANyuQreY/kHr
QgfzHOFgIRB8C0uSLWn0oXz3Zhdd9/FdxvH0WhltiK2o2lz7JoNzCDqE+MjFZVVt
lO5DF4iE/6ChVOX2XbHUjY7YDsiwlwuxCcDuRT54NwE5D4rUkGQ6Z22Ip5BiaeQO
u0nlQT9Tm++x4gcTGBimxgR4aJnZQFbJGV8ARFGlYJKTYi2fPiBRA0cu+wkvHSDz
bpbjKkxrxygjV4tC4vQv2OGapqO+mXedqRneiEYAr1s4oT+Sslb/7jPs2qtnbBqj
TSiJLQLxAbS5GPwTfhlss2+4JRQOZ5jmdX+iaF588dDgmZ9GU7iWMwH1yLa36wTl
9yBTth4Dz1GD2c5yGoy9EpYptIhkT2+Cz/k8GGK3wl1wmh41CVoNSn+6C7jPH2Gs
L4bJJNl7dRe3T1VqBzi1j1C7McqLqpZIeuylH3iXGk4I98Nrw3YzDvlp3FhwvSWQ
lspSEF17imphDoLoSmfVKQzi1iGyCkMjpR4S+5aCf9ZrWd1HW28NHBdvvzC8BjBY
qNZve2dn92i0z33W9EOQdYkVYoJOqajcu64Pw5WeO2pxp8Tbsx0wTns5yfXfzqFg
wM9jQnAke1mWkJlmwMgGcdvHhq3mk+mJ+y2VcRR+p+DADv+2OeudOhkx1+XQ7gbc
hX1ho57wBuDCoTFgy8zJcfo6KtX7Ece4OfGC4/vL5nKdYe56ZLZQoOtp9mIxyJ3c
hkD4QTNSXgAeQ0yVRirMF1GpBttcyLWCu9WqjwtsTwAP9TlLSCODDIVyTaP4sZC5
RfYd67/NFBo2+iSRRVuiBN7Vb9wEILnluHU7XJCy/r8cAk+XHtzPIdcsuNw5CcvW
ZUB2f8TQK9jL1d2LefKr4hccF9wDP532tZcVGwcmuaWpyj7LsePsY0J4U4UdXOUy
`protect END_PROTECTED
