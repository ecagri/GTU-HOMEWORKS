`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2TK73mmmsyQJrRp9Fzr1rfOKpaGon/R6HVYNbWS7XHufuxHUidoJZMEJdqmZZduN
fhPWHquZckUGnhfw9V30wBQIEhnOR34LvjcTir7i/tEb2nkvXfZ1/Xzd72VjhUwX
TraeRT1ddWJlyzBBiDb5KdeJRwrVa7akBBT+7wldaLCgyrMKnBpAKawjbaWO15Vq
vEfEXATch431VOwGLVbQo1UOdGk63P0x0//pA/LixZbtPkh4+6Pt1oKzFkbsrVwV
bS2zr4rgHOme/TPJhXS430gruREAKftVVGabDPh+QuwwlRhpCI/s00ts2ByvfhJm
zSw5X5vTOHhGrBPiFNzz8VRZmS4azIOiJcMFjDRknpo/DgqhmTSPtol90DTAOVE/
avP24cAvxclHIE/WiZ2X+MUtns4EQxTNP6/DMo30CAQqtYw/gdgbSU+7qZGFyGBy
t3joPNkhlOn6bL++aG/5NRPHwV7eqYY1EPIktMMcLObQneTEKDA+keROObcGbC1N
/wIiUhyafyYK111Z75PAmuO5lwIG3ml+voL0zPIH3Sa/ICDSyHhPFSfgqMszhT5w
7GaxGzcMC8XY9Toek6mQMzZSxNrtYWNbOJdEbZh+vwD5HlXHzsXUJkDdcow0kv14
rzQUq2EjqDjyG+okoVJ3lHYlG3GtWW+3lJ4VsMyRNGXY2X2GEmosS2v3miXYw0LZ
XW/uFKJh98JZWQHX7Afr/5nswg6QZevMJAW6J0SEOBEQ5clXZyuZP7QwErYDrz/g
RTzeryppP1p3DkDnEVKM+5bB6jXF+3OiobbbaA9IDWYTOmtgOoiU8L/PjTOx68s0
R2LuIfs9fr+4iS0hSMeTWCEWCQBO3pGM0huyz1v2e6nl06M9uy6K1g0C/hA0neaf
/ZTnSdEoutMdufxuN4hTsu19lkUL/ID54NlIsnymQvI=
`protect END_PROTECTED
