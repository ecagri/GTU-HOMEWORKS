`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U4jgByWsRS5RHzuvpoQGB0C1di8/UrMBXyDuvd6nhFtT7ClaTzvK/vI0UKjC/uOd
wHrfbGVHuQ4jWoVlyoY4ewi+t8RRILIr0JbsGPk345J6refVMKM0e0wTe1HBHSPD
Hq6RBSOJMi+/etgKbpfxGCHxCzAyslonBBlSrWdtzV62asGnaVJJQlYTmhaS0ltM
SG0R8jqpRhNbay1QTARyU52xpL3gh+Jo097qUONlbT9GajQNGk2ePBytL85WAiPU
vxLvCEXIfwuHWy92VibyfYYpgl8iqLFfKkIYwpyKNIO47bi4AQ8TYjmxq/uiVxUK
pv+hFOQK1u9e3uQwtoip6odokA++sbaBVu4rcVDnPTL0khLuAhZGuJp2qjoJi2Oe
PSUBLXVveo+ZRjr5a0IY7hd4eS72AZs0WFiJi1VsGGeXoWetTVV0s3vBnLgG5Wru
XRLVCb3cck3oHivkQxZbeYCnxfe3fqXQcUfrkDzB7QGefeDHDIginJLI0NqS3+WD
jV85txpDxLGhTl/cRZbzPg8n71qAPeIEOSdWGZenxfAFhMRg4nhpEza4GXjB30wi
khvNlQs18JsRZv2Z2/sKSlU81p1cbU9vsysQoIC0II/ILsjg7LJ03LjD8FYoS04F
9gO5cl+gJtE1lobDeejf8VhJZUBrE327CH09EsjZhcloGILEJpRiUDB5fUn8ngPH
x+jqjs93LoqztrD1mfrjUA3iWQZt582/9Hd4VmSc4r2HwW5sZ3B0lwJvB48Rj+cZ
UuR9XGLY5XGZJJ56FW8Ep0HqYD9sj2TnRKqR5vwOAxrw277LjDkfbw0O44Si6dms
gy7oK0uIfpZATttgWuR1IV1/XaFkqbwky/Hw7rnJUF3kEy8SS8Hw2SaRyH00RprL
N1m/o4SIj9YHA56zFq7CMVrccJVjBHViFNT9LRwZEpYSLsZM0mKMcV6yo7xZfd/5
m5I2Q+Gb0wCHXEpp+AdvmR1ggkbuZe+FcsRhD7PnqGXmeqjlIjCLKt/ok1RoPbDY
9c39OnSBhj0YX6yIh1D2YscO0hK/4uaBt+2jERe2z/gqCN+joePu/YyXl7pj1a7E
CaM8iyYznyZoYS3bioD9W195ENkB9qV3WBLHohVIVieyArrb5o1REyUhX4bp6W23
LANE2uKPxpv90KbX9k0RNaCRClPiv/r1wW0hOgOTWvbh4G1JMv/A3x22KeeyLoj2
ez/N7VRMNzL3PiIvXxRVrpkoUge6/xgRVOBz6lQHIBk=
`protect END_PROTECTED
