`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hsxbEWttc0J5SaA3jccoTRlMk2dLC3pNmpftxXSb0ymOGfjL9H2Zw/2vyJNoITJc
YSLeXfStBBNaBw1p1ZTsKCapC6V2qA4Bg1CS7+zhPpWxU8a6WmERMlM3EiGgAbzR
ilGrwI3Vbos3qTSVH+/TKN9ZDuMxkF3U6242ra6GAnnCXnxCd2MQq4TspzsmD3Zr
JoJB/LNZJ48Llwo2EE45ZR4tP+nNubhU/fsTpg/vmiJ+gSPlZifCYX+yE9DGbEJr
U2hIpKYmkLD0huQxBIQ+3HkXa9klGkTET91z4nsMUEnfSy7ADsWDjiyXP4agKHmY
S8vXad86/kHrdF1eZp4hEM62EDfTAp/FhL8LLrDW72WxZhlKNvRfSmW42knucXc5
ShA21ac7BGG2X7uzT1R38AqdWqu/pElsMQqVu5ZbbO9OqvYalZ8NbRUjSaflrYSk
biad2Me3Qs4G4W0/e+ya0YHAqtEEW19AONE+ip5U+TD5WdqREf8D6fICTL072Ib+
MX9RPv3fXQl73uN8e5vN5raVShlLUML8HIqV3mBFjgpHu5n2uYqor35DRmt3CUsu
K6verSbmug8MwGu7hIgmxYqEPYaaXXKo27hoIc566fHfXPc36+PZsKjSnmYiav+o
q1LdPIxwbRus/gB+qEjX1kuTbg9a/q2VKAsRfnp1Mi/aymBl6lVQKyYWtMtINjwQ
+4WEjSArWrDnEQ51bxUywE/M+79vAXFa61TjqodDA4molxjDHvLJQWjMMtP8SjQe
fYAUOPwTr50IP0xfEKjDonU9Lunj8jbsOk2S4lwNiHz4gZ8mqCNg7/yvXrONDGqU
KGFCURiDGy2DIG/DTHY6Mwz/FSq7IZ43HS980zfQkx4Cf58CUF5bUpFvSc17fq6P
tKI4PizM+U7cKkTiCovnf2v02146YWt/mLYZPtX5U+DvC1ZmJzW/61GYDwoPyAFv
FtgCAAD3dOU/Y4hlIp1aybf7LrN7W9WoyXEWrx5KEEoF0N241K2Vb/4UcSMaLIFr
e1B5qpHYbi50vL+PGcmJxZOpd7+FelS88UPgMEsn1NT1FrYcGw9s5iNrUBF899ab
sn475M/xSp9rVaUJLQVKm0OKDxe4q8pLeCJTQXGbyspoWfIdmFHwuE5Z9SAoI21e
FBgBZcQsdMgUuUdNOQyhrdbsAPabQ8n91Xj/KfTYMTkce5nhEe50BgSA0hNvcHDP
KNxH6OdCS8xkKFfFWCMXj0lsn5IdaLukWqhtOcPMhdiZ3Z3P7uAVOSiIQe3DxWiW
WSoJnMyRMrkUBTIQKjMppSirZpIULioQQdnWkAz/pGX9cIfYIUY8ITrUTeYcQ0XS
rtfTBEaBUMyx4TMTE+mQMjw99EJ9A+1r5guh71n9Eeppkzh+tdpmGrHSojJ9x9QB
CFVjRWkpqMGntDUB0g6qXITCyItSrSZiIJxcUQ/Cew8n5J3OpjH+RrYLJvvca0/a
BxYM+0IxiOdb9LoYTgcS9yEY8Q0m4fY0P1jVT0tE1AgWur92KjZeYOoE109WmaX0
2kz3knNYDA7xx9E6Vhg86vCyDEqifebWiIbCqh0nDrkM/jVpKWLx0PTsUvzcK7Nf
A0GbnZSONhpj4bG5D1RnUXIMpi+ErHRAiiqeF1Z3Qdc8zh74P/YqotnIClDmq6Yw
ki4zfsWgaEvy2dkYa64aBwRNe07/QTfDrW65Z6tyftRkcHuzTlrjITpZ7fuAKjK/
ZbjLcU0JotoGQ3i4OQ4jkclfYo22uDdNpdSHHrp6ATJtAzUJ/3fWGAE6dxQiitWS
yA6T4MwezTihTaChT2e/d327ZuKpngyF1PedZDAPwbbEPKVTu1l0DGQVrwsVvz9q
Jq2whM9zW+ZkyhG4CrqsrE8DAOyNkUlbow+uncfc8J/EX8sVnBZQKZRNRpwtZ04B
yRf9dAb5ECFi0c+Zqv7qCqNOMB1fOv4UZ1aQpEyAs8QotRJUFboi7Tp2Yqfu7/kl
K+6jNLcpAAxval++jMw5QcReaBAF5YivjW1C2tp60DE369poUTVE3KlSyIjvfqx9
Ir5Hv2Uj3hHSWHGXA9dJhdHZPOImHFq2MdvB1DeW2mKkoGPMVduYHKIZWALt4t/6
/4XG8doyMeLOo0EsXPmN/Aztmbf7bbvPx7h4XlJjfihlQ7NhtOlxcCJaO2tFII31
EVuhyyOdxb13r8vwvMFYQaF2A8QY+QIUi89TUg5t1kNPY4xtw6jKtPrPQl4T10MB
Y0SrBDFAJo4diW2N+p3NdsLqNzySFpX7dLlL8R1riULB8t9DFnqJBxxfE8U3dUHM
k3kCyb5j/YuAvg131tB4WxDSfhc/NftXqhbFrrZkr+iRe4mAQFG78vDdcopT+071
W9b41JPDwvDMW2RrwupuBq3t3YoUmARr8gyN5JKJF5JNETA7bSzPGeg7T1/8NOoz
a76togKt3L3tLKs7PpPAR6XtIPkjGs575FrsMpS2QHAdFAhHxNXnEiExkHeBi/GV
JpNsXwoldP2f4klLZF1N4jwD7RB0ljzdxGSDsFWKFd4C317lMY/Irwp5ZbbWx1rU
MUje0CL+1ERTojYl3pn3nwAuovyiiMNQ3DnjkremYyqh1zNAt4Im6xdTqO3IQ29i
dz/OyrO57opfOkFuCZBUWe4QvEdJ2QGqbcDAjeLCcpc6lPe7hkad95hrhiouQwJO
+P6not3T3Id2o0CzWs8bfpKNVsbjPxdq/lFSH71Nq9tk6GeBQZUvmiCCSZYrGOfF
B5crQiqOk4KRb5OGb+vYT8+AYU6Q8dCWyrk1WcSghwKXGZRgQCOKmI6rR/kvm1DZ
xvBv9xnlN3iY0t1asXR770vcKbhpeIqmtbTUrImYiDva49cB/duyA8o8XYY2CW0p
2NWHcZC1YV8VxWwxUJx/FGIaVk16rwtql8wu+yeNuMXXwjAaoOT1r6K6cBtN70Yc
kR12d5dQ6tYCS7zrpGjuvSOv62i+wYZ/femBUPbBavEoEZ2yzARPN3Yup53Tr1H/
s9scM1fKkXmONk3DFltTg4WG9v7ZsCHc5UN9MT3owAjOdmZ1/kR4XfQkAJA0/sLv
OWIr2VIPn0ap/JCYQqyUo6RcwV0sZ/6GwwZ44ScRi4U1DttHXecn8Cu4OsCNVEIm
gF3bOxjLc5t+4JSqNNLitlogece3HYsQJCmx6iQpatwYZX2VVropB0QX0LQwuaeL
HgvAvueDqh0NHa80zPqrZqZLGxWd4GAPMLebQMymzYPilIMVX0SK6iiXJS4OyAgE
3Ttk1BD2lXis7F0tlY4HBLmMgpo4hVotYNltDH6XLHW7WW5MHopxqJ+SUxdy4a86
xThy0sxEhL7aoJ6Kym4OnZ91lboh9Cw2o32uh2v3FH9r0dnBPO260Yq7dG4XeTxi
niIO+jyEEtMe9pDxgkiDBTXghYmXtq/+VZ1MBj+s7OKdoaPeRuNTt08+wHI9p/SV
WtDxsKE3kIObCT6HwALjUU/PITRensrlYH4qjXGpFcKUA2FCIrFIWJJkIPLxtwkT
DSB9tfEdfdYSRZl48tO0O2xZA1WTMh6TdQdDtsPyCrG6pVAKJxrjrjWTD5bafA3z
j7EtjYdmujDhFGHmF3gUiYYWulqm8fQ/BRwEXuVAupQh/eywExKcj/3ByMwHxgOi
ZXv3NumxZMISmFSFN61LJt/MLynGJxeApkQJHhQeNnwQDcOPOiOb47mxx6+Ai3U6
qjyN+tuxPGJge1k3ldGHW8nq0fTgpfDZL4Rb+CFrEhcGaGQdl1c/BgJu3ZHRBo9j
p5Hmnn5A4s/N4YbXHLkPS1wZFVIlpTvBk4QkEW1liToKsyIszYulrJvN+2aIMC9s
Uz/wHecSMNkx7ze0Tl/ohhIZ4FB/nquhfR476TIp1i1VKYtU5CMVOMW28Pxf/eVk
6qHpTuUf0h3tCTlZFOlNPrHRCufHBLzbJHiiiJxmomMv/ZK1fDzLYYGxk3sSfDh6
bti4hLQzEe1xmvFjSEPfuZLbCHDHkDiUTpCQ0+zth1HU6OUWLjgGW2un3KRIZg9t
Vs7sPeIH+xiq+ZKlfQy8SyVEa547QSD1T3LXgjq1bYdRLyGAJVAXXYzPGoHajkYH
TctNvAkoTPSTUXTVtKCRvkAiCyd1QLLxSEN+zXbLsF0RG49VmyoTHgHjMTKbGE+F
leYIhZNWolzAF8Q53ZoUqNkD8ABIWAXPxDXJ3d7jS+KcY4dOtovDCYTjz5cCUaGI
tzSPAEPogBXGPxIDVbHE1xtYKCyAsch2HLOSd8pus1uOB98UFKpHznW06U/hY6Ll
+ofQ61L5+FTDpEeSsFCZ+w4BHtEIBmeMgdIEiIxn8IWoVE8YB/8vsdeTei4soqas
wGT0tgbvHugugteRfFgaNSFQ/GoVWqDW0FQx+79t/fOTbilaJIpN/V2sD3YFFpPd
PiENGr1XQvy/UHKNrpzJNZ5p7cXLj2LLZuXv1REcopD099Bl0dtCTLFiplDD26+y
SkqHPoOODaY9jPmIK/RZnU8PhqXZ/K6+AzPvc+5cKIPP4PD7ZXEYg5jCF/4Kp+PQ
n/K3XCSZx5rubJjl4rMh78DIvKHEa4KbQUUkKI3Ir4lJgT4oxDUfLXYIBEQesh7O
j6qJmqr8vOVEpekqwqB4rZQSzPIxO2a3mBShzDDOLsm+45PTQD3O9d2vugkJCBbw
WiwHmQ2DuIvkAZkhf4Iv4K6sHJdaNpnDw7laMwmw4LA0Lc0Htkt4H2Ly9jNFtQ5w
qysxytjB8uQrS+j1/pPEJaBIzi3UzI1PcFk+PqoIsdTsqu4NOOyevv+g3kj+euNX
6Ik8N6Xo9++4AsGr123FdDccTw4A181GDWvEOFnJ/Vh9TldCJuNa24nP3v7ZBGgr
sEu2MNoaEJ+rT9zNZrFe+M5D0VaX2ZHaEV1bwiY2UvUveLX3czQ7xnEKBw1MPBhk
r9ppmhU6l3ay6Ze0Zn/N9F6vDeR8NPnaesY47mN23nhXg4U8E9AG8JF3BHWOb3Or
znRw+TJQwwwrQ0sWlYRFX86lU3WY4I1jdxwOIhYeXtzrrfDpcazj6STDhzHBw1dg
uwk/mN2j6PeQ8b7tVQOkSErH4kgDJI6SPdQg3ezng4ZjMFkt6660AlshHHjeHr6o
Tn745UGvPtcjyQJy01/02wzE/XjBDnhgVo57jnPc7q4AQs135sD/eyR36aYZCArG
Svk21IYSd9FED28yZZG8JXUNaQJoguYD9XF91yiPXPxBM6gfr52vYBBTP93+PSi0
YJgUEaOypouqsXS8CAwE+ViakZZ0IhEWZBOd+uWS4yN5H6blIxgARw/cx+g2FJul
wrlwKmQX8/kKKXpvBMMFnX+adj1t7aVNR5vWc8dLx1F4qhU5qBZBYCTrX6IbNuYr
K9WIpK7gRF5ku4tCAPCc8iCPHHj1W3qdWnOJU1uL4bSeth7F5DJBD+/wvjDX51AW
N/HG3FqQvw00VX7nkYkV77uRqpylQthbK9oBhBm7E8zlD6ly20eqkyi3t0TLNkX5
ooZWEV6/Pb6mM5ng9kHCAcimFE6EFNfGfA7g4fYA3nCjnD6doG4jlCzlevL8Cv+U
3gKr7kXjiXJl26B9py8Y99iw+tAtLBOaiTJqgrSy7Fqg6sz99hhuBBLAEjsV4E4I
t+gMy9l+wDEsjFL/NmN8gRIAqtwv8MVRdo7DF2gJJ4O5205qnl/KmPIYvuB9WaMG
1in9kWsRwNBKBT37L+YZu0I6lOYkJgJvugIcjDfVAZbeBHRdCSBJXmv+DnTygGbH
SqoWhi4xzQcno74hXtz3e7fnRkPKhto26M0xcXjh2RkDj3v6uuUuuu1LtD0YPWxa
NCKRxaDsScGgXdDunUXwUmFfwCSjedLuZ3AMPPV9LbQ/V5WNzJU0bA1WhnKbQtGG
lBbppFN0fPwYQNJYZjLzjvGfqn4w14HpXvZlzI2WBAot3Ywt0qX6Qb2HVnv/b6ik
cOgWYvdbypjK2Cha+BEz8VJj3sZ1nMPSYV5j4UPhTKZoKHRdnJLHAXqDjOeDa9Ow
`protect END_PROTECTED
