`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tuqqn7D0BARGfa7sUzgXdaWuPChA4w4uloF+KzqfKod6TzlkFTwwmXmRLZNm7J1b
DcmkT9YkajpcrEd7Jr45yAJddmcNnyCOM+kmWJnd/csREwuBODy2lOSVDLGmwLxA
T+oLGW8JHXSu34MMokDymthhp/D6ZP6CkGoEcBDQkkHYD2oNCN+rMDCGqwSzwm/3
xemQgl75RKaVQ6Whs4IzGYZhdUnZEpioYA/rEQvlOOd+IUlDp7zfPiP4KkH1uueo
qgqIpQWcCtd3vCoKUoKceMHOJRNMjX9V+y8IAvc9nq0Fy63krOo7FAZggAzd9lJT
a75tq9ZOVJSXzudDlimW5D6Wlxqm/w/1zgvYVLvPHx+cr7z89juVBOfIt/qoLWee
gNt081+suy59yVPfVk6OVQ==
`protect END_PROTECTED
