`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nq5+dBWTG9Lej9x78UcxzPIm2fBaE5Ug8HrCM0iibSS33XAo8EG4PJE1HhIGtKNq
dWX+c7K4JltKFL4qzmyMwhX/WoIni60UaduDW6q2Wmu6fxnEzITb7c787nkyp38V
O2+pvt8Hh5JOVl35Me8JbJPtShP+SPx3kiLzMCPTuKldR4wF9qSyjfQ+LB199QLm
RNO6SbBFzVWDc75drl5vES0LWCMI+XH1TUbTFS8QmQ3uOhD+FDB7qlAVUQgEA5Kp
07YElR9pTbBnuNahPDEeAT0eRUAEaJcNgDvLMc21uHQGXOefWvXjJbkjTVNTFFzT
jeIzGgFKnHn6qjABBk593C9OimcfC/WjLEgZriPwfjs7SKAc4OQNK5wHOUq3jcYP
na7VUCmMjM7p+B1bU45diMo15F4vjuY99A8HUJZnmNYRaeF5Pqbn0mx130dc9GNg
G2tPDFBsD6VAVWqEeOKoGWwD7lblXa48vpZwitpZuOyuZuebCEyMD3FClVjEoYZv
vvaejDPaVm5U6K7mPUjox+XDEcZnCqhPH0bGbyn5QLvzQLn88QS4kYKpRZAs7Sb7
b4sFdUgLcxpV0XBwz8Fg7K1AZ92HZWcCpKTpsP0UquCLg1b1ezD4YYgQt7NacUp4
tcJ07SYx8Q2NeMWrTjwmSpLVt4VYpn/wGoOnt2ApA5JenZCvWbbjXi9V7nEqhqAN
1EogHinhQD0xVN25mABjdZ5QmB7UbM+pDk6Cn6P3imbpjWq6DDO/cFKqR/nmTKFZ
cimQSOlR1jN9XEp+Uk+IXdH3cMp8QFhJWzAgRnJ9pj1cQbjjc78K8CSX7utBSe/s
GD9/WCIsNdw4pvU9j1MnY75cKv/3lXK3hBj2uWtk1NMVn7NOBoPaUyCMpK+U2h9U
w3xj2YX+aI4gELcuKGEw0u7qrtbljvP2N7k8CnB33Ig15AN3cJHia7sTw9lrRKwY
onrpPXQPGLl7BLfMuvenDtDCst/Byr7UR+FIAfqung/PudX/MYRrC4EiaAnfZ5gS
jtCGWA6hh9ADblqxS1rr8lf8tGIY3kVRm3TFkaMgOWEKwvAk1L6C2QNmlLkT3jBl
yJQ7cqOBMJpqP6T0Bhyf7TwSUju74jI3F4c4ORFtFm2xm+M3esmSexJ0oZyMtHN9
z521wWEg7D2OJRUkEyaPBYt+0dQw+m0K33Is13fVOeN749ae+slHGvwayrwKF71r
gz+kFrjb+0zaKU8HMeazA8KJOuEESS5cH1UeG+SkZHRA3rwlZi++gM4r64dW1up7
h+6/b/RahPO3n9KYmiXw0nJzL2Aq7MjihNTbmmFFWThmkUcoBjc0R0Su23uUktWp
gbf/SqHnvwAr6lvIz4Gn6IBmBI7AubyEk9UCGRBPsUrKME13re3bwSpHg2XeY8o8
1pR1TQk4XaFZsdMtWafDzQghKvMfGLkTIulK3rCwpoln90E4OygTu8U/8KhuUVku
k0/PD0M1OR5U2UzE8pQzQJypxAUzzrstzGGYWkYvhLG/EnOfqpTD/Y6Esq+/YAmd
rc/WGVVJdAx0SbhEaQ/j5NNfGNvooLgAKCM7Lk0LVJjV0RTiPMqCb9jGxzAuz4Sb
x6kPop8bWCXzLwjBWTzfiV2S+9hAIubZtB4ZvYormPDKIP9mGNCiHdsRoS3ZJeDb
ZHqqVQdDrbYzoZqnprL2zwiB7iUvH19QwEtTUKyogobwFA1NnoEk24kWSJqVc6Z+
V4kPVpLeEusKm5fMs4JomATny9jVhYeTzjPo5rBUcDkWnaB6ubtrbuUuFUnqDRP4
8wLwcGK1rjkmsI+AjwVcXq7wQCRPp27Wvy6/ranQOi9WRjGDYbaJgMLHz51xXHad
4dMG60NPOdRo7TWdao6gOhmWaHwSNu09PTNwLKOwb0tGGwtYBubvzAFAT59Ff5Yi
1DMHCe+oFEvISRq45xY8iIPZ14OxD2erz5nD0iG0TbJOuzSt2ciiW+yEyuhVqQy9
5+hHS54i9kW9dqeqC69RWBw5DprN6vPCp5xj3eVsmM+hOb1oY/11qOdmXI28M37T
68JvligwB1NfjLatvUATm9N/p4pk2BqNVwS8waeBMcUZRN6NofyC4JkbEaRo9nxo
Rwd1miIOwJJWJgG7nqexJag4U+HQOgLuEOzRSXXW2kcWCpB/9VsPx8aAt3tzdJGU
AxRLZk2iOSLzxU+/2GvvcijqiEjSiY9ORX46fz9WcnOKET6jLd27U7LCTZ+d2Gl5
zb/o+DWl2TJ7fvdCx/r7ig0Cc5OkS3YgzpwsVfsQdfk+1CN3VZo1agej2wktFi3W
ykJ/BJgAuiPg0u3i+Sc9QTOLK7ZVl1XMw1HZRi6U5V6+giNxCFr6B0xUDda67T2S
f4M5YR/RUAWKI3GesweqvU6nvYqvcapz0T8rz5DpDH9PV82i4SaT/RXwyxfGiYdF
5MsZkG7ZkDE/huwb5pqWrSjdpxPm/ZsCkzhVpifNi8e4SN8RNd5AbsqgrAtI5sFC
mSZlFR9GDXuIjPihxjdUuiRRWfLfD4zdgXJbLykxYEwVu98UAZrGnDMvvs5zh8Gc
bj1NRIVa9ZAlfb1Iz7gxOAS9Txjl/a/1dI7coPqEMxkB5CR8OIpZja1dGvRfRxtP
kHHakiN8bGUTRX191nZ5NWSnmu3gV5awxGqHmaG4SNoUl7KJ72HbOvg/J85wbiKa
nbx7RjjHanHrOHEGKwYAPHksxUlSyn1gwCIE7r0/i3cmgi6cyqhGJzvGYsgOdRN8
5UinxFPezhWHNUyPWm8Ig23Lc+2GHQrILlc83RgazlIG0LD1plEf74mOTKo7Ta/8
piPcqrlXeQ9R737u4BMwu24T+7tLMx+O+vHk2uQBbuZxTtEF66rPxHSmlRbvz4DR
vyHZhJ/8mZz7W5TFcPaGLGcAdkYJ4dtmuzqbO5/wGt3TzjfsziXXREElldUU7aMI
NXuL2JIN53RFehzTGnur04LIh3XgF7m3wpWciuiB2uQUfriVnKNm/oQznJS+nwws
sgnn8nHCcX6YWSXtr7dPojb/8o8Fwv4dpiPhI8braj7eLmAfz9L1tsAC3z/oROyv
dwaz/PwAEcwKJbVT6USvRkTyUSfWBOWMnvTH4mGcuN12t6ghhSaIlG2xJWIwFGN+
Ex/EYGZ8BdMbRkzFIo396KGjGr1k/B7lbukyhyscjxKgJ6PqrNrjzarSWGE5z2KB
dGJMpMXvv9DBhAXhwFZV/phLrj9Zs2A1muLA5C0mgoU5AIdsPUGqDJLgZ4tnZkPM
ZtPI7wffHHL5IsIPUs4/mbbbumAfSKE2Upg1gD++EEw0pN0TlkTO5gXJKEKemR+H
SMkMlBNy1VTdUUWZMUUcGxpHDEgmDnkn21VyqfrGMMSknY+Yhtw+j7CXEG1fsw12
cdqItWablXQwl0Lv+5YYGhMseMuuF6poPn016MAC0i4scNgKlgsutfPxtuF+EFRz
e00M5vV0aQfsT9gbWTXMhEnzdJ9QbunqB3/crHP8DnrMsRwC8Q9OMU+lvWtUxDeu
3j1SvwMmuZXWi7rwd+uDZS7kdAArnBRLvdeCPA+juxgpFIPbCJ8vZUyELtY7larL
81aZ+a+MjB6li2oHaSpiZJNJLedt1VnbOIq8RGwlQeg14j6dok/cAJzOS/4TWELB
kUW7BvqF8RQKhNGvTTIC50bibG+Dt80Fk0w6PKwcJLpReI45k4BnlLzYP+4IZPzN
F4esE8jPJppqYHQg9dOWI/QtrdvHtdYDHKJbFnocA4vQoXM5l0gQXEWKP+AneUof
H/opGStkfQ/GIr8+ioUMekACisw1d4Rx2kkvYtgrVPKcHllfFuqRn7joBkxhDvyN
YTAZzmTDb/f27tcFn6M3MnxJr2l363TcbXDbG+7myJ8hZ3oaj0aaQKBVMuRSRiKB
gzDAnueedIqpYehqm/L8I6ff1GbnHOMAXo00VlUPOQB0JigPRtRkByB/PZgezq9M
Rix1JBYgD5/hRUDCdAJSO0F/q7pCdCwvvp1bmcv1r7MFwwfZDP6fIHn8IEIxfoxz
N9iApo6gIEOICz70r9efXWebiQVMwSkrvYLZms96h0mGjI79ZibL3QK7dz4GSnp8
zyFLhQ0eORBPpQoM3PfE9UpC0XVtV2NdlSXXFpH+BPsfyPxitL3J6co9Je3nwv48
`protect END_PROTECTED
