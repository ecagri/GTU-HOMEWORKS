`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OvS8MG13zQXZqSv2x+Suq03bd+SIzeu/2FE6gfcDGWvBwPb1lfTo+nfU23bCCaK0
m9BKNo07GjSvVDUpOh10Nj/bHLQz6i7Zuu0VlpdWdBJW7zeAKku+ee+gwMeT4ZW1
F4DnE2/P1TQO0j/yH3w/nEQjvhCvvDISWav+7GQ0J/0w7iOVqyTUNkTS5kgsddUA
2v7UKOxMpshSywE0bJPXWgxpJNi6QPfTHVsh3Jvrijjoy/yETmUspLeEHcjBKd1g
VIDOu+X1ILOhchPH7SlKmuAUq7s9l/Pnts9FETrF1pwHOz0cTXcQ+Nch1HKnq91K
WdZWAy2WSGcU7oQFvtbz1BTjuYCeuL86kPsShgIcG6JTVo5AkIALLMo0pDbHaLAS
WKrb1QmeZJYhL3KZQe7r1o5f2RpaKZuW3zGNgfv5JqW8rn5JFxFeXwWgQK0CzmgD
g/+7bqrfx+tcfsPQlBVpLiJ20T0Ls/Yua+h9eCmQSmKC5n8z4McpYahkDzJE0cD9
Hg/2wUeGSQkrbw+b3SCOiE3Q6PonXgLp2Xjg8UMzNLr3r4GBdNXRGKVcVB6uHFkD
sr88gLhZlpc8Z9DVJUZHMdBodbF2JAkcQ0k1WY0K5c6rzn2riEfzwMYTDhj0CDVF
pnuFxLH19mIL0SvzibZhjxFp4CVS2oGvDrEi4227Mf33oWsJJrOsVkKi9vwbhFUd
NUjAtdOaLvc2n2aUveZmpBZtQ9BiIj9bnRbg1sYfoQKy5a7XdUxFqFu9YDJF2xsC
4Jz+IbvLmO4n2di2uolVrhhuB7ij/yG5LvBsCX66dXtqLbXwD1OkpevV7j4YOtM5
diZSbXIBSq+vYM6IgU5BhuyAD1nLJXy1WHD5sJ9WKvlN33KJF6mYT423V5cCiu0A
nU/UFG2Sr/ioKIGO165gxDHkw5+Dt+hJ/fcCxfwZf3ZK1yO+pIeQ90dOR9QOUmjJ
qkUG/Hnn6132JNlr02pwZeZ8sLKhfEIQXZ1dN+Bbt1MatqfSKM1mgou9Z2Cm8ATB
gOZwuV1WoftMGCCTefov00vouyXy4zSifZNEwoQOBew+4wt+prRBhYqlSx0JTkKi
pAqNWLVi1mQYepgSaGl9a0w4uMu9DQmeASwqC6OeVc2h4uGnfUS8AYm5j0bYQtvR
/9jhZL7DPItF5f28Yk9GIvuwim7hBDHjnP5ttRaNIFDqD2g+qq/tr5mb+DW5cxUw
17/IIsgfiNm6WkPgDpwGfUOdP2C1he10yy3SF/+b4SzEKyCraKZr7zesl3WYA5iI
t1oANRonmaDOxzEJ+vYs1k6hVLTW+xbohUp21wGnlDXLspEWrL9ACkFic5N5lOpX
xBqodqY8VkGECNOBHi50Tgb/t+vRrbIr0PdMsSIS+9ezzsaHr+WyI5cQTQ/4mRdy
ouT5GbiXO10KKqp5MINizXo7Rp442u2c76/GBAHBNlQqiKO6pHbc6gr4/yIHR/Is
Y5g9gvTmSqWEdH45xPJFbsL6f2spZDva84Q1N7Wi56LxEeP7N2RLo90dcv1h8Fng
UmdeNwsdFy/aopy9DFi0hsTu2p3rqk+9/sapxEY8S3l9yTv5En5LiBMybklmNuRE
I0wzCnwXH+8STZX6CscFGBB1oS6RSVKXAUpDZmIM2gcPtiSP3/YcvlTBZoKJHdC2
Hd0/DvAnzUfH21tw8NADezo6shEAPWETepCPWWUPYPIABVMXbLhozsSSbIQm0JvX
fCGIVEVHrpuLjWzPipy0nppsNxxKpoydNRUMw0Acnrd6pnPM5W4xsZCdbsKvcUM+
N6/eG/mlUfRGDkExmEfwSo447theietJZKKnczxIa8/XRjHF2w7g5Ae7B6ms8ogJ
U9SJq2EsYqJwTxG1RL9/EwXw0BNxaLQt9O4I/ENZgd0q2k74ZGmPYO2upXgPegsc
k0571OIIseKmOKL78jE/RsiXZPvF5QJfq6POYhGfic8wCmwENQV3di7xYCyYRkEZ
a/tRKfb/HyjDYiRHGcIv8M+fj7FdDl/9yWp+IgyoWTdXA1Av0IH1s/uM/FiVMp1w
CwzxmVPP44sismGOWRW5NQKn6fZ+vuKEOCrZ3RqVrfqndu4oMYcLs2cX6Vy73Kr2
xDK2Y+yGdrxkxhKkv6ysXLO3oVfrrAE5SG1TKnCNKkqFCHexoruYNie0T8n6UE51
/oiwGzSe7Yrl4UtsC8I5zEjyU5+vv/46wX0c9mxcL/ek23EW+TOiss7r3/dok9w1
r4VUkRSVDV1JkBPPZSTHc/TpJClpJZlX83RK+EzxCaj292m8ptNp2/AXN7On1sf6
bsD6r1yTGzo8Lu9Xir0vNu6DUk3XKBWbWJth3BG7w6tC5inb+7kWcpcp1OaigIPR
VXJDkAkS+0lX6so4mGk/1pzc82d3GDYhjmIpfBY1/CQeeeOOmeTuUTrp0XRW197W
o0tbwyOwoFs8f6zhiHBQlwl4bTxVTk1PFRO2LeLJ+DFB3gkfHUBXmC+WmwqyW5fo
Kpjc3N7oOjlwsTYJQ7w8ORh864ZO4eMEaN8p4/BmSmU5R4ITl+GYs5LsMbXwHxhF
HWxkWj1I5S9s4Nz4TojPlRrFWApieE1tMeaHLFS0110FicmsKtB5ew7WJjfY5J+Z
Pu3fYagmnH3bOqVeDmhoLnN+Qsaik3HrXA5oVzPRwkpwaLg7QSdxnOdv+03JFNxK
5PSAzb9Y5Q45KAeDRMMBxpli+zh3DG3+nmT+77GbEXbDR6crDE8bbsaQacnYUo7f
0az/aNJIoQKK3VuG9TNc9HbQtWLBDWM7SUZPA106+Sz6Zt/2frUE9Wn9bnXjX68A
w1MteVetJVZDBX42AaoydvcHUgoMX9obHxSf48y4JOz26LperGUvgkjVRDiJ1R/q
Uq8Y1u8TJlxUGuTO2NYcUXzyX25NmERf+5bI1THsjXQn4MyI3Nn1y3klHgMchL4C
a3AG7tpKf5iFh6rdvHt3mwFxn2U6FDgpQxgjBWYypVtjXONQl2go1vovpLInhPgw
rQSmppu79BvFI+r6/lPOyr4IKiFj5tUtvnnZfw8t4voLesrgnxme0wZB5+zGNcLg
PjScMcfAE6Vy+9a9BGpWdqcs4/G5S9mV/JjtcrkfU2z2u7tfHlDod+n/7Sq5liep
7Bese/fFs2noH2Zva9B/SSyPoXkD3gwLXQ4HhJdbEVy5czWbwDyBpGf/V6SVkXFC
qR+RBKx2VgUbDJG4DhXxuz1hL1PqiG08UOmfXj1jv9C+Mqz2jfTZgTWjsE55UCr0
dFkJSLCQM7U5J8SY4ypYOjLjwN72Nmh1RBI6FrbV4AukN+VtVJgWZXJuP2uerosD
y4gKCvlNzYCg8/YGm84QMBBfsOCcd8SNZnzFKSzSoaZGmKLfNr5ha/ESiZ5MvcJx
fnC/ZRJlbLTBpM1kEOKKnKwvMdfif7FSur3vYjiTy/ubqiwG/VlQ0UKZg2L7q3PL
3TDYjnPCDwSDSBh0mkHjywW7x50UYPCLKUTtlcd+qfNc7V72SdLBMMN2wU/iU0kx
26s34Kvb/i7iZ38LWHX9vpyBctJr0QgC2GK6LJ8sw4mQVbFIfTwXtHWlATr1ye73
uaVqPXm7x/FFqs2n3goZBecmnGDL3zYpZURhMuoGZeZLV1woAAj8jpuFxlgz0DOp
Rm7HUkYgu76hyjfzjEtpGkgdHkfKGttjA0wp3GbgurLDHhsAEPURozWUG9ZMjJov
`protect END_PROTECTED
