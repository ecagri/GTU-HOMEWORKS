`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HJ1lYIsLqpcwqvhSIuMBWoXF6r/muivOhKE4INwkH3dFch/6c09ZJEnmsczWX55V
HRLqA3brGLwoKfVL7HGBhDw6q3n7bejTWFu9YIumykHozCpk8hBn7FX02kx76f6/
rbTiQ0Q+uP9KsXE6JBRm1CMtBlwVZSNusZhXB9pbha+95zFG8GoFo24ligAGE+ER
cRvSeZ2sIUlPxdsMUJyjtNGtV/L1f0d44tkLNlHXhaGX6uF4SKgVEbvjPiVzn389
bWhvlwmzSX3T4zh/0I5oxYMw2wjq9qgZZGA1p75pTM+KG8NbbFV3k/G4+Qu5H7x5
4CZdvo5/k+VacB9cj7vtzYkFl6RWiDUE004zxdDNgQz5IMrSLX9IF0ytLF9fS8rH
1gwsDb5DJ6My+qUJJLs2g7KBqIBcAXhivtPpi1ZVymx71/YzsgEKZX8rGxncn7ix
slAcsHwGtP7ypZUyrzh8sB2Yqo7BFzmvKHK08wnF9GSe6c5fyXQUFgwQLZiIJRGT
1bW166qiCAFcU0BMA5xJ1jgs7sZhOMrMzaFWog9k26QMGWVEm+W5SMv7mE2GcIqd
PdjPq/rII7L3MeefO0bhcE+NVlK1G3CSF/NW9o/87Tmzfk79eJnrUuYpdtt7zGGh
S4TJUpnXpJcJjMtYxEVmCNa+0Zn9ORR0kH3DVvMqmB9fKahJtikWBJ0Tzn65Dfpj
rZi74D4nbg+1ABCcUmgl8Pf9+K0Ha/AhXmDwbLEREQClfOnuNe07T9tsXpJ9FZCc
jwYscu9JyqRKClzFGDSbsv9lACBXh6MrL8QrwEPfskZBwvPq/GYGBaxCdZV8KNC9
dqLgVNNw0SVjMXYR3gFp7CdP6svsWLlf52Ta4AHpHbcAxpK/9oDNmRhM9uOHjrcu
+Cw8vfaYOKFdzB/CTu47lLEyvq5FLHIEI8j+yj+uM8onFipGm351lzgIRjAvwWgU
UcUW1xkAf7S2fokvalI9Cbbj9m/cLnBjWPTVq/1a1xCij7vQXqmkwlT0X4DA7RxE
S92UXLZjr6hyc4JSGGPV/xqrWGM3I4hIl1NOwyLzn0qLmJ8uxD9K34SSu1rUVMxA
paMlaJJj4qtQIQ/A1mCEyxpDFb7MzBZUYv8HHR5l0hIxSFMz+fsAq/3S8arAo/T7
e7LWeG6PUqd+W5RKJ4L5WMiN2bFT0QrVWfdGL8a7Nc6GvF+bO/LGGNLp6vdAzMN2
gDJnQHf0pxOH4Ch6DJ5nXJqzGd3Iy/XVjmSZqxGI9VNc90foCyb8wkASpkMDaBF4
cjHxSS90mypPwL0oohfLDmEr77r3KTIVoV+kTvwx2T5JP8lGCmUrhHF+tGbLlHYE
Bq+nLi9fqTItLxnXTUaB9IvbE6k2x/j873Ff7wtWKliRwa68hDXYB35FkmoRy+CY
GJ4gqVxlha6s+0Wdyc3TNrl3TOpRiOg8iZeUqwybwry1TmR6HuJ3etgH5ft3NqoX
w8X7utZJwZL1eCq+pK2rAncPbufmCLuUY1TNua3vB7gtRjfJB7h5z/igW+Y038BU
LezJG3aEoC5Yv7FPqG9+CHelFBRDLf1xj4+Gi9uFKTFKXXiavqOV5Ry5Qynj5oq5
8fadMvszsQu4vt6P+qEvN1lLp7UI8r6uYnbukvvLQqkJVPZKvUkVu/61RN33gpJ2
OkTwsG84VSYBilLDPmynW8VmchfKSi4a1joy2Ia/uETNhqNSguxx3+tm0Qx+NKzo
6imsiZk0lwfweEYw4ErzoJby314yQ/sK1gOvevdor0lEZVMAZFBwfGpWHQ7M56se
97HoNmuTf/EeP0C/bw01o5rs5S5zGNrs2zHRh494Iv3Yj5/1dMP1EZ3pPzPc7z1v
9F39Y8xXReUK+DKbA9nV81MByQFmvNhHZ5ZMEiVBE4vjL6u5W7WvujDFrJO0tU2B
RPV9PDuQR6fMbYtgDel5blpccDSEmWAy2AYtRat40AAuQlNDT63HNuNRlHGEyw8z
+mXZMnv2RwTPnUYIs63DM1sbShLTlL01hC1rQbW8iKrE9XPdcd4u3shAnYCcgE5O
wmRbm0DUUTcSTUktO5hUeSXkXiZzb9zg4VGQejaEnL9B1Bs2Q+1tTvBmtDJppwKb
8ip38QhonmhqoN81GekbLTHlRbRwLFd+TJFMb9YilMj//wH3MAqAjY3vlGqxUwCt
AIm3w8p+Y2m3lUYPMXw5duPj1DQ96qe0HKgXAcqiXDK/XQou8q5LJas3Z1avNhPO
E72GbW4EYdKbVAT5MR27W98cJn+FuhT6mBfVkTHSSnn/6R23vs8gD/QvhBH6FV5S
8eNW63Yp9AANxPNBFeVnZh3ZUZSMerCTyA/oEM/slGOOJswKiATqyTz1BXq3kJ0d
H/uZAj8yhYs0W3TuppcfiNaiiTd4PPRfrqM2RkjOhLePLjG/l9wgs1sqOlH3/HaK
n2CzZzIrVWFSKnHHX2PFR0bc84b2bZb4Xi3BC9M00FQXwODXyIUKhFR+0q9FhdeP
3pagJoPLZB+/ui2jJ4OPLKPDxHQCB/x1vVYS57Y0PHyw7D1J/zH5+TkNQPbDdnzI
0KMCaHi9cAU4ENFzrnFo6FmuuYgRdt7TxivTA5IVLpNY4ru0yiOzr5rDjV4i5YTg
QPuVEROaPlR6bP9BuKQIjFmuevr9nbITidin5T2QpYXglULTWWMDFxLlrpXN89OX
7XN0kYb2U+nVaOLLxvyrH1NCGVRkAcD07seAsRa7vqJhKdhvwpjVdxjQN/7xKIHc
Y5YaFYWUAOD3zzYR6sbpOdrWqlYeOJT6wqaqgwzmK0oO+kSM5DUXAEli+mxccILO
lnIsvZ27h1frguFFgL2T4+t0qiVOIWpTx9DCDButohK681/4N5ac9w1HzgijUGyV
1bNlqtuMPxH0aWZAlO4JPVqVqGBw0PpFLitdzWlpkYmmnLYFKpZ3vTAjZCNU68lE
1HdIKRSHZ2PzwzOo5VIuk6IS8368jCNP7qgBwCXjVrjQHzG+NExzW4PXivp8B4v+
J9PPpv9qb1OFP7ghQzbHOjpru7Q6lF5Ga09EFUfSWki+SovqwxQUbOdoMa5WTCzy
u7R6D92AGFQnstr5j9Ch925Z6XXwQMCPQOE4Y7cv/MlO8UDqA1tzTEMppo+mUc5N
5BwVrW8Q8DOaRXEtJ8MJ7Yc7o1ugLMuu7siCBiEV9s87/xwOGSG3EL7BmQQsaI1r
hsVWEuQB1kp6zmSKiXOl+xpbBo8g3EhR2SrOxwVbhCQG92PPmH+0E1PlzkQpp4G6
mTVPFKEgWPpwY+7vrxf95bdz5kJC/tM4dFx44xexr+mv6qQtEjp2ohEl9PA4YBed
3/E22R3ZGJcR7x5e4roTQPHVFsYbBnjmxAKdiVmb8eSFbf3QcP6QIHQBVr5Vmb0+
++a9PgSimAlvmq7iYN2D0hcRWoftkDeAHZ9LU9y+IWHAEhXFQVVBbU0s/0LNei5d
LHtFTzz35zs9YOq13IryrvqPuSnw6Ubfembpk5Z7KoWkk2FzAOTmFSpn3VHQ28rf
b+GABHfVJ/7VQOoYtc8sPcSRq7Ixs010F8hOS7xX7zkdMHyn7PU+9AhIVGKMPyOx
07DGCt9w7HTBaZf/R00QMhDW89WcAyMg0S6IcfmUYe6thMpGrVeHcRPhqSjMKnXZ
OdjLw9Awe173zBbP7iMzuzqI0zu5ZBOYR/1m2w4+5nxSX3owcZVkz7z9GjmlBk9u
x7Wv92pznQp58yYO2YmsfAlHlhdkCEAsLiVr+xaHqKUBgqh1m8VOU17S4f7DaT25
lk3kTMOuZdbUk06N32Fr3u0IGdswWphctAYDTpQalUGyKsWfEziKocdWjEA7fTkQ
UXJQoXJ4acibhCI1Xv5faknFzZM2jcropH53L18dFP1xcPwpskxRPsvfaDuBImgp
ffgIOxUtOXi7iguFkG+mCptETU72I2w2ivbHeKZua3XAE8bDKFqUXeWozFkBa9ew
TD3mSQNZU2xThn/ncwjDPDnOaQvmHxdhn+SfS25Z5LRnpMRvB9K0SSop/9lDK8n9
9F4Y3P1rppACHhXG3uW9HYiFPwY4ipIhnRLV7J6ky0rlu6ojjdiyo5j2Qy7aUBsL
1x7ObaqUMTbI2J5ffdiyoDUnXcapscwUCXLbU+XlAz/XMQrWKu4Dn6r+w5EZiboN
IcUFnAI+3vPKLavHl+pb6srUguxq5KO0nJqGh263WzSnF+GcafexI1bI8BvmyzCN
s3oxw4e9OGaV3ar57kPitXR9l3cFQuq7XXMfgop1+q6qRhBRliBOXc3by2M7uGwx
0dMe6WMXtMAEy3AzNMaE/8+1zEe/+t+dB8seKpvY2/hST+nC3vZT6N2pojgTbums
25WE28G/+93qoeV8QGTnvU9zgeKcOxuurVC10QKEGnNusbTblrvtjdre0YGhBqVo
Uu1vrQDcYVxL+FIw7DYF1F6iiut1SJ7yGDezJwG3lWKprg3dXvRA+X9VF6Nj2awz
2lteU9XryY3xgJNsJhqz7PTsy5KTKyJLfoH1CBU64S5u2TIwZcsa7p3rbNJLuBbV
VlnRzFKvU95GZOEVInClupgBvIfaka4WWp+m830Q1LdHGWX0BWqfa0g+8qbYSQAE
CGKZIfSoIBv992q9/PXlEDTBsoLcQbss7jasjPCw/mB8erBporGfmiSa5TDen1c6
OWO5R/FrKmSS2+AuS4hu8gWc9bbIafpSdz4dO01jL+f2NSstjAaheBYdXb35I1PZ
v9t9RHq+STnSgL65HnyKFeJ6bNb+hoMgHhik+TSmYP2MYVD4FYk9TwlTq93gJWcj
MjbFhkbJ/IsTrdg8OOWM3PtPanV8qL2KVzfCGhbQP2po0oUJTGLUcLr0GvrmOWp2
r5693VMT0CG+VeV+5y+NEPvTVXr4CRpdfpOOVrPRhYlkiZ2pca7lFbV8ArMTChOm
CyDIrFWgWYkpAUHhpJ9ZxRNvI/oAHv4IduYrDDYcPNTRDnx3sZO2J05RwrA2Ck+e
X+pweuQZBI7xDGNl18skY1QfaJxcvMifO+7FL1TikyOb/Lv6CEPvDFPbgVfeL/qq
agRaKlGmLHjP8LVzR22+bjMt4LGTapj1g41Q+7jXBQKv5UtlwmoMEi+nPyAAPzDo
Frc9IFP7Nqpo6xNvcdF4JgWwE7SriDn1a0oaoHVUoKWAVWwwEHXHY6HgIky6NFzw
ZyRRA+pw3DUKRB+LYRh/nsdatfXwnHAhfHUcdtXnJTGJIVjcxHCfZeIOEW7W3DRl
TTbXejucQJM/Bp1L0kk7h8EK7zCoa22cv6hNcye+5h9/vu9+MArkT6JqEi5em0/z
wEq+2F7IFX50QAPr36zw4NsmrHRt0uC7I6HMs74ox0pTYbfMUrnHoTPbrvVDn7mc
ncIIiSfBbjy2cOi5kuzeA+O3Mr/rwlbiUSXe0n57AISPPC64JJwBsZaF4R2ptUwe
07P7EKyIoTPQkO0lbrOFtDi04bWyb3OUl6B6sHmnum0H1Rh64yr6qM0vZdAIVQWJ
DfwLkEvjD5NMJxvKq7AkYZSeXXhegXmyRW/Ck0sjdkSZHXfo2YGWI4z6zVgDbAWL
Ku4510szJDngaE15HYzTa9aO9ta4bZqN3o5Pjs2pGaPm0tiJc4F7AMEsdzUZTxGY
EASUzpMkKsLUv2Si2nSU7V/NBguY931oPP43Y3UY0VErjBX1eUsakXd4Ng9uyKra
9KFUL+rcTtj4378WayId57ePbi0MjSpCMqXib8vTvux0ZcCaNbIjZTzVJXd75Gzd
CmW4653vTb5foF6p9799uIr4nQVrrec+UPmDy7qeMgNWvqh/O00vIPNe6+Oc3cU7
Z3mQ8YdayUT66mA7y1yF236yvlCM1nAno6927f/18hodtae22Ed1jj70lNQte/JZ
2XTdSmFKuC4omrfjL+qh0Y/62l1vB5v44EY1XNIlkUkr1uLbkEPzwXg42GrpCSCZ
4L/ROwu6cDrWlz5liPOVq4jSdOyVeSEld4Xyg64IdQr7YVx5usoDCS8SOi1Utkwm
nrcSS386u13BBSsh2uBJzJVAy4L+di5lu6KEklEE02qPOkZ5i8XrgdYkt+QcY2WO
kiCpd53Wn88GbMX3+JqGOP7kw09WpgKMjnT84PxQn2AYqf0ZJsoBlyyL3DxJyLGQ
m5eCIx+BkchFZNMff4FmADIyYee3L0RgyIsrW4qFtBCkORh2boniQ39ZfyCtoJfQ
j7BeZtow4ypomfhO+EJLUytxnLNLFuOmLUOay06CvPXrPgtzmDLkWNcxcbjbXcKw
Gk8HBbtEcE+zaUpOKY/P8IhIxbWXVz/GTs0sJzAuYF6IJ7CRI+ifqHVWYNyBWszF
j15INTbcLhV9N0mJJxlY8sBGBupCzy6+CGo9G3pu8G3u5Bc2QrzqkI7D7z0PiB8W
0xt6S1oCok5d09vbGxd8Y20sBKVgJtwn2s0AefJ/wbR59CG1cjlHD/dxg07f/Ruy
afMtQnd/kfrWLWjBfUG1DGJGI/xbXyeCow56ZjJHVkrD2muy+qfaJJYgQSH3/uaT
bL2ZqkqqU9tZEcCWdNkVWB4oN8yAgM5dlLFFIRd28ggxUkB4VaMQVStQjXHlIcZ9
ZAr1W8TIHXuV4lxvtDbEUdS4HPli9kvhx4Xe9dgkmP7zf5Ol3iVLP9PSeQUEgKtI
mz9fhAw75aOy16ciOU9Df0pTEyoCY2dnysRFTRqiIClbLeOQDDD6zlsrohYmL2dG
lVkMaBZoLKgV6wGg/2QS84s2Rnk0h6B3ZkWIHA85FVRiZfXIgw3IdMtYgCTpUweI
4QJGAk8PuvAaOrLy8p2kN0fHki4qDBnOTfvl1geZqZkxWQzkkiEoppgshj8dipmF
Yo9jUz/9qz73wA8snagVHKE0vzlF62bHQXVitPputGJtarhK4/qSh5SeWqa8Je8h
WRQOa6qfJrwM3d0vrB0m74YDqLm+qu9grM7Yeo49XRxNKmoT9ZcUTCLI4dpVCbDa
t6u9ZPhD2WYokukZkrO2NxXEnyamDZIE1vHF9sGRI8PhSpHl1J7m4xRh5AtBqEV7
afGrFRGmuHSodV7Auc09r9KXYB6NJzwyKavDzxH7eRvz1AtCJqOfCfzHBM0nzYM+
kMzYuNU+bt/zuzrcZbabhi50A//k0fe0vBOTz1WF/bT0KaQTW/p4xfjIbhmrBk7p
vEpuikXVnKd6Y0+buUy3pR3En5QmcSj5oHsZUmNMHTE5Qu4v+INZgseP2zUleXNo
ng2nYOoVH8ucw/rePa+g5qFTBMPsAKJ0RH8+T5iPf3vWJS3uFvJnTbai+6+hOAC5
xyXxEnF6N9w/qL5/a9XrtvywT6QTyAmoplt/CIXJBy1EJurnElz1KveH5jpMl947
cwD5dVA9zQIkiPKhgETMBDegzY1Z2HZTVxek/7mz0jOZlHOpDX7rhaYACYzhojLi
mWYs3OxRT7lH3H/OAh9ZtAq6oP2Dv+X7+vgWOQFI2M+rXNQatEkmwKoLCyNRPo59
MxkNS+bQ4VaW6Ws1qO+e/H4Ail/Hz4KppQUnIayGh4IaZSuwcW9S8lnWQDnlJjxp
atGUEGC6BDMACcKnWLNEQNP9/qGCoqx5NrlCpqbVaMk7lgC6R0tt2pTazsJazeLw
aa4eefKJd0ddfdutoiGbJRVlJk8YW1BLc5zKihJUmtV6wJuBh49xO/zay9hNzJ2V
gmqGRe9Jqh7BQCYGYCJBKgcD6JFHkrIiU6IAinej6iIFOdZyRPDMwAB8gEhOwkkV
qOScQ52npNLaZidqKfdOzeR0DpJ6XdJL6yLnKTPL94a6KZ0M//pMo5OMcgvryXK2
4R9eptA+pZHF8S2j2LhL+6Ne9PBmGxDkp11K+4wFQGG/F53bHCARW1GNBbCFAtS6
GY6RXhJAXIMjrqlottNLR7ZFnYGw2lHWdIMJu5IKL9SsIMQhdhZOdjOFVa14yeoB
KcfUraqFo8HUCISjnZ0Kbr62vAc6UZmQ0S9vgik/MrBYaxQCgO6Z2xnSruPDpyQD
leIfb43OHiLounPTdY0XDw+y0GNLqMTFU6TLlM9yLYk72Rt6x9Gxq5Uwg3ETJdYg
2TSsuhxDYpEOmNBuFdViOCR6KJtEqlwqhIUs66ario7x5xdUs/lVs+Ei+atJ+UOZ
2F8S/eAVg3YuI8NlnIqEreCEMlate/flnL5DThaz0Pa452IkXyukeg3NDMBVwLJH
j+iIXRPNaBypF+oOoQqF5YTu+9wO3tPsBrUvEPvtStEBiy6uUumJyyoNB2NlD6QT
v8o80AlGTmbtFrLO3PAyfONwvLWqID09VkSGMJSpf0Dum/P/wCINxFzUBhfGDXn1
GKjbLKa+7hx7+0a2VmJXaUGbRkYWnWl3pZetHoy0uOQpkhafjH9+AXI8fxi6vLkb
1O5TELeYPoB9C6ewO5dU6QyijbsYkjxrjnGWRqe9pB4ZzsFj9DuNVwIQurI99jFG
zuY0GFGjyLZ54syN7AFL+5OfU3XJxvzxq7WU4oppewMntZv+k9Zk8Qeh9axE8TVD
qfIVhki0v6ToZa/5sPNwd4N4zyqP4xe8geRjuiggCCXJdfQR/0moBN8QMkMFNr9J
xiL+csXvenqSeYNW8LvVMvdrniLI2Yk8OG7zTTloDSAFtx5zNq5mNDEZ+81NVOx2
GDXiMXuimFjhHMvkEJTKhy8h7mW8z/7uc7tbcIiJveBSdlfpErDY9TKN1ZCKd0JB
N20m9nI3FSbp2UomuBFV7SKSUp+91NJR4n2k5oxzxKktzZCxb5ho6p8a0raj+nze
8kv9WwwYyOzvUlv6uIp8bZqEwAHX1TEKuO3N+8fd7RSWDks/dXTEQSzs2x8nDuWM
OSuqvKNzl72idxoANWHXJ93efwFES7lwEinUpAh0qO6tQh3S2HOafBk8YrmClOnF
LbLSG5NwehO1juUTzs7VPSkUCZBl1V6dcuwtiBIROt82mt6xoT834Awk0zbzOPaW
N8oV2KHlgrYPPjC9WblDPCQ0EUNfTGPbZq/oqCWy735g9S03Ru7zclb2H7lqI7wH
AbTM+/8Zr94k9RjwP+65nZGll5s28U3MyMkdCPutlCchXlE3nHzPdju3bmjyB6Kl
F4iuCpHoirRy5JK2k+Yf7B+3G2shuv+lGeIvWgmNwsF7NEK1b3bMzgUZ3HgKhwB6
eSSSaCYP2pDOZaZVMzae8YIpPKd1hbRcL84RorQTeJqNpiTRWt/SmmhIqDXILl6K
Dy6HS79ChgzfQFaGtihDI64SG/uiEl0CIyIMprvuwM6y59OwGmIgSy0IPZGXEFDu
SLlZ64QKW5nPlRlTsgX2IDNPwimr0VDMnd90IMFhf5NzKnUmdpwC8XuQnnpPR845
ghx3Nn13ZLOvV222VD+ZsqY2toANt1L3hdxrA4PfZK5C8mqjbzC19O58xOITj5f4
ufWQWTJG+XiVRG6ZgOCV2NIplMe9YJXHIChsSg6/GQDjiaLF9DkKyhJlKKSYuw2B
AmqCXU8UIDSDIHIkY1JIXX+nZFxSSPoZ5/x7o5YLHKx0vmfcbQuF0s+p41D5u8Sf
J0noDKLzYcj2f/N6x1gBRgq14ficT1RKgTE73UpX5nHP0Bl909ghw+oUiiyOnM9j
yisUymXDTbZV9wtrNW0FZlN67s/GfQhHOIurPz5UT3d9aXf+YulkZnDrBDeGU779
3QfKFjYn5icLaqrKHc8GCwwCjs+6H8IfiZFwwFUAkzMVXmdb+LM6eUUQhUNgxhPH
zbs/oJWaEOhGObxplfHPIqtD+S8QoxtpFIKTqEuFb2JVZdPGw+ZwmGI3IfWEe0OA
Ntdkhj9XMmIkmQzZSqMFLj9kDtTBHFMuM8p01EdI9DRtIG05SIYtWvg2iBS7cVWc
FX/8g8pGLDMv6s/b3oZLdMFzMdsBUrzBZwmWyWtpPApBe/scC0PLlM/4BGMEtse8
EI9R/AW6LJDSEvkmkEHG8gyD77wUm/LI2McgP4WvoYAomtWEcjii1Q0n8AZoGePJ
8iShWoeAX2qyqDHcSyp55jIrAYdRIoKaTqZ1kn74dTeaaCK24rN6xMRRUTz+47Ir
NxiFGqdMauScvblOXDN3F8MprGhmHENpDJ33yVkj0KFrMHeiMYhi3RegW7RGy8Fa
C9Cx9BObdFAhnf7ZPXdu8baGNQy5w5Ibw/yMwrA2JyWv6x55pdTYAxnjf4tiCwoe
6HgEpNuzr7zfcP6U+kA8PnWYJBmO97/Auwxb5A7/r33UuUyQNTfL03+WFAH2V7C1
Zf2lmFmqyWxoachdEjqeybBtIz/ulPxl8PLEtAcrVEXYTspfmmFGOgfJSYx9aDCk
Hbv4DRKl5D5tCrUttCDA0Gp0PstDDUd10iNsCCNDvATnUpAakNEi2p5WAGEGJSzp
fXybTFRFbId9muU7XmBx0u+MGRL52K2+807grdx/cdqMAU1ko+LlqflW3/OGh728
QrZaaORrF5ER4TH9DbZmbrlJxQoCkqv9QvvZFauGxcH/4SJef4u0eJuWbxGecdGo
yNDFQYJdTXamV0PN7iqoEnWwMzPFHTxB990RmFTfZjt264G2rJbNan3MM+07YyMj
fiHJyn8a6SNNUzPliG+ghjevrWlk+UgPHhMu+ucVLa2l3nEpFr2TiKzbc8+d8K7m
lTnFOEFnswuxetZaOhjsMX05EGvS1QDnr7nA1XdvQLGYi+6cX1eBxECZBhx/zGKZ
NSjUzb7U/3C2S81KoWLeMj4jSag7tsmmmWWcdW3J3V7DjsSx0ecbgB8QXJbimMht
2QYu2YW+8XU6+HeX67XsVLNSztSo2Csu/08wNVhldyClTphuEgDF0Dt0r0UxIkRH
iuHSr2ktHPKNSH2yu+4RFEHIXih029K3NNA9piizaNd0+2xHQMrYOGN7RhNp3FZ3
dAzspmYqETeW9ylSlnPozTRvN9Bdu8p8rW3ymK93SfUa9l5ndYGQ/ccc7ELfcxBL
LCMwzNX25l66T2K+Q7CGVKko/YmITMqtp1COOZlM/WUlsO6WZotR7a81KBy+62fw
uXGqp2rmZjP7wbUW492vjgsnHkTU9oD6NiYH3jjI5EYmi9s7OieKFqyDc+oEJ8Sw
i5gApsEVbwrOuTMteBw697++FxgHe7wY+jYvtD9t7RKRyDPRWL6UiOFZvxPYA4DL
DmrRMwn7IC1Z4PCXx/JG2AzgAUjTpa5gWimNWPUM4QqGO+rAuudxZLXiQNq7Oxe6
rRPT7DY7DAiEEI58r4hiHjJpNhPJUYjPLbzGZ2aTTy3+tYjxKDi9s/6OEMA3kerI
KAuhy3+vDXK9PWyXAiQzXuOuua+KjDfZI7RF94XJjwpWRFx5WMiTqFvM+trDggI7
Tb78U4qUl0pX2QduZIJH4ExmBBo4loudaF13SzemDa+VPK0VyUaVOoFGmRyMFog1
t0zU/JaDNH7p3liLnZD9pxPcSlb07kym1vdgOHL1LYrozMaCOG1qOWEWf6p8UDL+
3kXIL+b4gB872jXhnZN+1dxb1sOhzJBTVWoVkxNU6DAdBLkJXZkQRlprIYWjypyi
Ol2ZjfVkd+xjDrl0/JAFsSsJNVOP/J4IjN/AE8QCwjITE714RxsuV5dO2V+lJbIT
4B+AbHEuovPk6zclPDBROJti7u9i0/tyZl5fxYIsW7GJfskbKHMnkmsIGw2P7syT
EONjQj2E+d+PK71NzjYhzaCuxgI6rjXFXZNbtojjPcIAnpfaw5wBAWfz888lLKA3
gsAxX3gj5O1OzYerfHXuD1Utf/7i9panPrX5YumDqlDL0oKdvShgqXhj07u7tas7
7Rz07gqzV87TH8iaRv4kESCAdLkjaV4aNr6BNVZ8//ffSgCUy9nc7V2UfqgnLaOA
Z1PX65izA71jXpxTYWNJXlWW9/7J+a0CkUzT5CvomYR6r+Y0TG20DPGKTiGicFzc
04DQtfGFmoyS1kukDcceIjLnmmRGQwhow/OEo2RS2ylukN0MkQbtLopmLPCD+qQW
1pBLIHHK3vbdx2WwFTTdAcdr5i/vuHA5X39GNc5MfQLp5Op2WfS7HcfEO41ofubY
P/b5JMgq35yNGcXQxc4Dv//Zol1T/dzeUgzSsWrAZUganq7Hkz+TYKVLJn7w88sc
9EL1BdnLQ3wGBbCF+1E+TJ5ZK3hHYxhwFmmVQqRiZKkrkezT+f8jbd40q0/Qf85b
5yGmpz+BM/FTgNlOSZLlwhfbr6roJv0BPLwYFaawSXAwKGZQR7FVSa8zOqmYTB6C
GJobXVtYg/VfgjZwI02RcjJNb3hLAy9QZHQopjfPgVfjy/fM2CO1Mq4RiVtTHD4v
P9zpEekzEJce0piZqNSDfN1B2SSzTBlZ9957mmdIcxLOYD66IUV0hx2XZg01VmRi
4rMVT4cjFUmYhV0styCNAiwL940LtW8SD+rC4yV1oLkH0cVDd3gMvQzzeadj/O33
w68K8pLXp5bfaeI1qWZFMPq/Kx8YjgjiVzZJ9LHXA2V+85ahqhy1mOh3h9gY8KT0
jort/etK3nrmyvO9YFutivd2xDnXPcMwd9W7/4EFmcFU/aycGniD0c4/0JNJSJFL
fh8gXI58KYrecebCFRRrm1cSto5kP+S86OqqP+8qtKtir3GRXn/rs9et823osLtw
t4Un2Kcr2yGzA+pfrjzIOPVf7puVidpzkvpQJR9/22sKOH/ZYVUfLT6+gU7I1qFF
Joyj7VGPvMh1k6xLrEbXXVpH47qRa7EBsN4Jhk7tf8Q2rG1XewzG9Itp9sN8Wd8c
zgu0upjiwrrsUIFhL1Ajb4nAeFJuMXsVxD3xM7wkcuU24hhL/BwsQHgT24vg6M/J
VyZCYDm7B13N0j+pk/4vupvV/iN4ijyXzbCdAvosV16RPx5q/QI7mP3QC1niVKG0
Xp/hgm9cg7NLG+oBW5/Zch5BmsIKUxzajilAipVSMoUULgv7RAonEyZihrfEas/0
kIsZJwQzLoZ4s62GXr91L2x3UGvr/ZmbZiSMIfwUp0/tc2/JQgeJXzgbiKu27nZT
V8Q6mF5YDhadg8bpJVDqbzqv1U5v4ZZbfSC2JqNFn+taaHSXnWfDy169ildPLRKk
IK0IAigrG6d0EdSrQQbD5r9TIGQBluzqO1teH8CmBOSKnx19eZ6+bO/7aS6o8OMQ
0tFT4T4IHAyabyQaJUmEVJbDp5XVAVn3EEVxE2jWIbnSsDV49TcHjWhusYDSy1Rr
SwcL04kNlx3LjVKF+7DRWRn9oNOGFWjQkO3ypivLLuY=
`protect END_PROTECTED
