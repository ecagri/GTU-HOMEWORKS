`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V20hd9QfEo+l5BUqARTGJJ69SQPHRdTpD3EK/lkDOyCM0wQ8qdCV87VWuckXM+q0
qrBH6DMGOyziAhHXduYU6+T3YMa70gEColVod4T53V25dsb22iFxX2vHKJa5XSdT
TMPHzT7EyCDMyR0aIWJbQ0tOFDJSjXJcj+0t6LKea3JxPMk7bWDttEALKBMgTkhk
hNWd+XTwK48bk4yqVOCAf+2mz+bHTZtxNa8N3Nz4ychtB1XosmoTULqvWP4xkCpZ
GU2BJC4NIKuq4MYcvB39D/YPnnuV7Rw6rkNsm5g368CBeeJEhZ562HqeUGExfJ73
1I/c/ksGvXo7zvGqANNy4UUMKweHVyucJIyE7cL2CzLH11WFQ3IQCUk/jGSrRXuA
H6SxkKDYWeDAn+o9H3/2l2tQVJV1FnCTr+ehzZUuROgRcXAqMc3x/LigZKxArBLw
nJM++xcGeInUWleV2PabjIQbDpqMhBR6TSrKx7cyUH6Ars3ujidF5XFWg2ntAq8Q
MHQ5GUwcPZuTBciPmHF79DvzmFLR3k/pxFgmv21eKqtMW1434TG8WDTP/uprVI0Y
xO3R7F0F+io17i0JZv2RBu3gKMV+Z2zpiK4BWe+fLHMOT2ZeGkizzhQREZL84nHM
BdzvzzQfHKwrhhjYuKKD9nB74Jus6jn7NTkBgxCm4ILLjR6JgIXg0TTQSNRdjmMw
hihzfWI5wGSAIdOW2T1UBzfyo/goaVy1bHlMI6vZFRA5q2Cd5G8x2AB+SjGS3XXW
oDre8A+MLWiKW9OWN/LBwjdpr6YpGbHDW9ApVijzcJ5YSbThsr8Icul4Mxpw5PmN
yP69A6rH57z+erEuWF6Qhetuk9ZJvAvukj2LYCRUMnylHKev/92gn9MJjbklqrin
NiTaJRuVLfUxNDDV7A78wXZaOb1BFkNqHvxwjTA8anblY4M1c7odBoW9i2F19KEw
zx4aM0V0zmitofvUBljePHZXCUAjN4Fk8J0gzqLCUt6IlQaMQ6PFpkDn0mnB5GtK
MIvn3ktclUXV0Cp1RIc1EfcL3WW2WGvOTHZrSLjYAgqJ+Mnm497IV4DEKuqiVBw8
kTEQF7WcBut5+DgWHHMN3aR1hLrDKu9yrWufq0nYS+BYOdapClrnYdlQRLe/WVLz
epj3h1AJJCltzxTSLcuzymVghzYRV3e2hdhKTedwhpnW+MO+fSC8d4VW0ccxryX9
BPiKc1W5T7z0vxC+YvJE6zcvMFwu2Sher/dmpGPaFvEH1JhkeTOg+wybzLCBXcG8
ZY/XeJRfu8+WQQvq6V/vAJ5hEEGUmyo1pNIWVCZPV+JiepfJNUhAjgFhJiguDuj5
mRQEiy8Yj9l4mnYbhffmGqcH24NNuQJnDxJlNioiw0qMx+VmE/J4kwIfYTvD+6qj
h0nzLsRcPlZJVMQCTN8xFcJOy2KUrGHEjl8pESwOm93mCrUBl0D8Ext+vVspeEUW
CQvTwH4giES9uJoooY9qYhFz9NWosTNgWOJVYk4PlYwe2Uc2GFeLMuY2pjIsBMLg
xy5dc8gpCizjFZr5pjIbONVJOXUuCY8s6La2TND7xgw1Zd4xwA4fjDU7G9Ve6y5O
WeQORZvJHMBtMUNw80ihg5mh9eO1Me9Sa5WdNmVe7t7xiQd3M4DCIMz8dQHhBNni
`protect END_PROTECTED
