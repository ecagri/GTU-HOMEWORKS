`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ImpHeFfe5yNHIhxINUtGKGxDsuvCsOaSCkSojUGYNOOwFXKM9BJP1tqrCHhwPIHB
7Z+nskDgGy1/ZatV2AG1MV+LGgj9wZZSGAXG1FtADaFNoeRY3eBI47cl8gaqPRSD
jL9ZhFreprRUzNLjT8iiYtIi0rM4p18Fdru3jNq7R6FKKZa2HIia8CRjh2wppSba
vLKLbk1dmYQyae3Kvz2UD4Y4mybeR151F6gBNHPg1LpMX3RGHyi/bbcc5tR1kS6i
sjolHVdCSYh5q6EhPuEdYl8/lxBGy/a2cx8ARsafqgzC3K050N9Y9enuw6P2yz3Z
4gjt6EwDogVVpDvlXNFfXj0Imb0Gdb+VFCzWtqoshTtWzSlWcr9u46tx5QkdlG1E
CvcGhA7wZGjeOiEH7CKloc32U5noRYrzS8fOc7LmMOsC7Z4wxPF9O8BxUxbaxHBd
ugJHIwkFFPLuSzAZX9WYeM5i7ubNaI3yoOY3OlUJ5YEQspOPa66FMg9BogmigdeZ
DCCja3OiGhPAX4KUXJkYhPHdq0QcbYv3PnraRUS0jiZMWYs/c4E9VlHNZt5gRXtz
X9Nf95vohCbsi2cCRLnkY9XaJeyZD7e9Xl6V1taZYIAKAm5szMCCK16/HI0dRJGk
hJNkHIcyJ9BgEndC/svhkLEPMztFTeJ/UBnACwxmcBlqlIzPDWyo/9/nszmQL+D+
/wiiJFS+UqCC5u6CdxaODqYUdQfsSeGKWvcjHAi5za0O7qSP1/S6/MiH3tlyFjQR
QgTpPT5SOlzLlIjcJqsXRnhRDSV7zyIM0VOlGUgExzd3M00VxX9GjtisqCXMDc6G
nZMnPJNX773gXmAygPgNy1Wk5/iNrviZRDyLqzeAgPlghkDdG3r00QzJauuJQ428
q9PP8NptOaKbrlrDpHAe5qdb8jDBKAwZ0i3EkzYS5rBPkClShn5AZI/kY/lU2oMq
GazFrbR1/bEeSdLmIxnOaxN7sc7eFWcX29epOmKnPsoUMKVDsGa9odmsI5bXkJZe
AUmaZWZht4SdnMYbyW1kB913K3ED1AF+LAFL5ZHgOPIKE2vkhkMnOMvi2Deuz6Bk
LTMzZ3h5tmUIsMGkNkjIqUJ0zhNCkvxnqHpBhgH7LrSEtOc1qu/pqXalRe79iRJH
Z/3HkABzXMDRl6vfEMsG6XWoXm19Mxy7Eixb1nbdr9cYifIzMukBNfk+mzpx0bg1
qxGMSSFfK6ZiOIWtFFPHeN9PqWMVkaCag8scTH+PPK/eqVEUUUvmZXRqTyWajpad
paPocz7/ILyWv4PTzEiOkcsZU50ibfDSzYTSR51cSAm6I/yQH0E7QT1OdDlTqD86
cTbdfYzVBF60huvum8tvBVHzTDz8ZpaBFMGHD/LfDQrzL1B7osmBq0tW3IyJOK3t
LUCg0PSyJ1crMpgCnU7BbWtI3pT5bMdzkTiaFspc2MB/6Y91Yxx6Jy4DZxmQgL0L
bgEmc3Rj6fMFYp4UJ/ew7hurT+X2UU/+fmmTzzjb3ceITGHx9W0gxOmgVJjfaT0R
IfnkBiFW6V24mLv8w66yhKtwx6DEe5jTnI4jqlTCOOuXFqc+YuGZJs+C34Ccg7Ci
ZhPBhM0ifXb0WFSIdvxydV3qJN6UmCMd51nV5iw8Sqt84W0+fCrhOoJbIrv0lBoy
y2u0vgHWcHYZr22YA9/6PF7t/Jm5mr4C73SafV7avaYTqlFnEg+vyrA2Gu08HKJ0
IXDaU4k+WVOGUccYHo7JSch2dbebAIKysgCYc0UzyL4aAQrT+F5Iu4cw8zltHw7U
h9AYJv4jhGxr7ex+gloMzHEMcnPV0IN18ZlbOTK4mbtl8KWtSOJlo5E3xnwuAC7U
gV1KfiCZMWmy2sYua45nj4dLDrt67DLYC5OgZo5fewOMbkVOSls8fMxrOAIUigsx
Ltkweh2foNqZqsghwtTBxXBhsIHA8Fpzo8bNuyIgwrlTjUXxOoA9t6pL/sEeZRcO
wuOT1tHdAw6KlmxjgW5Hr0/s725EV8lR6dJNpvIxCC0NDhWN4BOOYnofo0E6v+/v
P2xzAK4UvyWWcNIQeUoQmuMm0ISjBZzePrs1EJ8yxowSDqgB4OZhTE8RaWR8qlZw
OdghxHCoJIzgCFRJbAlUPmj7P/zrIBzEVd6/WcxWYDDYVE8+tnt+UgtkyGYmA+2y
64Iv50EyOWKNhH7eEKHeowQAf/RGe9FcZ/YhxhauZcj0xXc0rGtfGa/2vkYx44Fv
vpW2fJkB++iMyK7ZAFSBLWfdhGE993QkPkMFemqmi3LjF367anh907Zpn4Y45oMS
mw+FMDyHUT5CSCnZEV25aQDGQEx3lhBCrafxiuNvqOBmRXlChuHrhGddkPb7LPG3
eMPba+oA9ns7vUYNJie0rfg9yMfEr4gUgY/PPUQxQWQLUR3GpqSPhK9L1lcMkeb5
ElgVsecxM1dzNVOYBioaCkgl7TQL2Mg63u/xk1WobxwzgTM+wLRvFoSgWFK3hJ3b
JUns0UCvpjvXfplVIdM1QOl/fm895m4ACcK7k0dTZWTtonoAvLgFPN1oTzEtulAr
/hKpP3OeLsW5rf8F7sykIjre2+qSq16x66P/Jvu6Sv+sSJjSDr3on6KjRfXKDLbH
chzk2hOBjqgLBACTxkg2lPFKstgRaqSl/Ri3Nr+B4yrKxtE/pa0BUHrJ+8AQdQsI
ESDe59lFvrU1LAr3QXXeZRN2Kqlgz1k7rU26Ke6FcXaQg01UEq6O3OTyOf8VMfBh
uVsV3Eckop0OvNF7d7kNhOGRuC7OYAejYvx1rEw/gfS5FS4OC0q63snjyqahaQvd
Bilw9C1zDA7vVkxyPHH8NiwwYb7APzXgY0/wy2I5PaeHVfAA/yiNE/Y7WQRrPWdG
qqE7/PryTgBYGisSrBfs+Vwdg557yL7YQqBtwnqg6cw5ah58rA6HQ2pm4zs95f9u
ZGkPI7GzLJR3HXeOaP+p5rcMLlb/s0bSY9ZG8GVnOO1+yLYEVBnkESQtG6h08mg2
LntYziou8ZugGyRBEIXJFMlrC9Nxs4Cqbsj5BZLRAOu8IQHU4z3wpYWxrxaIi35R
rY7XNqKL3mTmCx7QWP0vU2O+ppCcoqDH796d6Ib0hDE3pEnviTvE/lkTIg52OyW9
oIWK3xp/ay0w5fu+y4YSrNJ2neZDUc8MQMEcBg71pV2BeqfDuwoqlJgIVxwWi4Bn
SJJCOUi+wiXSUSXqXoGrWSaAfNN4jGd4j7DwqFJwV1tcq8lzyrld009BLchCO8Fh
Xlyf1CCNE0bgIk5wupKh9XNhFCcHWpbuDiMsCBddUY8MFEKKNnLhYtA+8SsvzLGO
+p1q5Mv3/8jDOlTsMU5jOPTEaRGUx/A6pMMtdMEGWKGFxmCTIyDQUKeOFW0PYo5E
fHf5rHBUMEn3HcNty0ITF4iPMG1hUXIR7Xb5gQw0VIQI9voUJ/7Pf7pKdridkz5e
ycHM2N3n8dLIwIqm1oiN0VzKY4Jqj1mVjEECQXv1k4Rz7axmIAqT/ZMT4IyD3vtT
6Xa5h9F2WSsKbnzRnTovLoMhGiGCjbty2UyxhuuowOTudXI9oKeP9ARUO2ZNc8MX
8DejWSVHkmk+l1MGzm8Tfzv+P4qtilZlN+aT7Yw54y8YXCcxEPN0hs6TevrGdDh/
46B6eZ5BGhNoIjREDJUn9eENbOXz6R7qvGLPugrah059BjYpw2GO0vmjnIat+4A7
Ow05N1+zICw+qr6qTo+ra/v9Ppycd4W83klJRVmTVoeNwhPbIYy4TI6Vx8AQXexr
eKqZEbaD4wizlbbIZ0+HV6KllNcM0tlGjE4mC3DO9I4EcEsKfxMR6NB76BkOS987
xQFa7Psf50RokevS2PhWD20VkU5EjTnAsyE8rsSV7/lQHBS2BhhhUAnwZDw+wjs2
vRBN+6oxNMb06TuY8is/Q08RCbUUJVL+3Zh4GSjXNBbnoyCjhEJm+rWbaEtOeOTo
w6++1KqICq5I3OWOVPwg54QlP8vJHkyh1GcDLhFkvgL77vEL6ghpVuQkvBxno3Jh
+VDtp3IjYbQ937qRRG5WQ9vpfD/gKP+/8Ahgvefq1kiq9twkhFl440sBKGE4LocO
HJw/yqpvE7FesoGKloJJhVmh+iY2pl0IGJbk4hco/jqKI83VRiGSdOCA1fn20aCB
StBll06ugj5AQHnGFIUELbhHctGEKPQ0SRCASp47wF7g7qdYCZrsaQBih0YWpRok
LaWOHtGu//D1te3dA4ksHvsnyIgRyDJIlFBv5E9U7BrMRwqIXD6qRddRI6tDoXl8
BArJYUrPj/+aLMpJohba+vDTH4fUr6yTJrdVgeAZ/3dzTkyNA5NldgV+PV5UnRH9
NujefxrroDOIVtN7RfWamlqTbPgOyjHXefnuKmIqB1LRa7cCh2J+jTguaCkmz8XI
eRJAWGsXME8tSjGqSBDVOxUB5dRTDz8fSSggr91HJFwvqogMrUDEuWE/SvuBHcuN
3Z8vTHA4ssktbNXUW4K2c2lo10cTB6p7IRshcSeET9kxTF3Dd6ycMHzVgZghoep6
qixGKPGXRMO1rnd9Km/GalB/nVy/h4m/WEVNrOQcb9xBfL4vf1Z/2jlAZTcVxlMu
uWXrAVdxioDwzpx/si1X3XV4FmHf0bLdAUFX8jEDdeMCCEpotU9aYxIfIPbgHaui
49lXExl9lkxNnmfDO2Obg/aI6uvNgAc0z4uotWIWc64JGCo5s+EqM2oFK1TeF9c0
8new0icA70Rv1TI9t2qefq5J/P3V1wsZxsYRqDzchziBfHL4SrDbbgmy/07q94L0
bACMD0sCvR7vwSnFOHgvFUz3qFzrvxS9q/mo+1eEZnFqUt4GRlG2oDU+nXm1ynJv
BFkgkz3K8k2w0XyuWa4CDdhiF5sFAl4VaK0TOn46XC2sd9/IM+8MhdfjBtUd01EW
YCfw1Kf2evbKuYnLtBO1eueQUhu4o31HX5v0qZtr8aRxwetM2gWpcFeeAgK7vNLH
0HH+9/Q3kjKy706OHjufo8uvILzUUTTRET9bLDwa2XnCxmJOmh0PgdUtMw84bLO3
yvoYLzlqA0rlzCwE6iDYrdGYaQXReNIEc6LLK+8Odvt2tQ2X43Nl1qBOULcvx/G6
Lmq40NVy40PwwQPFmGUeCbiZB4xzgU5xJxMIk4hsFCx3ZYwsGC8026YM/zyIcPuA
vge9TGEZt4gu+/St+dBGUwMALpo2rb/RlfClipJcs26buvu+YfVZdb8fxCLqmeW3
NIHUXM162rkqYRBFCtjb49lv3wHM/myhXJVSghPzjLgIlFNGwoH45GZ9yhj1s1Ok
aHSYCzIxnI6cDKle3rDMl1t+AT+xAty3GIYjy9Q7X2Kcrm+/gePPXggZLeeGMH/Q
nnXHYGC+4RIqUMt6mrMlXdSy7mN/yJDJsDx0WOR7dh/3yj2jymND8qILj2K9AAh0
otr8cSHDFPVfc0CAo3VX1kI6gWUrTNPQBsMIaJ9oWyW5FvsaPt2JGQ1W8LjyvByV
E6Fvm85LxMxry+ku8Yu9O3/UWzYOtygprltzwS+Wv49DeO/MhXdAW+7gGVaV8/u7
rJTgoRoXvpqM4J9MOUXkQclcZptiN0ay1UeGun34nTfitf1CmAIrdkGICVFix4Ar
DOP/hIwqEle43esBHssZORGwVKRm/myiGlVeFqRMyLZY6g6GSoE0B1LslCp5y2mF
sq8LXZTFvFTnPtrMFzFq+c25hS9GDGD4cZHCFsChLbBFJHRaHNFuq16BH4Vb9n0H
aGCk6mrtXjkAscm1JAQ6UH7AGhoSaZBvnjGl3DF1GFd/mwa03yWAyaszFTGSDZjw
Ezz1D6lC1DAaQ8sBl/K4Scsa9l4pnGCs5z1IOasc6GoZ/olUy75+AXCq+fPlGS6V
FkUd5WSXx9LkQF+rFJNX04ykf9ft3o/sYBm74j69HJiw24JISUTUn184oOWiLFpP
XJ7OtgEgK05FIDmkDdmMShBO+fQOzoVPCewf/QTrHq7NuadBTurpUgE7OGE5b+MI
Wc96F6mJPMMyp78+oT/KWEsiNESi3azCm3b1nXDLnY5H7n2RjJnxeYodfGkq4Uz/
G5oZAa2JjE+cTC/w0e37QpgcGXVVnB0ng1q0TotE0NoghnN0/pOVIvUuaAr2Vd4A
ALoIXdGo13DPzqsjpiJa5582YjLeBY+1rVLIWy26LvBBdpuBOoIDHUG3m4OhbgDB
ibZGMMT6Bzd/UOZqL8CGxv9aYgR1OrgfHMSWCk/eDdgFF6NHY6Tc0zID6DaOYUO0
4DtZpDXAQArJl+txnAgPoRrmU6UE/cjzb1qU5b0cQuW3zHx28PVWRgL2p8wzIq2C
3+E7C8Nq0UAsEW+M1WjRsY2S3ReqFGmMmhTJXpIC8nfJTvmfUVhlOqZWpeHdJx16
iYeny71BSvWFDMojHU3aG73hqO+rAvKXGhbO7hSdfyyN9yKFD/OdGiqgD2jdvHt4
WKHk5t386Or7dIEycm0bZTHztTuFujEkoJcgjIt8HXjjjC9LXH9jCjLr9U0eR05q
foyJd+rgI5rYbUVbrTrkkuqUoo2JC20U2t7IUKNWxHg3zUlgjyeyJlCHOP94oN3b
TZ6mt3s0INkIkolEAFjenlIgjZqpWBV1uYDxTFJdkzCBSqQyIKQe0PiwbznfGO4Y
qhIqosOYy1aeqx7z/kLNGxQbCvzow3t8qVN3nh5fEgFC3NybVONmEDlec2El+H8Y
uslwANxLZLTaMGk+NJZTrb49Ly7ospZtOPk/aMhaQHOGSDY2/CeuJuKdt1TSnasx
0J4hsG3zobf6rtDbRzEvW0Gr624DImP0piyx4bwBKtAgoBWI8Bo/rS8KuDJarzI+
N1o5d/lbPy652Bza7kkfxTWw3Ji6VEGpqdgJFgorp1mWYOuME3S6kU1F1Rimr6rV
emmEHyaHzWtPLzS0Hq5LXsGE5Xoh1b0A4v+L+WZKtK7LB6PKOPbuWjUQRB6lmA/C
O93ok6ku8v/0p9c7LqvwMQMX4h2f5QuUTO6sib+tA2De4kojlBlMQ065DQWHGBSD
3SRJ/VNxRWcZBt+7y4Y89G9XoJFA+AplcihXjOE8vfqBad+8j1Ssz+YD4fmD/OYb
OoT3wFvhzMACbfQ2oVypDNDPXZc28+9q9PHoa66FKpsMYDVv3TLiEMApS/1zYfKC
TFfZ/2QNUoW3464Ogy2Jo9iIkBZsuX/S8a8wpFEllARvQuh+C9qOTx/5z3t1dA0Q
bMdjyicAUYgGn0psXvh8nAqm+5DkJVmr7HRA3lhwbYqb1p1hlFDD1+KZj/GmsHCT
/kma3ZIyvHjKrMxTnQtQkxXGGsbb52hx+1B6nf1c03RUSQzue2KvfgtlrVTNUKar
UrEYlkxj3Ewrdpzal1iV5jZap6jGDryK8Ny64dje0bh/0evhVrkbaMwdG2UHKS5T
SuFsKGAH7MOsK9RBtEhfxt16jBj4EWhTBUaj/4/DRACyeEVqOUwHLKL5XZj909cm
uGOC+4vFIu6p4s6b9zsAGfzQ8nuKkjQLtYQbrgPvfVs+2suQv61Yw1ARHPtTco0U
sLAfsHf1TXGVWoubGLQlnukrCsLnEVDC/SuRol1v+In9BOK8S3gMttxTWo0ixJGP
2QsRSIYQKVL+jyc2VNQ4blGq0+Qb7Z++jbwevTNHzVjrvc10z3zXNH7K3I1FJcDo
5tL/TdN6He1JdY2I9HQ7m+0FvSBxvyKjgh+mHExXMnS4bBLSJREApjMw1VhwHxur
/T/OzRyuaA3w6vJJa+HeyHy01GI2UcMbaGfHPelNTlxXRftFOPfmMFuqkBoazylC
+l6D/PAdG06cZ2Ncfrb5HhojVBuylNUGXhEq7t1TRXseCLlvZzTVbu69MNLAw3Xb
8O7le+1tq42PEitRWWWhZhQbWVPd9pFa3K1QrioBJbMkJ+LxEhkZ0aTDks4sz1it
J1ta9R8Ns2LcJm+k+ZHPaxRgabQcoeXUcVav31i8TTc6EUTf+sAFOU1NtkaI0B3x
yAD0miiFwd9kvqIS/E9StBVZcDm/LVPCfjWYAYTcoVM=
`protect END_PROTECTED
