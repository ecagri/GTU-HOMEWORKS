`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GPSwHWpgCjugFfcoJmlIl5s3ohL8MCs1keu0wvGnbQM03UgJdRcVOImwAxjaGgHN
CqG6p/k28h0QXpmH83QwzrxoXYYmJ5i4z81mW44pMSWQWHpMLgzfe3G9vuOYv6S0
2Z0ZFPumfpENtYF/OBdTVLXE/wCFz/mc8rBMw8/k6mPj/a6LyzT0QZaP05ReDXbV
QiRvL8cKACsjf0Hxz2RSPXS2y5kWZYZpnmD7NFYfeFZr6WiLi+jI0NoufsRnZ5Pq
8/UecfamHmKWI8m9I+iKiBmBKCstXqLKWFXnZbQgshb8Ra0oYJwt8/vQKjPz/HFT
v4E305JjdPkR+wzYajE3OMW2FVHDebv+2+91BbdMo5mgiKBOgh0nkYeWzLVHr9fi
1vx85qCnvzaJiRRcpaT5ofgueBRkX6QmKBVP21JFWaon3Y6f8ZxY/b99NY8qbObI
Jc8PDrZVVzN8cxLY3YvhGxLGwkgh/0p/LqT7ZbV+aKEhMXUzjDthNnR7VMjm4ll0
aEfaJxWcyqT2k2GaIjD8ya2lvaSuuDoy0cEUDX6hbTr/itCir4kysx8Hm7MMCjCi
Ie2AnrgyKctVOzaCAC2l8A==
`protect END_PROTECTED
