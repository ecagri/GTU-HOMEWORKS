`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OmhDmBpx8gz1sZOfL8BIiuBiZsubUewAINbS7zeiVCoFTvQxGGPC/fAPNUEDHdYw
HsZ9jVpbPq4dGkuTKymv7358/kZNZGFgbTh7ME25e+NhLVlQdO1ddYrYqfPudROG
tnruy29a7zi2lJcoCbGRY31dz6k/3TJbRPdOyFlqvLcOwW+q1eMs9g9ES0eHlaWg
/Zu3MZ3Nh1WYZGpTGZR4yrgPxSGtJ+HkgGeSeJfzz3qZ4lKaA3wXyuMvzMuk5uWs
CfK4lKLrLQIa1plhA3mPGPLK0pdnNGMxKSBKkEXbjFimkzI+ovreQv0+BCVxJJD+
Jn8eEpUP4omiQ645dQgbG/McXQ4Omb5fnKbHBfFDWmQiITheCc1eJD1OSjp7sPU5
1Ev8h4wA3G0Py7rVpRXXEZ6ml6dp8x05yVvHH2KFlXQ1zNZHYgibLe77bLE2S2C6
BPBcahIF89Kz9HsDy3oadEDnS6Xtc9vPQuBdcHPz7Jnhhc3edH8WSKI4/z30YEy4
GSSnx89R7Wg37Fq/BRn5tobLQIyns3c3iv5QvurHMG6x8xLKOC5JVVwD/u+Sjcm3
i20ncum0ZeOdCcPH2kXRG4leCMVdzLJebIHp7bZ0wRr45T6BtGAhueFHTMHDRwGu
AnwuJdWfxoJAyVeeIlq1TO4KaUfpAYYC3WzPMvGPRYoCuj41WwCX0C1+ZSyFYVBr
SW9i8efdYH5Xpi/6cPru+vuNcwSoVrE+7zzsDzLkyXQ6Er62r5/ygdKqNvdvTvdb
MDa04UkbEdyZ48pXhj2hz2FPebuM2gBMqQPG7+kLAdhOp6IiKpSPrTxDCE3aFblT
53gctljAQZume0FRbZoV8UgN1AF/kiK+w1h6FfmOgWg1BspxKxih/0lmz06Uxf6f
kiLECE/0wGIOJZUiV0tPwvKS5U6fVeKz6AOnOCQyHPDW8O3bzxQgH9yEe0a+gOeX
ghxNFsCU5XF+lVfCKWLFsoM8yma8c37mgNIkM6UWArEvu9be0WmRRLRTNFyxMJLO
MPEcq9GoqDpIVb2bVw+/lQqF1lMUqzzG4Wh1uqKx5GeaqdfDuU++RdwzvrJ7TeHW
MdAar+LMBXQ0JmRBQzfuJ9VeVYt8dYaZ0/fwwz3xUvxU+mtHhjKza81XrZ5jFhOk
QMtlN88CjRpKghoQaQkYOdEJuNJRUlT1Kp8K9kCj9/5739ARU49VvlaRae1ka+OM
GA4q9hd+OffMoJmqDAT3PmNBKP/dGntRuZt1/3UEwbd46OUSoCyoxkFxvHZJK+y8
`protect END_PROTECTED
