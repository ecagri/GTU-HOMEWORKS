`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WmgQ3CJlx4h5dZZC0b6wL2cpBiyBNoTYS+7X6QHMx/av9SyRLGArFslPmt07X3C/
ud6S/1uX9y6p5VQtFfid8H5LGFQQynSPp2Yp+/eaX6oMyyajzY2w7pOoXQrQltw8
57Rc34lDtizjqaBT0WLP/svpFwyHrpvbBRl+9L2BRvjg526NHKULcwJ0vf5EToCc
Pm8ztjowYjTadvpfvglZ4hwjlWIMYVHMLwIGiv192YF4E7fQYZ2zDYT3xMLC5A//
FElQ9tU9ADD78yNPbko/CdG+Y0HP7bWIDdvIg2ImwV5rzG1NofAjOPSfLlPZUnNu
GxpwjvX5O0PfZwM3u3yjFhtNFixrluKJ5G926XutDN5pZxbiwCueDiNOeIDS7lDm
zs108NAiDGHle3htbvgCk1ksT63nspY7vHr1mmM0kjN3b4qT33GZfjwCFJbUNRD/
OWDN+4hMxbYvoOI8Hv9h69SxuK7dTgojoL2OPZM9uOOX31S1avP5kntWPvNgOWj/
hnhxUrbQN0vXjmpe0NjsO1c7gEN/4lNkcet3skItl+ayS5jA1xYqKH3/vMwyk/XL
8crIU39ZGTV9WKy+Fqm6iuAJV8ZxcWyxBBRWG3JM0h0820jGiawxzFrysTv/ZPLZ
cKJLzX81ztotrcGwOTNfWRKB6DfKzJ3w4CZO7G0cDuLGfO4MmGwQ2NuJ+RMqBBso
yqXf4emiF6UEApX36koW4KNQT+sBo9qQok3ccXy5w2shj6H/DPlZHVx8S02idDr8
DS6Wj/tHvEuGdJXp3GzNb2v+iC9SJh7jWIfjqHMs/cSxC2gCdI1NBexjr/ZtHq7x
zUe47lyRF3QoGZD4Mv1hSNIxv0+A8eogB8bvBgNn+YR/mjo7AqOqUAjnJZaA/rnw
7txLmolejKxyCwdCI6pAjT/EdcH+5Jwzz7xXwt8t1OjNSUC4jghJtnW/phbkK7sp
pRiJ28uXhHjWanuqmbqe0AyCBWUP4cbX5a7bjBA19aW1DJOgJjG5ATKEVe5yaExk
kJEhro0jWQpoA1VptoAf9ZUPmBoq/6ps/puwjLBDTng=
`protect END_PROTECTED
