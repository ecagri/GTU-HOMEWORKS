`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JWFOUJfC43/sUevHbEP9d2/R/sRqWwj/69fIonALUmXOyms0+YJDs31O4wS+yL3u
F1zLLasK1wZrtjh0/LS9NRPODcyJH4At9JrPMWmXwBCa2dr38WU1bPKEUtAYj7M+
vaZjRKWtOUPibTLmf2J5WcaEKH8U1H3WgMM6Aa1oPV7qa0kVf+A+bCaOKghttwSv
QZxia0q+eaT0QSkqTnLhxQUs8rOWraVpaMemHJd5c/LNpoD6d7F8/6epRqkCGTJi
y65NptvelEbv5tm7s8f7TfNPr9ZpK9DFVQSpv9UJ63ip7T3b2RE/xJ8Kz4lU+BWw
TTdt0alYSLJDdAkFuzMkqYS2749s26vk+4/KCCEqy1R/qGI1UFiSHEFTg1XE28qh
HmDK48z+2pOB0zDR2vy81oukls+I+1CBVQtJW2rB0+4z/SrgDrKNy9giItPsMzwU
F3R3wfe80wnad3vo8BJ5+Vp/HcQhi9gOREf5UlRG6gdMELhM4z0CD0HsMrn7yI/V
QNGCc4vwhw9GM+rcJuOn7M2foovmXnlpVzLTHYOV6HFxYY6vCcEo1lfe1ElUt/YZ
oY+eOoDQwpK2EhGGZuXb7/nlulzPR4KPdW73fDJTu1ZZbCOmFUQYgyUiiEEPfCr1
SKcT6s1GnTtv9pxo9bQBBVb/JqkiOVIIpcl4URsNGdLTziv1VBPq8PhnPErHXE9J
gL5VPZLVCVKhyIDybVzwVbDq5d4rczc+nD4ODorX0B3KdipaW0tFuFGpc0DNn4/p
HzqL+p67Ckn+HqueucRjzCwpFIKRc+flS9Gx6MlBrVLBNMTaGWSIdzW69qcJt7Ph
Wy/lOC7tjiZx0NrDVedYUtEvNt29iVPRZLn9Wwr+L/A=
`protect END_PROTECTED
