`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7WkImvH4OA7ire+4RAlhgvwvmgVNc/sR326GOYNAvWD/3A91iOWbUifz6/n6jta3
+MbpajrxydA4EkEcwRpF4Dj51HgJ5nB7tvp81rkZ6LCuXGrIPLrwG8szW+3srK1F
ETVUSf9e0Yo30BMaEIWARUfwq2kf4gqs3zfKyyhR48V1GSYBEEb8gSgtWzE0XY1c
oAnJmsWBc3Xxa/IkFCMWQ9qm0t1YJ7fz0jYVsgUVTMgYRMHfNllwmM52FMkVCHMr
YXzwgxLKCxOUBNsgFn2mNfyrHL/a8vgKXR+p68CNaL+CoZITehLdlGXBNQTbCZm7
h3H2LpFpYVLfnRaWfFGGP6J5R5FagSTxBXqGTDssbvLeeTDXZth5IthB15Q2CbKP
KJNF+r9kaV33dF2BOHBxts1vAtZSPkDehet1gUG0WJHRSvkxPK+12nCW/LmvahMe
+dLQtXSz1PQBJ5LfdRK7rs5pPi4l7irHMLC+pNAfEyC2aqePi3x1Qsak2lJjd88Q
Ilh9mGGkwerUS7Y3cCKJemEpzamcBglvXa4u8Ns+OQTJn/fc8cDmvPb5pSD1fcHR
hlRl+YMP4CICKqrw+W833fCwq+OPll+WWpUNOwA5S32H7Q/5+IRkXnLfdqObQgtO
m2Dcz5P/v8+TYppuyr4qt5DYa3QlI3p4ReHWla2BSV301jQkr0r6DiAbu7yHFLmW
Z8Pn36c5o1r3m2Hir31HJwhfQFAgjIzcFLaFX5PQ1yZ3vtwmGlwR2nLKDIXtapoi
NNAO67xzQcnB+g4eVPcf4IHDQlKlFU958+tZyvTLtYOJrshmDIl8wZGkqwsml4xU
rQXMp52aS/rOfzJTKgZmfmub3AfKi3hOuS2WAdDUhF1YlIl8K8MbI69LvJ5OwTJH
KT5xkzRwBbNtsVLje0PIykVAWkOvFb8Lp/6m2In8oMyejh16AgsrK/uA7qMWbnAQ
T/98avfv9IvWVUp9pjmz+Fff7PcuLyPttWHg1osWxTHq5QBNMkSVFFGfAus8Y4TH
i1NZPfjmdIWP0m4hSyFx5CbK5GTaqpk2j2xUMlrhcQHJIVgPmmfvUkh0Uu3Y7vgf
9/WvxFpBl43xi64byQhEc5i0Lr2+vy/L74Lkn/JRQWAHWrL08FyLx9G+2fQyP3tt
prsTEORHq5eKz+LBHeO6gvgaEKaehTHshzV5nG+4PyQb5yLD/9sUptnSs1qVfgAz
/5ts23UMYIONJm/kne10dXcffyNTgJxiDOCGrT7aX8gqTvSCtB7ctznbKpk6atDK
83I+TyA6+Ht9JZiS4Obv/mxwHEJ3Q9ac2rcYns6DSKvY942Jk8vMjF49iXihdqeD
cTTnj/WYtbTrLlAGRjwS7+DSRRUurPXtE6adLLrxqKHG5CcRrlQjPSXvCvzVp+OX
DDX3ptiGggmfQXfaioKaGnjLRlRGHp5voCzmZoEzkiHDxNxn5zO555dGLIAh8Qxt
x1+mCcHOTpF+dfDg9gbQgnla+Gvgr/nFEpc0EaTVsxf5+GW8G5JPDd21EPCDdsu2
x91Yla2tv+tWd+Vba0UtQwZub9vVV0TlW0dZRQFxbCFVa2d85i4PhFCwHgBP2KlM
dmFlVg+bEvIfFUCCgr91NufZEsbIDzK0vk7v/q0dnpNLkHVlUq44ELwn7h26mjgH
Zgyxbu4MqQXmUU8aG/f47+Hk3o1eQWW1jpUZveWDMTUI2GrygQzNGt476HOpyaAz
a5N4Bq7YDLfBIcOq2Z3/CSyAQjO3LmzsFpsfwFEDAyYzM9ap3fDDLVppm1PdwnVn
4N01C+F9LDzlE+XCO+mjVh7f8HSorwYbI9llVajtY8kTcNyLo3SMkOQUw/DO+tv/
rowk1KSvlhhxHwXmfuho+VnSjvf7NYqrsIX7Av6Zqp2Il6CjhNMcx5p/d4Pqq5aB
2F4kL7p9lcQghs97aP8A9gsX1DxdBXEvGUST41xW06p5VrLKAMnkd+a6JxK7/2tP
jS6VxhjUF1tYH8dDI+jXkPKKH+jpfr7KPgHf7I4dAYLault/nAkr9ZxtTkuA0hGM
EzCDJM8jlRGeG0tfJDaZKIltBo10hMeKrOCc/b2TnzgrYcYoDpzQxsEB2eBz/2C6
hgGeO7/uKKPo0wGHhy+JDcc95HR0DHws4jmMLvdIdWdvjmsHwLFKULM8c0l6z6ZA
R0QKS66XZplT7micXZFiJ0KfT4NIeL9wBNORmCF0FmYqensgvrZnF5wmRZKz27ax
iCfX0Ng2XUw+PLxjUTJTFp1k0na4+Bl34smB8pDd7/3WweYWcugmm7UE6nOlgY2G
kp0xNUvCtpO+F6gfpVtY5QYFUj1nA5YymNwaMvTFob08mqEe/xjMciaHBu1uBcsu
S/54YUkMFsFU8k2SVDqN1d5uFuw+5EFhouGNk4wbtnFuEkTVHCWXM3RS+OxwOBxZ
4no6FITRDyBIcj5KVB3/6BRyeVvjRotKX8LyDkpaeUN3H/EcQ2iL/YNYkfgyDSpa
XdxEOc9sh7kMn58Rt0mF79X8/2mJehHG1tmaBip8hjGF8aj4SM0ptoBns83yr3W7
+1E3sz3+IzMhtq7UaIrNiASo9cJMd3iBt3aEh5j/7xB8MfEgLMeXIAYnksbTwOsF
K2xxY+WkwUk/W+t/nfAzMdy27nq2KqonUBMIfBvxxoLQfOpjYd/UBMYS+HVP7keG
9+KbW6G7uIJb6m+3L+tsK/Co+bMY9AtIYIraf5qIoqm9KkXhG0Hlnu9GQWP6t8lo
BbnL/VGzDEzhG31PRAS+noA/8jdAlNziVAEr6Du7VrZqLfUzgLW0y0fJKKLUNNxt
Y4A58ar56EpmBCfg75JBpYJb7SRj7rmJ3opfXh14T3MiQ4i+F+j47lTmPt6a1q+8
qoX9XW0yo59wT8t8PI3BRv9ee2wh5fplyLkU0zfN4qV9kWzUtHaU1BQudQnOrZMm
JUCwRAJB0+PCjmVBoEhw0lmXmjutwRyJso8ICElZThYeS+gsowIdMcX2IoNWCJ3V
Kgowq324c76W4JpWF3uqgf3Gr9B2DdNdWqPmYf8vEDSOoE31kAkz4rio3kFBSOSy
nJceoxayjPJCg4HYEwlKY+2CoQ7o4PuC2dBBRmra/KLunq69ijrua5ftW3IeLzkA
mCRCk0AMzkoeg5EK6R8s5BbUt5MpC7EkT3UjOM3A0FgyL4JnZwv7JhuAJY7EEqo9
pAJzuRn09n1eSwBaEXDOF0v77V9WBCxUSz2J617amP17nLVupPeO4VOKxmL4EdDE
tZYubTIDV7mQq08+vc5v8zVeESgOuB3p41mnElJr4sc5TmTJprJ4qmynaL2pAF4/
jTUj9mY4VGS4/uxER8tTvY8uXDPlUqyb0Ydnvp7cLyHwr7FuWaGJBEeszc7Y9/Ou
ybDpwh90RNqM0M2WCoLIqY3W1PBH/lYO2NTs/v46C92TvKZAXlUa5f6hBSmuDhtZ
idYpDDI6WtaufKZdAz8i+IDezuxlzrHNpZDpal9hHU2SP7p4MlqHgLSMRr2zGRi4
IcpTMUhhJXUfge55UlMM+gqotT+gUPBi7UhILv5gXVjjg3WYbtYaYNrxjrfMyf2M
R4QeF6yn1C7HfimG+/THOfHRnR/UzeYo+IeG/9D1RDbGoj2Pl69LJidyU39DbfRD
S3woJap1xpJcAU1/s0jM9rxLRPP9yEsTJc32U6oxXWj9LBtWv/a1n04DvE2ZrX0o
z3TLNfnPXQIpNt0mFT9BpT/Rju/Lq20oXWt/4uaNDnBs0kp2ePd84pOftogEXfiT
o2LhjHoxadI4k7uOmJXS13nemB3RBpBTeBUapA3GoUHwCALwL+Z2W4cC+yeaGEWo
LJJIJOI1KalsML1D5sGcTCfiwIYWqOcPTEgAGLA6UBX6kOOZa5UWSF//oTcHQjS0
5hF2Go8oxLZ9XAaQEUFYPnob4D/zSkuB8x0ajqfYjrOJvdSMA4FEKB3ApxTu/MAV
/Gb+G/gYA5BVGWwaTpmqqTxomS7j8By00ReHjrFweyzgFLGeqzhs7jBLUbB2uJHI
PdfsVhKlWbAguZwR0v//ipasK4mRNKB/K46RifzUnWqlNLAdsX4DjDn/qw0GcjzH
uzWdSZZRfqVnNOmXG/WPd6Qdgs9W0K9xGwyKu6OrKbt1wByrm4QQueegEA7nQCOX
QinPo6KoW2ScgM95sl+LFt4y6ne7pnGHuhAWve85VvZkFP0XBp/ezb093MymBckl
RK4RlVlFyZQbWm+S+jEZhTGZE2HztW5cV4tCqVYdn3c=
`protect END_PROTECTED
