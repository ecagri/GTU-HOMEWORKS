`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lJw9QbTWuhZNrLmtDL47RvvyCnw80N2KWcbjtk8OZEAux/juAZnbX4a7gzbcOqmz
pdBSFcoE9JIa22VyFsEPRCcdgXUV8C/4veX6bfPtS9NeovOAYn41Obet2I7iz7ih
ExmnIn4LtqAqXdqnScsds03mzIj8ZFv7Khy869mEhme3KoNLP6yUXJJuduXo2mKu
r+ebXL2dBHDVIUWMJ97ux2Lpmwf0tnTXEv1OedzmrWmdFLHpv79hQaPhsu6kDnlN
F9DsmTxRRyDFk96ctf4L7mXisfbU6TSdYzdQkSLYhRK90zn3GC1pOUiyrtsFDn88
wJE/YD+aEqAHvhFw6U6u6ofaCJPrfo51Hpqwi4UsGtycJ35kN5tCy27arrHv1gsz
WIZo1kZZq0LDt7lZdP9VupC6xAdRhBPY66PXx73IjFJUE2k18q4E9m9TkI7R7CPr
tBxs+NGOArVNgUOFIH5ewGE3wYY9jQj560RBwqFoA5ndzQASGASHEjvdbWodr/yV
UAOOXO0mus5eT8VFfh/5nhnhp2DAd2+L/ZlAoQZnD/NIIzH+nIAcFT045Otu7+F9
43X/tGyeDrPcBljG7lv9oQ4JBCAgghjzWJjW2Z9s827dVgO5GNn/05+DrQF60zeo
x9Pzsh57iGx/Gg7mV+p/Z4Ln1ocEjoQJnnPnHE5RdPKdt0E0x8zke56mpso10udX
xkKA7TsiN0vHpsfBSVhJNH9bNsjX7NliNaU1DZXMY1Holpyv2qmVhuGAEZoEe3kk
HJo+dOJC54fXZFROJIsNjBoD5SEupTmGLqNQWLFngLpEJBTN6x0EsqFOiRPJgqgv
MKQqVjF3ZeOR2CgHJ6SUfaMepLKHFm0/13wfle9C1WMtre4wJfIpI6qwIWq2yxed
Ax0t0OY0jkLPFaScEfpLyku52M4ERdNZATadiS+jgnYZeNanwYxsFNpOOOPWE+KR
5uqsm+1xUbNAugJqD6Jm0rTUyTBcJ1MC01RhiCmIK5UsXaq+37NaBQpnEhyWaJvU
VCdl3D2+2FSVgnjwbVxwx5O9YwFpChqpCmrc7qw9SMEus4kXHXVl2R8uzZEAfsQx
fB06Y2ebcUzBIaPxTZFMGjWGmYPgL5yhgDFwgFyvPgRk3jJHHpq5TDMw8ZoFiZcD
0m6lY6JZ1Fltd4qt4x9ogA6X1b4B4ZfoFQd6xYEgNZHiqvIhcRvw0KiITGS6e2Lz
JgxzwTjC0VHnB+opW7HIUOhkVq6qvSUShz7kc2PH2T6J7ciGjgB3AwlVxCKlg1VW
6qLY+dolmmfKBr4MkbBEOwteb5HVr4sNjYwrPXhdv7lz/fT69XUWjj4CrB218w+X
x6GPk7oUxwd+fbPJl4gC2oF5PlDKwi3NTDzDNQOC1SdAZMlwIUq8kx7skNm7WRxw
/fkAFQ/Yhx2aipPZrtKCG6L42vw0I85z9B7gVpcp0pHAEIv9GvDu+J/MLLSFJMUm
o7BvyibAPnpsHloA1qjy4LqeoaJKaK5HSnP9KX/qTZEqhLC69/4/0/S8DC36PZmh
wJ6OuQP9LkYMINvo5RESZ9riPUXrfEHTiP2PllZnp6FeNx7ztAqiJic/9ZMNqNSi
uBKpBSxzbkPvo/DQQT8RzlaaLN40miseqrV2YsuVYOYsnbp4qqCD+3qvb+ul9048
GnbAga4xepangnBFS5KMHpt0T4SuHGpcc+urqyojU+DFwNZ2B9hZHIY2I7nTA/aK
bOSQRufwLrjKS658K29wZ1/sJjAMTomPTQf4HsxUiwZT/ZJdMFOmhXbhTDeECNf4
+OUnx+q1IoSv9IiCHP6zMYodxI2mc86FhfFFSu9KHiRmYG0vjQ2aOBxZ86uCtARG
8VjnRTCr1ZtiLr3KQ8sEfNrBqt/lH1mlZCiSWLrwBw4MRuOj1NwAqLF/y4Gf3m/u
oYAF6CJqqiIAeHztYr9bv+JCpkm+cB3uHPDxf/gewCka15F4qbZALX3B0qnUzugr
oTrzbUlRsze6+qZZTh3bvXvBTrhfFeUblbey+BhskH9pQ21PEXqvBboNWZOB3HzN
8bQiAmyfDC1BG7RtUllDyqv19NVJ7Ij2XKI2tbdVO1bcY+daIHE+YGhShVSrN/X1
sEHaHHfyyccuxKVQ1NgVLomWDZoWFrKEzTl5GQu/butFF6wsHfa3xv9il0miqYk9
ZGsrKaODswDgwaOH2ll59jZqsTNVSCwJDxSHCEYeVHA2Tu3H/Nb2Zj8pUJHvPUZK
NNHleYdtNlu75NLX15DIWM6xDkqCmRj4lN9rKBljqIeffGg63JhjzuuumrtNrUu1
UAxnmm3+c8fB8cqTia5aJT+m5Mm9Fh7ro5a45vBgh2+NWMmPb61TdUedEpvzL9IZ
8rgg11fD1kZYQiQ5xDy+ShYXsG2xd9Px3CvbiUN3A2iE0cAcViXc+8eFnO43HkNL
Iu30w+x3rUWxq8sDiLKqdjcKCbx9mVjEGqy474b+WT6ejG8lO+8mURogi1j2eYLs
wCEiJf/+EzCHCCQYYABlv77nF+CXmKiGEbQfR5ExiNf8hqGAxaiH1avIpY32VLy7
LcT0BzLGO5guIoM0MyWaHG9ndOPfO2knpwpYpHug05TOjrrCdoWkyRVUKFfbUZ8w
f9a0c8K63863jQMAuCAcs+jJQKhFZd7v9uClKQ2ACz3K1AaaBT4U7+6T+HeTNXzB
8rDlGKNIhnpHbVdP+QiVk9/HmKw4NLOTiKq/w6ZyazZEdQjE/f1KTgpVedeLupmB
t96XO8gRlPwYzjfRBRJXv47fAIrdeLkllMzYX2lAuX5fLP6SPuQC4+UjnClHAHXp
JCWXBIAu4EWkXJsrrAAGq7HQ01o9/hxcSPqa4Tpqbc0q1MCESnrHwnJAYK1/Wvnr
OPjapTDUXCslX885wWdgohP2VgPjr2pi7lfCkO0X0NPcojIYV3KOaf8TghFS3i6U
izYc2V5nLXXajmWz8g6FV/fgqq78zcKZHeh45isvBsPoTLtIEntPkYvt/UcidV8C
SEXs24DWxdKam2PNY7pUn5i7NvTuYzQQEVbmI7XRn8JFJMClhWE0sJpwtK0bTp5h
FiJnB85ABsYSEMCOiOjrb7qIQ2Mcf4DA0p4p5CMdNB/xUb9bU1MTPef6jFskiY2e
10YBEQnJFrLy93uccdGbEkZa+a8m9G6U3dpPVQgpzsKfGcNywLf3qtAARAYAEUKb
6b0mxcerfCxutFkeVxMbm6Z/Lfq+/qEkSh8FPfunrUTcZDfzM26Z2697h/or32+Y
lvrm8iCHAPGiCKzMbboPakq5TwiTx4/m6B5XCvTHELPeQLbiIddwKPprkXOJDrel
TxZ7lYMQmNZD1FKmCsLa4lngszyPPEYGpYOqQ2APlRbgwzp0VBoH1YdNUGZ9w409
lyh4CFCLJuZJ5BSwC0HCDdUedElzVG5UqmMF0kOB6PpTd+tEUAzrue8BDhAJ9IT5
ZBvRBB0PdNwsP9CqMZQZqKiufAgyGh+8EafjFQMKX3GeQ7pfk2pAmkcalR+vvT0J
36FcHDRN2LDcwf0nqP5rHUvWPvfy6tKRxycwXnXXF+2L6/kEIZUnT2LcrvPay8W1
f6TOUG4gBsOVeTR8xvLowbLrBH+8/NRzc3SDNHgMq04dad38keCAXDdGDZkGmb59
cth4ll1lSgWDvGYu+BMo4dwEccAXZFZHPke3n802Rg8e+3iCzA4PtwucStJPIYeg
NDd+bWs4VC77EIovGAdEX2S6MuBveWFtOLmbRcMTueQQ7QLFvi+nmxBFg6L1Ri1J
X14a0ccuahdEcxDCAyA2Y8iUmUixhgmxYXg/fF7bqEa37bUyPb7UldGuDqqyjRpF
F7DMjCCJZO2RZeDXUgeVCoarB5ph2jMqx3p1SiZXvxpIdtDmA3+vK5ONXZH82nCv
07B+g/4xyv+A8ZdwKuggB66NXYF+ztiiwwFFz2oYtV9B8N0renNBf2QFw/Uj2dkF
xNC9s7ecN46H1NDAlCzDyV765IGbQRqT1inmNIIZJwszNDU31Hii+DpWz4JX3n/n
Je/lFK729LmP3AJ9vw/1+Df8gvXnhot6DQkaf+Rpc+KN+zk/go24afNjXUaIdlak
dDSuzY7zMbEUTifrh5WK3QQ9BzTazEMxSJYgwEr5SS0ILAGjjLlBvKtDsADXmrRL
ncn+5zd1221TdStf5pFcUIvu/M5LFoSeMPgq7TxRiIg2TsHup2lgF76uQYerW6mh
1tyMkFxqsIXgMNvNluegmu3zVB1PXrQ5yAp43GTGC01N0aq0TI2Rq7XR+NrIa6vE
UlNEYhEBp0vB5+MNJ8BsmOM7Rh9T6YoP+oKhPVl/AN3nCMjVqM3bATMAVkhBEyYc
de/Xkc8Clf2w/KItfny1VnHaaLzQMFt11iaL2jr5cyE=
`protect END_PROTECTED
