`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+gNbjF8gOyh0HovS9NA6a0vl8BwF0mnGYnhwBHo7qZXgE3a4Fhw0LL6Srgd+yV0G
kfI6IFYS0fbOxAzCwTGiI5/f/qux7qafZco+v6AdUdspRRVevH8dIwCNaxFflQBu
dA8qeMw4rHCUM3aJ4e0JnXj4uz6q7gCRIySPulQkM+T4g5EUxfRqWlnzuTIQ+nOM
Z2zrqnMysAY48NKYXVBNxI6pUK4JKHBl3G2DQfO9kYSLYSfobAget6F/X2Q51L/e
wAZPHoIEE21foX6OKzmTP9gzLTt8hwCaZ9p4fRx/6M4T3/eOgo+ds1Y9yip+hsIm
arqr26Pg4FAB3X4xeQDSNtLeKlBsiZbupB+sndy1It7gktW948sBCBo0TWtmgjFf
qJIv/aCGjoOBZqR5/BNu2ABZde//xLQcJjs7mXQqMJ8DoX3tblP+GqB+qplbts7V
q+aRzviJT2rPxgjzAgZv59s76DfvpNbw8LVB6lBAvd4xhoT11Hb9FDQgz81Iot5C
hEgxIGWTUVI5v4Sm1z+DEGUaWy2Fp7i0libOSdS4hgqdW1oeCtB/eoipQxa9ddLh
T59JK77/+S2Ps7ZVX/9qMpZykR+3+f/fs9DrIkfnHW3ASDEEqpgN9ONCNq68Qfs9
YHTyJhaSjioZ2A+rpLI3MA==
`protect END_PROTECTED
