`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ltM3LKZCr7v9Vh/LW9LmEr38rVm774HKJtkYK7qNzJ0CbJV5Q0RRrz/4av6/Fu2e
rRNDbwLE5F9DFDl5gZzuHhoD/xbbP0nASs5xn6GnWYjxA46bAxG++Gb+H22dg0AS
DLDdshrKSyWRK4hm/tinSY4tWqqT+p6N150DlVoEqfmbVuJs6WzRJoyUR8hXaV3b
Vpe/wvsKx1EfJK+77kod9ItyyXtKlmlCi5OXeGE9j/UZRFUD4ncj5l8ByVJa0vnx
QDDbubCc7V+R8Bva1MD0e6NFP9zDqzJ2xskeUqFsJOTXZXO9B5lVd2MK6nwpCy+q
3RzOPyn2qswDaV4xb8nN317mE43xd9VplDUqOTaK0l7KS557oX2albHYfFsWmGUD
MWRwbU5HQsOtYhuIgdNfvnIyMEvPoD+XqMv3g9ZWXIYiMda+Unp34cptIqn2NyJ0
Tk8w82nPxHXbel8ldihXAA==
`protect END_PROTECTED
