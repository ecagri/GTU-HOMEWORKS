`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iWcRe+0tdHZ5nWIxbzkNcK3xqDkmPpd9bGaSbRDvvZrau3aXgPscbqZUIVRonsIQ
REfCvfDOufTM3RmXD4qyZIy7VvJ88OvLMsQIhNOB5F+Z2NhnQQWF7Xs7BpLo9RHn
ipzvWwlARapFaZ798xM12sHWEd80RP5XLK3XzwDhKDRQl/LA7Mfe37+KH+I7IagL
3NbCtwpQLjedXaZTeoUEZAztoBk9VXWCR7WvyOFucmEZKNC7+8GCJlaQgrhb3L4t
1nWXg8vf46rmuPkEe/gw5IIbeQp5p8Oe6xe61Y2aPlHYxvNGHddmdufVkNYo0nqU
SiwnayRw/7feBD69RjiQwZVoor0l/Vh3jh/9mLyeByv9xdAgMPBDvPCiL42s44/g
/Pjm5k65RxXbUyxeMO7mFLiP+OwHjJX5G7vtPiiU6BURQ3yMIHafWrbMoneXKVFy
KT1F2kBifwXR9IPBDGZeu7Es8ToXPyCu/fD4oYWBUlWHb+QxVU+DKDbBZXKlZoGr
Bpzz0DlIxcwbWUiDCu7VIThmIyztZARRp0CgBwGcREjcecB48eFRFNV1yqWJbrlJ
H9ROhkbwoWWrMmOsC3u83HhdP4WQXLGznKlaxDowjb7d3j1pYT4ZQ72jgh3hZGGy
`protect END_PROTECTED
