`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pAnfTC3FS8WGnwTtG0hloU3oNgDE8RpkuH/pP8Z4wHaNtou+o9sRG+HkcE+rgjW9
3n8t3/M9C+C5NergsvfjAKPWZY1BA33IfaA6JcusjUcoB6zroj+A0RXnkEE3Ca90
CBlal6FLa0HKBJGgxNPkKDtSDNLzHbaH0TwXNRH20ls/+UDITaQ+JmkMWLzGshVf
Y3fqnLQKJFuUFF1iGQp3Tx/ptfFWoZl9kv7CtO6DmYcxODo3TWmFDx4Xnx0OTOPA
fmVVYs59KrJdf1c1ZmnhejYRW6l19Yh7C2PyqAPUvzRFp9bMWXgvgNOQA5b2o6PR
jK2WxrQz3TdXytDHR6h10ST1koaZJBziylmRdSPLpzIh/tnYU2kXfxIQS7NiqdfP
vq0u88PowkRV7Q1yLZa0l8ctKIHQkimm0WbZ3IrvkmVg2t2bs2bak8nqELqXHxg2
X9niPs8z+c7dbHtMf8ZJY8iuFOcLWrjX+bf5cMX3mSADe3qn9o3gSVZWBft3jNDX
0m6XTdjGnZbXx6ojIdp2KBnY2fPrVwT8w3+MM6To5zmTIhZzAYo6s/VzaL7bYDUU
najatOppA/gmKlDr09OiO1cUvjVa0eOsS/uRsIXk3yjpHWsdUgcc0cVYZMOJYqMJ
gt+QQdD6dsSFEGVVGjSC6UTtNeJ/ni/+yyPW+O7JzPrVrNa94HizQ6Kl4ufpbM+5
jh6M2Rhz+60nkO7vPomUye4ML+qVSHOjG3kI6Q9/OIeYf3qQ2I6JxaE6vWVIxqA4
3kbnti2DKSjNZrQJ/flqL+yalEsls6yb7Cergwh0piSUHvs6PI97FKz0QFLuwHdR
VIJ3mnHYIF26QGfCXTTRl6FkGngqN8SLTZQqu86yX6qgbUBfnXpMI8aXQ6V9g4Nb
0PinO/bTpVXbt6/KWA/xkQwXEGDlRuZZwRcD+6n+q/CMzNc7BaALEvSoaQeipJQt
ObYp+SCV6oy8awcxNZHMhXzG3Or52a7JasFeNIi8iwmAbHEV6RtmcmQfWxLHrDWm
bPx6YoOomixDiGji8+w0JKgG5LxcZ3JxhXaOnuUcxIiaeKCTjt83T/eRWfRe42qR
9rlP1MBvawxxXyKnIcADrVZ4bMXF5DSD1oSvuep99nW5esZyWA2FzL6gTQ6xVDJt
bdXplWA2Y0cNa/1e2KKm1+TL6b4bZ7D4kLCdB4t2JcuKnAGgQRz3qSqnqvTrVSy0
KPHMGKl36oKzxH5s6caw3aFf3JK6afDu0cWbDlr2/ug8C6DI28jhp1v7CYanNWOW
65t3IOgVLNiQSJIyuCk4mxhVCGHM/A8e46nwi9sPVzFWuFV4fS7uxbJNN6/j6TnN
RTj193H39ScWNcEtDQJg9teDJVTiiuGIWJ4InKo/XJAw0EU76NUV5hbyk5RQZ6Nt
xfTGwHrWGouTkEANhKaIFS3pTgjIFSsYPWb3i+7AAyM+7T8uNKAm+p+ZoFGuiIVn
IlbZyHpyZBYc7EListWV9UI4HAg2oJYW4holenr5+grUGPlkKbUu3D6+cIGxg4UJ
e0TIrQvVxHLuLM1s9+vSuX64pqb9kalvrJU9b62ipxnS8FqwpoqvaEghPNFtGQZR
V9X6zaTYQ3Q8c2QQoT/UWzw95mPfqMYCnRpv3Im1DhT8SlvO7t2pqGBgeex8xzDE
mNV5ZL0eRH4L8a5/d2hPWPbY2ZuU1VekW6zJNNLYfwNbCEqa6fiLlyEQmBk7JU7i
pQXK7zM6Q7bnn6lveol1z2S0MVmfRf+BXADGkiglKv3i+zZKv8w4P7oFASe/Qpyd
PwAbWeBX2PwnHBTI6m/RmqrR/Y7mxYfPVqO1kRkmNfXW6TE5oRH//pzHkr6RBRqI
NXS03jMUC3wUzeKCuLMvcj1HmDtUuE89uvs7CZO8XXBTJf2H1HU8PK5vDk/Nlp7h
R9/L/W67kMKX4ftVWjY072rQ4dy6nHqPnzKJfx0mIr/QUbs2YXwYxJat4ubfK+El
BJ0xKxUyBPHJ6W7CJ+2W/LMy8TewQA7H2cu0rsI/n0VjYBICR1jstY3N1WlnQr8q
vLLNh1xMWVBi1RtnspflhLso9NG1ALiuoDpOT3zKwmS6UYO0MziTa/KdrrDyuHfr
Yiobxeu6N56GeMXdIiWV3l7XoIXNdHdznWyHcovPjuh8OYXxsfzO1OqtGSZTCEGW
smROherAXwWFnfr3nSBUNtCjIrzg0E5pAfUPVvoRGxXZ45Gmt8LBBQ2akE2v6zky
/Ndv0suREIL6yY54BliRGkdz0AZnV86fSLBq+S6nkW6zJgzAhW9vCEtq10yAC48t
w+fuSS4pvdc4dnulfkaL0lQGJ66+ghClWRpBVDuRs4omFCxCnwuAO78yy+vVnDj/
P52yBgtyqZs6jlRHrSFf8EWIUa2Zp/vo8tHoC3nzaj3cthhkusaWPeyvYMgzIu8j
PfGuDOP/46K5OurK57t/YsVlXDqD7yL2aUxzKPUyGJ8pxQ3n3nRSa+XnGooZwMPA
f3++Pi/ofVb/kMROvLCYnEwrJdc/3VX8aEoxkkhvck2z9WuU8d4yHdAsbM+5Kjyo
qZlqnjbHxc2IQethjwPxZXheQDOZKPtBrmRnSPncxbJBm8cw4ssSUg7AIHJSDnEN
C9LjkVbMHiiUqw7gWGNquZO+P+JPr1Pthl3cx17XYtUGiMipMP2Bv7EVPgbRy9qv
CCIqwFVAAuOY+PC14gm/MNYnwytzGaGnb89rmgMeDoVje359HvkGrUkRgUXC1G06
xhK/oSfXjEzmjLKLeXHaNkWeS0YlEY8CWg4JrgW6m/V4ac1cg+5tY4olTnX/rEne
4WV86+1ZuoE0RvHhfwA636NQtRH80BYUClwP0juyhAsDQmdXbGsBd6uAFmZr2W5e
ExRx/7PyMRuXYxxn+0RsRt3TYDLEQkFrpKZt5uik88jBIrZqWlKQvC9uuifXwDp3
01rxJSZASBM7Pw8Sw9kCLCcl887l7rpmxi9+HR+7rA5ndxK0z+GMINXtw/t1QqeD
PggEydcb2H6o87df5QkvZVNE49pmGPHDLYnrSqRfCRe9hi9nJZmO4i9SWa4bikZ4
9S2lKXKjr8mut0knAOhaLTfnN33VSysoyrHc4lR0Vm2wKAW6YdLz1deIFU7OjmI8
gu5blUnBujUc1H8o5jX4nNNnVj1aXN7wyLrLT4sLZOB/zP2VufV4ckTcCSf+L3gM
vjM3m/Xy3qb9aXp4KWnj31ijto+hPqMVC76dgiDcceAKMZu8EQfD9SmWdgHJYIKP
Egu5d+LLFHDOk2H+8s13hdZXn+73j5upMZdN9GXofrYq1yF11WI0uERQlQXnZhdh
ffwgpXUYq/vSBHqfJrW2DVJ/3NSX7kOn9B5J87OxLMak0uIQ//sCqPvJW7sFZmn/
2DGsIYwzmy/EE6rH8rKxPYyQWh3KsZlzta6wsj6gLKIPRPuWb751Gg/5nnJ4r5hO
uXYbKs9pfawePvxc1KhbCX/GbF3WeSAY7gs7ZgsMe+S3hUATXJnNW6WzOpP49V+o
rrJOVylRZeTOTgn8DKestQziFrfIHdGf9+8MhNYhfOYHduyO93f13WBVfeWIeWyP
lmFsEZckyAzvQbFhYvHUUvRkp/GLDKtTgB44MClpl6dDh2XkU9XxU2N6UjTNJQhU
`protect END_PROTECTED
