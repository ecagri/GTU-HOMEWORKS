`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
660WjDgw/dE0MUsv6/BDp+mw2mfM/E6x007k/CNLnXZwLWJkFX/by4L8aHrYbsiK
D3TDTluqfo2smmZEvs8wJ3xhUn/nEdJF5SeYGcYtqaFXNLpl5TRyB3xdKyBaBiu2
Y28+YpD07X28plsTEsuX2j0xBwDmrH/3oT4DrkozuCy/mNxP5AWlR+o5z/j/HHwG
GKjo1KpeD/U/GT9tVcxwU9skhli1GQdITX4Dykbs+xAN4qfA+9cD8ocxH6Cok1EH
jhRP8ZGqOYPenRQfAgDwsnNJ4Xq3NZrHWl/crU0u1zG5I82c3oEW+EHekpd08Zu8
JFm9crKf7CJilLzdJ10Lmei0/2dIVPAPennFWy+KQe9iriKZWJg6aRCZHcauJAXu
taRok5G30uBRGIXkSgDFb34DjlnsCQ+stNaoenG8KFcJg7d94pAUspY2JkNxVTcV
k4oekhug7TX5RW2j1Cj8Z+8sVk1/ieLeOiyzNd4fUe/LHFXmlzZ4IME4j/Krrkhm
rBvb6Fm1VCcKCnUtYAqV45DI29vIxf5UKVapSn5buHeC4yPTmgdHq8w1/7xMq2Ad
AMQtQqP7U1vDu1xECc2pPqTxTcblJDvGMVTrBnwaYFw+Zu2F8yhBfdcLLaOQKEu/
NO344F6VDTCR6rI+zfYdw+fU2eBpUfD8ot7b8JJBIBl9YgXMQYUC4FZKGIxFoTbc
iSiijAwGF39MFUpb5KkA94U8PqsAFW2nPwaaoqr8dzVatPFwo7xxT0k20PL1M9cC
qUc9VcloqsCjGTmg/SffzldindeMVyxnIr0mFqA9QO3jcxCxPhlP+4zhRpUtG5M3
vXfFi19n9OVEFX1/d7YrrHh/Slza10SbP22UjV4jQfOWI+ilhmegMvvYgtiaVozU
szSQ3UJuAPML73SmNE1w93D83jYonYmU/VdSLl9aZLlEcFuD8+xcLPAULGa9Q12l
AaEZ+HsaVzF6jHaE3IlzkGzVmdSvUsDKTJhMrWU57nbXRv1KqUVndNJHcneHMyDV
ct9NetTE2diTOmOJrdJBcJxgJku3G1McFlNf0HkBx/anBCvCFpUXGmuFup3DS2ww
PLpBA1zNkeKBDoEzXfxUt3pwzYXllXOkNI7tNm+sAKyWFNJhjh9gzR8bbBZNP5pI
jrVaK9G+zYf1ToQHCoCFGFXrvbxnIv6OzRVgMXPMGHt0tY2tS+NtwquudGwt4qhK
zp7BnFTUY8QLm3RvroogqQ==
`protect END_PROTECTED
