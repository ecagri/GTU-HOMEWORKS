`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JXiZ1P6lzX4CDchdSW5E6l/fnQB6S2LddX+woI40+g1RcJpOL+jsI2jF74pH8//I
ECaQXPTS6vT+T192B0VBPX7cU1qjD5euA866VbvdeqHTgCPmkLIeYLI7QJ7TJEYF
/C6eYN/bZNLvp3bMBQ0DeWjBY1qfbO7vOE3xau//f8/4XO0prQAONYIm5hnc08FB
UYBmYKMZZFEtjlGLK64KKMnvBbyl7J3Z5B2OECGplJ5yRiWTAW4svKxDjnREcfGs
aHMa9trC4ItG6kPrbL05zKq7nPIh/pnQyMAWjF0R2ywc8dXS0oUREbDLexqEtsqP
CgSt4BErgq1ettWMmhz3rkihRc6rDpsp4YSN0Y4ZJGogTL9vfzXO6Q7KATAQ3tfK
yPA/Fq7weXx3m3L3+hmj23z6f1RmXJd/swZJYAAMRFwmSXXo/Sj9D2Bh7PQOrlOC
bituWDjh/2oSb8KzS46F7/R6ztXjW7UsnOFCaG/maL8AlRMB+N7drMbQ6wvLctYl
7K+1FO3iNqgOOrh2alvEUEyBrdUCzxrDjUj9aCxc0Kh1fNI2gLczStlqPAbaR5ph
Dxqh7P9ixtOUtYJlcTmk+UyMCj9zxSUbht9CBqW+w+g1BMYuscEeMzvxi4zQOBc4
`protect END_PROTECTED
