`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2JVTV8YKoqtTUIKsvXcQsCptOJEMcYYDUUn2/MXKJa05ZzC58JMZ7/x4xaGHqJlF
2n+1z5FvDdwcPO+xC0owH2AemqAq8hl7/jkLftsbNvgH5298YvSaJsoJ2spKt8vw
GE6Ivn1nDq3g5jhWzNH9SR2ubQvWe1uPw08cyL9uA4T1LNSZmOSWgJ8bDsgBcfyE
ebYahytpLFdue4Xuo2oSuVKBPGpjh07heFoIjKb2XHrU+LYXbnQWHROAMUepwEAO
+EMFoqxcNBAmsAKUgOo0NP4y1W61husgoGJ+0nHIxpMf/3zzLzsOD9Xnygi62d2X
NHoDRa6vG8qjnW2yUno+BPHeSgJF40nyFNp+IdERjKF1YRd5KqwwSd9nAw5iuAuc
xiUdFAvsKb4zKMEcQD7HQAzXgTaqe63v1W9Rwvpx7NPi0am3LaI6DCRLyMuv5L3q
Ra1a1XoP0lDkt+qRzZ5Q7ZTbzCjNXFZ67bI9Y91TU0W+IvmSKxlXtWDuhXZlgMPS
I/9p6s8j9IampxvycfI4fEhAFOijWmCVhdvph0e0ecOxzfdcElyFR28TWFFRcLer
ACAS0S5+b3/FNz2iuSEaTN+GrVOdtx3QKOQO+Sy6mXUKJGNZx2Tdu3w2G4Tl144k
hEMhVsbt/O6uHh/9WALCRi7J9djxqcv9LwPYen+F66mY52FdCO+wrd6Xyp7NEDfI
fhtgzbUK/AU3Ubr+58Mq//bwVAprQoZJz+Ul9sBtcNHbL0E6VZ5a6kO7JhKez9Lq
vXRDRLxvYayXvSKqc3dDRvw+DWzdNkjmNdUmxUuzHpQC/Cyc9obIX5FMqu30XiEW
DfhEMZOhNYxn9IhGkW90bBj90QvaMAbXK3BVD8Ksvjak+LGG2h1Zvlhg8I474XYu
gM5UcLilmwGaaLaFUGAhO5hD6WJCQObzzBooi0PWpHR9CHzTKZwzjKwSHFF2qeV3
h+51T/Ud0kUS2rdL2vzZkjiQ5UMEz6U4BWnt9JyybzBlSCVvvB5q1R6wZpqlsAsv
Z1UIYLCcxxkJuHn7cWBBjjHf6mvfE642tNqYlIsPY3usy+2OoPhWF2bZinH04eWC
VYpz6tEKpPiBTPYh9CY0iBbBMKU0t/uTJlDUFFpTO3esEgofG9m2x3T1HKqU24rv
VGN7yoAHRjP9GfQmW//j/P18NyfDK4QT9RMhkKlnNtv/P4JawQNSTGhDsgKgzQ51
kiQlbEipuowac11Bkd3nBGmwpFqKduZxJHGhjXEjhpMZyxPvIr2b7VJEPhjljTA5
Bu5QfiRl5FZXGG580v2ybS5evRTwXUaBIIwA+e2E6rdXg1pNnRFJJ52rGYaW4EFA
pZcr9ttdIEV8UGXxjD8Cw4fcKRgY3IuO4oeAuI3WJ5xkRwsmxuEWTyXpl51CUfxY
h1UjMRDDbn0HkS/51gDxLDLH2IAHjfwSe3L/uLkkLQ9IhaOFB/Wdam18kscRo3Ep
wAzOZ+Sk4Ecup2BWBc/V6OrwiN5Nl+TYVUChMBEbMF8GB+dNY49dBeDA6FXMGByf
/+wmqNebDWD/fMEVto/01aqzmt2M8Vm9BgB9hCL+YAmWBEaFq63qBYI3MQaLzuD5
8ADefTHj3aIyGwVvkAudx9CWTfwWBfVwkxMQDTcm2S5NPMoe1oRqFgIsjTCZiQ6T
8VpA4mD7Bu7Hz5aCLNMfCRTb9ek3U0krAOFeRI9tFC5+lf6Ahl2LOCB9mz71q+69
kXSh/tL5a4jQcTowOTAW8s5QyCSly1fgysQ7/VQfq+R7cVUphOLeNya4DOfhMLub
F928aqsF9XJESjcwpQTnl3ply8xF7iqcCNCAOgxqaxguYrrikOmRjXEsD8f3ZlPV
CnXy4ejrgA0MIee0hDu4x7WFaoYDWgfvWZCr6sOaKH7igdiXQVjbqyqpLbqiXUW8
AudPSbwl59wguYkf3mNv8JLN59Kd/RbyRjxTIZC3x5LEq7nMFyOFDtsjzIwYIagn
zrSV/1wuGQFP5pXjvk53CG6UcjSvT9mf32FqU96aXDbI4X+vhIcd2/MFZWyGy8CP
xacCqyR2gS5e6cB/a/Hk6+2OeUM2fD/k4Z0IvAKh5uomGoWFpw0d0KwMsn5lhXkP
tG4fN+7/EsUkZRJiwcQqIEPIj6dh88jOSJ5WgBgXlmeCpy+1fYFQW8iVHJlE2Z/y
d73yadZ0A0CSdmwyYUb53vQtjMiqHMy6oFhuNetW4A0cRIRPCCGtBoySeayddVrD
QvPRCe67btGaRGnAlnoE1ojkpGrDlDrPL9khgkvyZ39dVuUtQQsYX2sZ0p0T0csM
7WPN78ismsKzgF5eg2APP78blMy5FyxOi3pnexO3IBOxoUviBGZrKPL27lIbATDQ
wXT6bZOzBJMXuK9TBQJfXDK55cBrHouMC4GU/vQVnFZEh8NnRwqcsfzMPDji2/ax
RkPIijmMbhgov+yAkDw77TryXsUj31h71qRiTzfXEiB8azIsHRCAoNvy/wcJxrxp
UcVUQiCz6NjMfdA460wAJD5Sv6lHi/d4Xj/Ub2eu+WXOOO/57iZOQhr8nq37FWK6
QseJuND32dJ3JGe/2OdOnBYHVCdP51KfMm+xoYl9NTMpLC+7Rp/+1wQpLFAzYgvw
JzfbLQj0JiuwFRprAqPtV85QkdgyC2cbnd73mgFOggbyVsGQ13YDpHnwTea7L4PY
VMpdjG6OMLjOmbvDCvocqixY2h4E6aUeuopct9+OQRlNGMl++38xaCHH8JEr5wQy
WHvcNArdI4GduyvewIpQANKP+IYaBZ+HXBC4WcHsuWLm5uepl7uV4Mszp+3W2Dgu
V5rE6a8n+zAoP9elHQfcx/qA3ekNByKBHMhUyXiFTkd1b3FP3ykYmYmZrWUb5syy
Nuwc54M1zjP3D2qmhu4XkQS9RXVx/giMIgNoRUhhIbXw6SdGUUWBRV4RVMm6fay7
m3lZeNgOuBNNWoH5BbB3Uz2LufkWX8eRQXCSKxHjKfaJxa2qWcKO4KcV4Rv6BssG
QY10TJRlnPw3jVJ+GyO4mlObLMB2ZM1G4H3xrzPJJfodGSwFrJ0jgDN3PnIgsOea
3dec5h3EWZFiV1YvH0YmS8MFpuA/3oh48xLqdQib7Dd5WEgKTM4/lep4z44xvZ7H
IoxEtM+YqZ/S3ik6vNbqLIK3Csz0iHQwCCw+MfVl3AF/ZfEqzBiB/w2vZ4pbKl71
ezAcfM1JEP4MO+ozual7Zt+l6xa+Ng08XM5PYKjZECKNaD6iiij82gAxHTviyW6k
mNcrL8rlyH1sAFy2NMyjugpzqHv16+Yx/MHoczRfuit5FPO8vvLqOHrIy7eM1eK5
k0iBCWgFURHVzHB2tCME2LC3AKGySUQqsMkb08v/mvZhvH5AYYuiBdAo72h6cR6y
pGIfxEuOnZpCQfA9MCj4nPuKvXl85MmEnOCHujAEe/CURjflwAeckyg8iW1kiIxb
PwkqQftnHeH4xaRQF9Rf/f9SAgtci8IG1nepZtcU+lpQlM/rSNlwF+DXyW6cEPn2
VknFTm0DKrZlJ5YC46xHTTQEBrlqsEXMsB2TZNSDFqcKmkes1rjhd/G7JPCjyt4o
9U3Y/SeAOFY1PmVHGU82W1rRkDUBVzIO0Fkyeu93KNaeWWY9VJmiNVBjSdCIhEUw
c41RXXKit10d6gjDbAn3Wr+4T3RL6P9i53/WswY5zP5ydQ87LEVbqr4QrdkSnr8y
KZu0th9fVVg5GYjeQa1Q2I6ZjO3xNNJFAIq9mCckAQsD+xBLAnHUlacDjkK3WNgi
xcUezrGlPrzLxqm8DF3PhlPZgWi9J/fSV/hjSO1iOICUgD86ChwOeKWaNP9fvZkl
eN6Y+ycd3nMuiw5YVRi2BvyhvftcU06CiSRZxhglkjbbC8wPhdjnNfwsp9kiGp1s
fPuuUELSVBINMp1Rlb3x+hSHZiQ4atCQyL8L54aYB0j/Dqe8E0cTcDoHPqVgBiU/
+B3mZDHoh0lNcBa0sVsZt1DzdCg1cxLj+bQHgMPVdSHGY1POlrK0zaGmBdkngr/b
5tcEu/apL9BobLma5WJ3iqBWmsE9MJfyKZFsAFzbCQzktsrbq3hehg5iGLZX74G+
e42o0jvOstBzYx66Grx2LYwAFFufmgJxklUKeXAGHeWA4XUtx1OcL9Y9LoB9uU7G
ng2Dr+cIHVJuqpInuEK0oTFAZV+aireYOIYuFGW0NnGRM5OONm/0OGdu4qthoH1Z
5f+ArGklBgiVMLAlcTOmNvdw6ky8li1dFpme+dGEwVSJNw+0z8758AHB7N8nWHZP
B4lVHEYD0wnUk5IizL+jFplADz3t2jkoHieCBovx2K3eCw0oilHHEmh9R0A26hhJ
jpgviPQVDIC4/fMxWiT6Tg4ap9A+y3gT90+tfKgtywzXoNboRcrS4tYQk7jVkhJI
CeKiJNXnbk9af4TfkSVAubuRxGXXOledejT2UJLJOv/1wHMF6B36ramSlgTTNhf+
muHR+nCCLf+/DP1jiYunh3EUOj5ywJOij4k16TAdfpNvGF95LwK2YontRvSHorW3
70aez9UW5P1goYS/hy/COG8DJoyPYravpxY3o6pK6dJEzbUiTK2HfOmDp5iViG0m
E0SlyPskpJZgoRnDpCnN6qSCGqidcpIJNn292WUDejTo0m2FRtnuMTeyKkJzo+TL
1XYTHhKufPWICbXuPw5Nwim4/0ALvDB/Ci2tEs/B7UgAL5RpWwjVubnFPsKsHDhO
ZhkSBDTpNZhs419zEhIM0DUc3EMax+cArWC9xCn1UgF2Fj+qntK1elRkXvo46kCB
4oCpGDrVDABl1uDBBbqx9krq8HQimJmvQaE6FSbAgZgDg5vsqfE0bFbsjjvXy25j
yUk1bEGtNEVS+N9KD5Q4+W1gLN8SIPmwOvyYp6nl7eRa9FjUGd/YgkyGiktTDZPQ
yXxstYE/5AVZC2ebExQhWKUIrE5w22qsVxuSJvQ6lQFlhBf6hVX4ddQGq5VSA4WK
pz4YFwWQwgaY0SYqVP20lHn62fxqMgFJVEKCd6qy3XnCDVQfWj/bhqUHfpbxo2Mx
f65QhG2o11daIiY/0ZYAb9EWr0nZ/KQDBP+Cwyz3uZinthdoUoq7q55BPqnZzCbN
ZLJUPnkQZsa6GkxqYR4lAcKF8Qe/f0OVVfWFG2Afo8CRvCGYQVmJohhGrjK+VxuO
qkARxdtPA+A3iwvigjZ5tz1gfxjxZVHE+miVBZ1xlcN1oTt0ZZCd5wKLGMadKcup
3LFMpr7Guvcv+xy5Rc9tjlZ0pADxbBL4opAgO/x/lKvnPSOEcks2NYe5M3Gpvj1s
rMbADiQwt4tsTWU8/QipQNp0WLaKisa7xd6ryea2HjVm/UuRJUcZ0gea3bOp8MA8
ell64OvGk1i+fh2oR4OHtjXC2B4c2DhmsZ6Dp6V0Kp1/wEa+qxacJDbLz0gkFwSp
GN6jLrLWW4US3NdQahdHnPB3O9/6INLzaePJ+MJFvvatlYVxivMBeaIqa5tSRwfu
KKvUo+cXnWsv5gQTCxsOLQ4q91zqz+GH4o9MjzbfwGc8KxbUcjF/3erRJ7M4i2rH
JagNsn15I7QJ9C1kY6gSr8hbS6aaWsjcJR+vE+g2nRd+qzoksV0bmdm8txqmwfyx
wqxp2jcA/OnZSkxEXVKGVecXss++CTQ8YVd02hoO/3bJghHYzbyczyaMtjNK/emp
1bdxgoOj8VGJsRT6GY8i2i4fesneRiTQCxVe4kriBez8hUk3IcGIJGKukhcjntEU
C19RHsJwMudU43G4Abr127z9TAYl893RFbO49H7VJIIJnHBQFxhgfNihYaAororX
X12BfKr+Up1K1Ic+1KH5YUjh8mZsFDTPJtRxWqK3Dorp3SiEil9P1wRbBifPCk5z
TkETkUj7fXnkEQT/T0z/eaFokNGu2DrwBe7mJ0U5L6kbnag9DlO3+7CxMqhi3cS4
sxd2e+VeLngW1lhleHBVcbAxKkwVuafuKRVr+egOidgjmyTPKmk2+X8QLo7I3K/0
D9ibqb4urKbAJNA464+10BhUMz7E8YRbalgYMRGDLTalyn3xGLF67PGerbOgG+Zo
IHaGk/wRBfeFepcTCiXrrVrE8Xunb7306y5a7Nw5g2NCzulnW8FF5PZDq13EeMLe
zAq4QWc6f4tTMD1fmbM0+qtdKMoZC9dDcY9IJhRBqCkKT7fnaPXlbr6ZwOZt0pz8
MjU0LxmhrfTSYALWj+EhS7xtzKOf4ObU+M3n0EnrD+TAO3Jjor0q2JwHv+rSyTVr
b/v2W1oKwbiqdNocncMq5NZWtlq6EG1mcxITOchUBlUKq5y8kkWjQzNg0+Z4bfxI
YdCnQq3Folpga/UfeY8ihjwb+Sh+1vtthYUGrbEZAidxZWzmQYz96nXOL4UrexfE
QqvoigXLroZA4MhS4e/ZgqYik54+BNL7zhui9cF3u6cEIO9zrYYwfHbWfIGkO+F5
P2vo2yrBKoDTR779QYXd2DpFgp0Gy4lP/fiH8O2iBn3yl4C8jMlCVQKmPVLqYIHN
Bs/ARNVBTcj0T43lD+HkR4xyDyKSS2CgIs1FRf2Q1N+gUG1rnphPKNA+tpHTwgf6
eFIZG1/A83FLmj5DnPGH5M0tsByo+I3Isl6w4YzqZr7nR0YBR52qUeWorZMLnzcj
7DFXUVTUThmoEsHZln+Rz58BiUt8f+HAzVISkzFUzGhJx/WOpDJCRpuqjscy4KZE
88R5owQT3Sx0COEXAvCIQSYJVxUqc7ntC+HgNi5hU/NzX0zAzHR0d+jveD9wqL2G
Bruby52poRmSjE5S1ldExikLc2uvruI5elzrtYs2yvRlszEUxUWnaL/6OlP5ud9s
lPhLgJ2p2Oyo6lWAgw/vG0dfGDr0gq7K3By71iDRJhasyjBtih4Adt2HkV0CCpSY
5A/KOZ2jYs//OwLEnOi3k4ZetvJ2LY9yesFqDjKiRumtZbX1TBJGUeGW5wTISZbH
ScIHvRKonSkD944BAjHlb8PDCwH8lTiQuoNbqDyHikLGsid3HONDWf/O0GFbZqQh
KqkmF6OvFTAhiJRd6VH9ZAv6gWTR3YYUZJNrwS1upvHwm8neUOD0v3/tKLmw2Dxf
49yqlebLKaIhhf2gQdZLE6BKd3LkHuIS/IIQcP5s0i9bekhGL60PxRnvoqRR+q7c
jdVsudcm5VdTfz9BcuXmaFwZaiM8qBhXyFwpPHF6puAPiferSv/2Sj43R5F+spMZ
QaMi3eG+Eoe9oOLEu7ja4CwbMyjJxzQkjxt27AR9oR7C3pimUiQ2db6XKQUDPqyt
e1lNXrxFMBU4SkpmbY4lbXkMn5tW231TX+q0+zVKYZWPguMWDMDro9suRTrs1TU9
j4c8rxIvGkI4HlvJBTPgW+xlxQSMWv4aLixtkOMjgsa6igvWvyhVx7DfNtyeWcWe
QRM3k3bOhKTQhIQlx/qIdhxqvXwyHsE2hP6uBQDjFMm57Ewi0dVv4Sl6Uqph2pQy
lP/YQ1LSOkqYzznjkPvgH2WFf/lbZ/RDmr8dTsZlqSvabKbRh1df2227IjhMSkr6
2sEPffdIo40FxIVXdijgx/RBAaMVpPyyyTsdSdQgiUrqmN+T7ONaWbv8AD2k6ZG/
4BvWl01ncNhvwGvOrFETMykYTxcd67Ca2nHrnTJn7SNF6IB2lfnHifjMpe1GgT1c
jTNx82cX0QnaH66hZg7bNCk6qgrrQRAuX/DwQcFdHOfbJ9xnAEToyAFB2rfuH/cn
p/1wokcXWOHpqqi5jIL5mMnqLCyz+1orDwZVmXstK5N0MYxbqDLZ20Rna3QaWmyS
3mbfQON75o9TN1JwzvQLSyRpi51xIXTpLQb5ZCov0CMhww8R7/+B0DqBxB3jJJyU
ProuhgkNPUW92uPVN1yzOl2muEYzeBwpeGaSYJel35J8DKIGyurbOw31RR3q6GWY
GjAVMT+1vtlOOO/uQQpa7fkOod4jpg58xMK81X0Amj2HSehUjYByQAjlZqudKgEa
rxi5neLOP8WaHo/G04FAT+q6fIjhBKMqiIxQtcKSWsYUt1jpnLhIH2pBI62Me1FI
4ciF6eZ1+aqxsPu1yrix3GFHJE5tKr7q5b1aWUQL0mP44Yk2sVoHZWbh/CalqSrh
5Fd52+mNsq73DrtU8NXacz4s8YZhk1dSd3wDPFO7ymO2FcMDpa0DMMfdCzctS+nO
ZVw6ViiTI5sxao67rAQSnDUN81JEIWvVGP7/MwumakhTLJQ9FT+IfNOf6JOmbWgs
m3tsrAn+7no9NmALFXQxjPHvM1zkR9RM10BBXoTbVnkgKqddBtqotqciTsXZQxoI
HYnWyV2VcMEurl6XpygSAPUyY+G/Y/QdJWQR5CAetSOZpCnQf6g5cL5niEddrT45
QslMuMUL4Tbq4QU3oA25goT565JMPRAhzAki0oeRottmK2ELi5pmcgTJjvSx8hGv
Fl7t6bZkTA5D089cwFn4UaMXzbbkng59EU6UiFixe7AHn9Ggf7sWmCg9Ca8RxtuL
MjcPOKC6/6g1MEmthvZbxaVgiCHc2LXSgH0Q/ELQBB3+knxYy1lT/UJEpSUpHr6B
+uq1il+LSdtFaBaGB0ssGBzUl8im2jgDLHK5jAzmq+Rj8fNTdOiIcSup3wGEixiL
AwBA5v+rHMmNoDD+6FRklMGI7XIeQCwclJU0M3l0ZQgYKC11ax2eIITkez0HIRO+
MwHE1vMnJIXMPYHR3zDMUX+V0Zf+zT/cYAederuaARBwpakI9TM3ysW+y1IMSb0B
9Scpo70QB1XC/i1wLULgQ7dvNPLX3lzn+1NaVNUyJUbmHhu8S9byoG/sC3T2AL/2
/cMVuCFocFh6gNJrtk3MdNlD4P8BJ0Jl9O5W/OyyhQinrkjudJxps3MK6OoAy0bW
puzuKQ318jRrH/7UBVISrNqx8S3Y7dEVCvlaboiyQNiLBjqV2T7ons6A7CKdtrAZ
bYj1qpI9s2M1V+TC4imRzGSFgadND0VVGqJDdt9eTEKQLxCRdDSbbk7EGGowBQw7
Tlhl18PixUOGf21p6iUhLDXLqBsYi8fEPty53j49MQpOBi5TTex/LAIFmCSFAD9u
QePQ53bqORlHUKFvQyZIn39C91n4blM3vNp3DFVFVXc+1nCXcC987hPLd6bq33Qb
pSmWXhp1Iz2RsOVJjDYbuWR1ou2biIAjt6ZmuG6uOTPVtOFiKSr9ogitcvaOmvCb
uneuo0/BKNbq2OOoTXhZFW0hDXoHEAfnWBVv+2TF9tZiYUqzheVDTQ2dMwmunlSG
e0OrkymnbHRF82tkQfk8CcFwpb1pmky8h/zmYQL8Y9vxw5YQ1jMPq6NduWKwTeYK
ZBLuabqKcs1SvcV18DFooXghWdPX2ydrs57l5MOC47dxabeskrzl8eMBDxX8LK7P
pYFeNdI10N4aH8z4OQAIRwqbrGSz30yB2pnsK/5zw2NG/gYh1IRmiA0U/+IGrkPO
2QiSNwf10xaYkKismNenRvcu2LnqfcMyZOhFV5ioOUQoG7lzct6cCyI/zlDNV+Z7
ZZLBXXGSUAAE9s+dL3846crecQ/jUbEwM9avSDj6Zd58B88/Qj2KKndgANJQrcvC
qr+t1Mn8gWPttBc6AeD4qSlUqj8zq6+MvdrkuLNT7kGXDKqkPwbrBx/x3GGLyLGg
8c8ttlyHwnHG9yKDnaYTKp9fT6Ro0fmmLgySc02Q7IxJTz7on1XY09MkwjezGOck
9scK6yrs/7MPkoY/gJbYdHk8NVYo4JMogquBTGeGqiPewTKpQbaC0xig+nvgFpDl
dtf3a46QbqVhXuuPE6998+2t2HBP5Pw7a4XxSNW0eceO5ck5vMo1wpxcovRs32zC
ETQ1UTaAGKZlHRuDocpQAbbQEC5EKB271YAew1jmOMYwm8muws9/YXItiYCpMob5
Fpv+Wt1sWfM6a608DeWJVYMYFb7Z8673n83V+qlkWvzdxr4ZpJjV1ZkYirnAuYXs
5ldgMc/KdZpUV11luGSv4VnFybhX4G56isCHmPRbG3W6g1X975OoPFHl1MF4QVzz
GyvJigfw5uCe47nccFZjq5TAAmrefvrXTx625wQ3HroEVan1nemKYp0/rN32ENjU
ncqBtEZAg7swZQ3mOjDaDTsFujZkhOoknJ/xEdb4AIwTfdIAa3uXUsrG9d3EGuxE
mTZdmMlezo2S9mn1sBIPAtw/qIM2Roy1GFRVIIS8+zFo7/IE8saG2dQr7fiOuNEs
DjF8n2gtK3BTXTdm9fnhkmuepgxfFVm8se4j6rdkg+q2uwglc5Q5DQa+2dNE612I
d8f1mlS3Wxb1AwusJfA3ZloCFJAF3/o4TuPlMMANuTNfqjlv3ZKXy3k+C7QSIvH0
8bqlG6cQFYvi0BCWMOwW5veHCuaFwNqC/dA4i9rvsAY6i51br/Ypcfte9d6EJMNi
NPQhkEeBzxynN2t1Nie7OeQ3UnCXDLzFOlfD/CPgEFUJK+U/pzMepjlz5MiC1vRj
vrN/RplDp0FyPcA1Kp70Ut1z4MWUfeGS7F3HMM8fLd+SY7i9S/c8015rwpCctTn8
TAGkRvuzjjhpbQ7uT1gQeShFShwxeIalPBPjyJX+b1ov6KsNeCOsXKRmp94S3BTF
P7OOti97uATPjIj16Rj0fyfdNevTM5ng1+tOjlaACdzBpi3j9OMJQ4+mI9XXQ75u
Bqk/ML7ceqxIZCtzQ+FSJg==
`protect END_PROTECTED
