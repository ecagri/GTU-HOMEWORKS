`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xvRGdl5d3V5oq1J89MzWjBji+zjmZwoKJ7kcPMelaEm38+4OnGLona+5xj10uVsI
IP2V259roPOZyD9zsUMHQxdnhzGbrBUNCogEjH/6JN0dWwARYpdJYwn7unErD6JA
jCJX7v6RaOOcxrcIPKNw5MUhmIPjcXVgwJgRSe2WHEZy+XZXJ+gpBHr+cdG/+GWs
Xrzz3SANYDdyL4BL+NZqS6EfouORrsC4E0eQeUAal9SKldIgfxG08agZg1Kpih24
TJgim6ZGvWSnhdv5D8i1L7NaCQi/CRO4H7AcRRvAJY5mQh6nwB0BWv4EBm436cxm
tcda8risB10mdlHQjzmcvstnHvBDPaFBek2KmjfEDEs0qUlnGq3Au/hZ9pZpzNUO
6WMGV+nBsUMTt0+RiDPTUUzAL8KlL2zn5qqZcqb9tpBKunVdrfI4kp7tnlGtU2Cp
dDa802zo0Mz5OLydqsJnKoY2P1LSNMKDojWwu2kM0gE=
`protect END_PROTECTED
