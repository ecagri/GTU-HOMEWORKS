`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ga3IHiWDO58JWtJhsgNn7iWpJCVTmeswKGOkxNdwzqAMlXbJZbLXCfTQ8k3X7jVC
HMdNrLiCArRHoPDcH13PvutBAHRlYLk29PSb/9RNHB6kuEWuYHGpGYae6oeUoOsL
egiY7MAyA45nFC6oa1KyoVbq9nqpGdzW6+LZ8DxMFvBkdyorOb48PUG9pH9l0MzI
ErfBZsBpFZ7LAaNhEzWM1TGUAU/704mbLqfwX3wTgt7KJVXMUA8qml/2VeVNkiaI
lwngIHGKQ8173xWwaQqhkY2wAri38hLD60mhyJO4IdW2gni7bS4j2bsmTMX/5Ues
tgw1RyrPq6B6ulWnR1AFw82GXvM8YeZNqsr3BYYwM4lZOVMOhRaimjTmoczfsvlC
vJGCKN2qCRhblYnqf/0jfL6MV7ybvyR9GELTQl2OpXShvv6dfdNBicBS7vTy72DA
bW011JIhOuSEHByVEmsIgFbzrN4kpO+D8MzRmONLnAlM3A91gMAEjIXvNpJe995O
4Y6dlcwhXBeWVDvn60jAJ6+p+dxy9Oukkq0i1QePv6vhiMLM05eIGlJlUEjX5inM
eitaj9cBQM+OKk8xWYg+dPIOtkslLJw3XgeF5tUESUcQAG1YxxNRdQrkYT8fxpNS
PCT81tDp0JwYWZwNyqvcUA==
`protect END_PROTECTED
