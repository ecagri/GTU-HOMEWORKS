`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A6e9ZXyuwNlIu0dM4LNHtDdeJkTmuu5YK6i19EguZyHMmyC17I6YVdn+Ep2bcBfA
XfHi7jJsjvs9YPma3n3GxRGzTDwT+m0LcJaecTElNJjZZ5ngMUIQSJCp6PD7wPbA
RE5d9xlH7928jsGgFurtA5paUQEHuYquUTRtQPiePvrJjx0fpOMNGnrtcqW0h8jc
BW0JJhPYMpH+W1X+xVM/T3nkgsDE7O6MPGxCmNXyjdjOzbhyA3EXF5lCaSjue/zm
VwBL1QJM6aDCxUVNafNhIiOROIJOULIvrShmLWl+C69Ru6YAPRwjr9KtuclKT1ao
srEnfqYUYAj8fb7haAM3vncgozyiZvdKoyuj08/s7ToDogH4am2qQ96qrWAE2roy
WmT7RsP3C4z3YVnI8iFbnNHckZ/M6kuJ5PHGoSNjobnjmpDa1wQLjEoS+eAOLd9z
pmMMk0RljQjADmjXv+6aEx22UDfEx7ZfyaNyjKfK2RzQ7YzwN6tnbLdwHtk/KkSu
NcWChya96ZNVcT8kLgCZKzFHmwsZBMlmRMcqoEpvrfOQzMC+bCKdGoLhXk8a5brW
n/4gFjJUVLwbDGjyFtuhWeg0+//foWhSwMdX1YWT23oUdhZJ/GWmEb2NqDPcoQ1k
/aoNCLcKaj+DoQYhLMdOGbn8xNFT6u2YeswfKsEZ5qw1O0dExD10AvcWuYBP9Prp
dLIwWYfZyF/+MCOtwa9QyLkqhniRN4b/g0fPLuLlDYeOoiWQEgaAF80xKeVpk8eF
qLwaGkvFlYLzlF84wmTqxCm7DpmqJXtiyny6GPk4409Mw2GNA+ejJOPW6E2kNXcw
`protect END_PROTECTED
