`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0gmA1BYOIGTzV+kPWKMjVwi/o1UAXBI9j37soUbe92F7nRr2NEaLbdfWBr5Rg76S
4RVGnJ0xy9x09/HiF2Wu20+IbpMojKI1CqNlmo0bSFEpLUwpf9LdLHvRShMwz3oi
rLUYiHB5dtfUGueuTKjx39BGm/sKhuazO2rgUd2HytOuy/ZzBTKkg8aILb9P/uMg
3bRO46dkcblY1U1UuO+ZXm3Vq8H2zFntrsq3QJ5FGgoBQ9+VJ+dm/j7nvT6c4xwG
R8pcbP/CkZV7vz2sbbQ0B4NrW8UDfgHE8Hlp4K8x/jfkAy3vC89lgMztBgz8UbxT
x7a+UlszFnhgdgdIFylbBiCVLH8agIH5fOk1+2DxeHqitqi/mocq9jP3Y9UiX+gU
dwEQ1dy0WEHhxTbeHv03QAnD6Hn0WuAVvw0VN0DSibE1EfhwIDoIvE8OFdoZ4cll
B59FdcoNo9BIBFCt7fWuLqU0hf8RGV+xoURFtJOoSvSquFWRK1VnaPm6D4FbG9Wy
NuAvNEChqRYMsCq1xuiP+njJyJ2fQwlNXYnmWBy9QYXropCOLKFh9083JdLk8Ihf
i8zTDmBEXCmWXrUKkcY2S0PkTzXL8EJgCoRyI2tI73HdauG0/TBZ7uJMkaB76oSY
h21q4gt4pYeI3TKgUjxYSiJgoqZS+eVhp66zgbE0IrY2qlSwsyzINisk15Q6WGhq
z23GVyD2eBw7yHN9BiqyFXD7AqL6n+dbRlpR7TWmxmbb2ovjbYmc13oBuYP2uAqm
bXUpzV4fCeSL2cLb/AAL6Kjk3VWUkafhfrtp4Af4EiIwjVUQtuWuU9SuNVRSpeKI
BY9jyzMGZLgcslLOld7aF8OHBTbRwQzbg7BvgX/dMIhAJIsRy7iMBfujLFmzKT0O
/x4qcRoGEzs4NXnEecOhjY6EGbyIYs7HL9KM6+01X53sbUchl3n/SnT0MsaBs9u4
M9LkJhubgA5D/ZSnkSX05zodwec3+wusl+jgdrVE2j55kPwg4my8seoVqSYCSVin
UvPRI1Su8AQz5jvrSzz2T+Zxq05FanhtNOIfszYkwGCU75Oy8HtPLZOC9bdIDsQf
77DXZHFu+EyryySvRxVy0gEGBCb8qsrK9c9PlRjN4bqLlG2N6VAlapdPLyNeiz2w
nkMlJOOD678joeedvIYZ5yNNHG5XgeBaoZDtSWYrE0FnApyufdDuapEVpXAeDdXG
AM1X6zm3xzvihPzPv+Qo/oWW/OOICPlxTBARXpWt7TtyTYNLsaCY8QrJk2KSZGKE
WNi1oaYNPX/ZiWh22T2KU5iF/M5dZxLx1q5CDrc5EBIXcbXX4n6I6n1lr9UajCEP
6aygm/Kipx0UCKmFEQYYpaduotDAAdzJZnc5ima6OtDI/DcKI3xfcK2XsuvFyYdi
fwk/xFvtuAcc1dsTljtEs5862Clc7bTUMh9BLEvXYIxkY3OJ5cMCh33LCxka5npR
mWDpCK0vvCjqud06cGSx90CAjbExfvzPWttGjz/lrrfEYyf5qJ54moRp+8LzSghE
v1GBmsLuODmbCaChhvuIXHMZ446X7851ISbQvFwwFedRwrh5x06lkIjny4YWBppo
d12WmC8lyTxiV1UcnQw8Y3ZjHeCER4WsaoQTYJIwqzvy/p0j1g/tcU/Ul0LfQ+ME
r6hu2FFSOe/Q5CUTPBq8bY/jjswvaGOLRLKNJDpLAIVz+WmbIOkaoJ4bdv+A+Qzo
ZRdY/AN4KOJdN1olFdM0pfTXRU9+IR1uJRsIZVdkp94IQ5A4O7j6sTUgbYhH4URO
v8SDt29rAASbt486zR3aqB7s1K3H3hdNIIHP324iYrHn1gm5iHKLIGBxrYZpTnsD
M5pbr8v6/LlS5ymozmarRx3bMRt3wDdk/HQxcjInwuHCM5uCEw339a6EAjnjvNv2
OgcUnbKjRpKk9wBL/zmoWuRSPAZIwQuvf9pkujXRkNp51Qgujcn7k+ljaYoOD2Ah
dwBRl8Hi1Ve00liN60iFPxSskD1IxhyaclZ4Z/Tp90Q8r423TBxSzkj7E1Agv7gG
B0wO0OQZJJyotHrlIJ68IWcuYPDTQhA0BRQ3jImvjLfBLZLjvnzGIdkQLtScqJvY
L8SVvgVXUC7yX4cBk+dKyutA1NqP/1BQVspUohu/zgP5iZ5LXOILsRTBDEsGUV30
w4+AtwperxvJ4GiueP1w8XJDV6YtgtzspzRebpJBFCAcUgA590rRmQssYZUWVCCL
Z8/OLJLvnXVYxw9Wu3DoQNiH3MDWXb3tXbcIrlYdrypSOTYQhwa/tkSg0uswIhDO
Oh2rlJorxSv6dykk1SDKC+SGRWBGd1A+Vr+J0RdoyO7mbjDkgTnpVoJ9P61lkdnc
OdgHTOrND7nlsc3CQNOO9QFEcVqcF5dteD/dVkxC3eU1ORofokqDgJdIuZE8RXju
/IjKywTTY1NWe3zlSjJ7uy367/O8GHuWATnWtcrCmaAjsZGW883TvRnqumvOY8vi
jbNqtsSq4glEEOJNQT7stA==
`protect END_PROTECTED
