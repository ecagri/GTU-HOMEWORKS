`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WwDMVUgLXfGUVblMMf9cQa5oF79NN12INNcjYjZrcV/YEOAyX06I5ggl+fpsaEao
EiKKpUsVcyBZG+L1lMyEAfNkdadrCNatZVuBgZZouuWhDIQMiV28nMdO76Lmt7Fn
LcIkzZ/aG2KA+BnZIwAuYrTr71ArNqP+gg1YVLFRbuhLdmvsLEEXhgo2bMteBfWX
kyCx8z1lTRqAapxcBkyXzQdGDYsiGUY4siI9yYj5dUCS0xcW45qjNp44ms6ifhk4
CTvaK3XT6p/dKaViFrcNyApGLRGl0d1+6vilU55DUjaz/ry/HoO/YSOuw6JLm42j
2ipQyNyJEfbvB8tDxplUtHOXMp5gPQKRBuJr9wW3LKAILymhUNEhVid2WZnrM9cg
0x8ZMuNnBQyXnCJz0XYSpaZSFfUroFScoFkUsXyUUmngcUXHZs7/ylZm8wEXjGCd
70qHDg9nsrGJESheQNcQJzcZwOrwwcjE5qgN+cAM0vUeCS9HGqRUCsCgHkas2i6A
6dGy5MWJYbAK4xzdDupS7JSbsQktupK3xCowQaxVkaZBHjDCVrcsZ+0zA0exhsch
K2Na25k6lUdtdJhOayS8fiV4FutoYJcSypv0v3uFvEJNcXZGXyRfw4H42ioRsZbE
/hMM3nwi6/lgDo1cq4jyQ0CB2rY0gzHatJqCh7fkYUu4DlYHbNL0WQf3UWeirc4w
NSf+Jd77uz3Rojfdsf5bSqaMpK8pfwMgoECpFZbFCIa/q+Ui/CQY+jCY3+sc0vFD
gB9E+dcTlJwg66x4TCCCBLQCZ7c0zWLRm9U7HMxkkRbC2D5MTLM0nIH+1vz/QUL7
b4sloEvLtoFEPJuR0D3E3bQaAhyrGkD55DAY8/K6/exV5DhuZY4EKFeY8fKsoqq0
uN3oklTcQfBEMFhS44rjVpn2L+pV+Ae6AdkIYhgsklyVvlsr98G01KvaIXnnhS3c
k/Zi8wjjoWatdWKiRAsXJjPPgKWvvvOxi5nGIFi5nqCGKckOacVEUG3lJFwZaYFN
puie6Mmq1OF9YN0AwqHNQqWip1p1/97xGPmA0IyJbsp0x2hxVr7KdVPDkopT06Yz
bM2s3Jn4v8o1AWS6cxITpE13HCe6RCXwJVY6+ZyBrnfd5n5GWRXLYAfCayH479hr
LJCzAxRkp3e7ZMIFEcXN1MGziHfAxkebaqzo49ShpiHsNJI2KCuf24PT0IMtIHX5
NMef+GepK+JjEZrIKsocNeiLlFIODVtygT48iwB4qL+YFIb7sReH6S2NPsPgFLyg
YmVPwdD9Qq4eeiz9EDDb8R6yDPUunNh7tCzJiNc6SccVjc85h4z9R4kYLv62buvO
w3StYLWc/3w2nZsFgnI1xyjkKQo6O1MDCt8z+MAc6vwCEgFNzdtYabu0Wg1g6NJ9
dajoSVCDxEx8DboTNOkpe1dBJP8lnEvJfim81dDtHFIIDA0iOjD6RKLV6N0MAjzy
0rvsSPUpd/MTukcvtjg+U1Cjg/N3AWJMfRniM2bTm8WtQ0GI3+GlxhQIesi+ywYR
mLRncY2No/3NqdZwVkJ3doGIybskDpaFOX0h1Bz0oce4MnAvFO/nzqK+ZkHvLPjt
KieUnybZGgftYlzSTNnOmRVB/IdE/8oxcYfONmPRYI7XLbwdGrFQCtkSqKX7bbiR
`protect END_PROTECTED
