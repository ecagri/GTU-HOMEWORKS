`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/JMWF76fb52m9mdB0H/lUYk8FkZvHQ3H2F1lXk2yKsR+GXm4zLvsOMAXdQOIpG37
b5HvPUjua5YOakiA4VWjVu+gu1tRnyV8Nw6NnomcqCA842Led0gjNOodeocnmG+b
u5rGFGjO12PsrRCy9U+iCpUJp9brOv62zBDbg7xFY8gD1PlAvxGd69YOpvQ+7UbC
nGwZ21WTc+NVw5lQwvMg5i6QxUVASHBj+JOCP5+aaTk5COb/LbS0QVVXdF5KJJM0
cc7OX80p1ve3cemJzD25XMNqDFBWugBslLJH/E37r6k0KjTVFpJnuUUrtSL4aWA0
V7DhMkHABkbmu/zs/zhr9GnGIhNFjhTWHAN1VdhOLnt/bgvEwIoyShz00f4mZncU
6ObMVuZvrScjbJOBnz2aoQymtTYRyijW3oL8vYhCAUOMWCPFk4dNjmlUvZHMyUBV
TuDWV/trK2kJbZJ91rAo3+dgiYylc1dGnC5G632Q1jKfTimbuD+3pcxaVSs8p5mu
N5/Q9uUUm6P/IizYec1VnHng/3cwtSFYb5gt3mMGXrvXX7VtEfk7AUvdc0uh+q73
sdLQO99MUC5hcJUPuIxNMqq0mKiDJ4yw8YYlYnPXzE773kbPXDuQGKOv9XvBzSnm
WqqDf8iwowCZbJIb0z+ESYn8H8n3Y1A8tl8wOK5ndboqhcI0px4v+W7zTO8obFu/
tJBRGnD6QN87ETVL2oryEX7HswS9KJBUrJo9sCcJlrEcp4dKvZ6kTcpr2FF4Tase
KOukuhveZP5txrQ6qlNRO1UfNsyvJRTOc55OLgGy1yCtiItzJa58+pv70idKGjM2
jUs1tVl4GgTLcOviNIqRL8gDAXK1rqUuoxlt80lhXXqraB6ZJEJblKDEhCcagn/B
AJHAW70EBrL/9h+QLRLaZ+OGI1l8uGWtv2exsYIXbe6CF/3XfxkZp/zoCdjr/FIL
3lv6W/PgGNt0kUqMwpmAjzTDdAqjODwGLNjW5U0E5+VEwIQsMX9kIu2yk1MDFSQP
EUnOHhnUavAj9qtHCNzYFKuMPsGejPqiPenar4qsoCls58si8BtOex8BrKx6YFpr
YakeqPt5soPhqPYRV4edyUadUUCLVjhQsJ1LQEDCismK0mhO0EDm4uIwYWof+PJ4
y6/6ZOz6uUscJso9/eeREo6eZnZBWRiwXb+onOM/Zzq3jofjmHP7PWxgUl8zeG+F
TdcIr01pLlWq4IXmZdam3/s3YQDMx2UBkN4yyVaBV9c=
`protect END_PROTECTED
