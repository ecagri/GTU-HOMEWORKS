`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
viikHzWh7Plw5KHYn8F/+jXqxylN/Nbc+A7Dno3tVKReG25r4+x1uT+c9a1RT5PU
4LgsyfZQY4OhqzwFsYEihU2dft9ngBJDQ16YKbgt8GXPEtW9kav/1Wuk1tnXDq7f
zNsb2SmVgAsq7+9h3BS4i079Cifi5t4B5CISUQ9FItELzUAroQn66g4wkJaufCO8
zRldkCOtuCr59RqZ8XMvLJ9EFJBIkWL+Li9eK7RK1mvxOK2pJ+iIUIymL9dtDjjG
SO1j7FL4+n5JNwtUenJzZICX79XvlOHdewyA73LOi0FjRHhFXE7fg2gPevAUmo+s
1M8nbQGza2oG3v7UzmZT3yn6aPgGoPabPKofKFnBsU1Im+myAUV0oz3k7IfEXGjX
zGO0x8faOy6YR8o5wzW5YTRakQ5rHmeJxsMr7P8SSjdYLVHIYTDSVMppLxqqpewW
B8I63E13jpBauTSU7WFe1es796F7m8RiKGwfnYatnvGy7YUWAd2dkx7Q1eIqbKVY
TwqBsaMzitB+TF0q7Bsz2PD8IzOK35rjUd9y3AlY76JjZ2nFy2CDPuVKyuytZw1m
U8AFr2BuTEd5l1Li67QWMCCEZKQrv/4zqcjdl87X9mpAQYMzWn8rB8+mHXycsptL
iiKOjQAS8qnK68apDPNZuL+K6RGYfX5wDmR0Ns29s0CVnxOd8aKbeIc90aGt0q+W
whS3iZqLtttsdAPMvKjsOHrFZCdm3gXE+1pKZEURrZpNUp9YumxL6xqIQAiNDwqe
q5VgdZVIJ5qgLG9jOEg/C5QWRk2copf2M5I0t0kz4xvvkeg1uWig07exO6Glyj3h
7v/SIVdFEasqVVqAdm9U1phXjjsSV7yDUoEwzM7XW5m58yW2R82Ak6oTVlxxjyNh
RtdlWf8j67Y2FyVeJCI7/RTQa9PtUy+70IY6djGusR9zYjmzfBXBBgav9ED5tUu4
YbcRc4LSdCC8P9ou71T46EwgxsovtfNRL9Tgk0oFJZjCi6fJ2xNvI/u8ijUC9V9y
YxmDjRMD3jRXROhlmijIux1K1JI0t9uvDGcL8Gc8mtB85AMcpeKtmfadviz5mev0
W4tIz58hutjZgNITYzZGBAHuRVe5nWslkfKXp++OwDODKsCSYsaGJE2DS6HZk2jB
9FIvAsqQ5YuyyqRkR5Ej0JcRuoL1cHI9z5sAJN1JXsZBmMVnADKxbyvttRLEikrD
R3oWxYoLfM4KHQkB0Br99Zz1ilCI1a5jGmGtdfgcdh7Yx17d6Y0Sio+V0mcecWY3
JOBaBVMb67OO3Uwtmxhn2KnWdPqm9j7LhyEOsJKP+s8HYg5ciuvw/Vy/CiL4sOPc
iXmr1cDZiZ1NMzpgM/hgAHYXq+nQ7kbDJU+5HDSiTEGNuKEODPM2ohZk6fS518WN
FMQEUVIBAjJegxe+q0wvcjnZVGFiRmepY5+PecqrvcHGP32q/+Hy35OvBd7RwxzW
xk9IfjylG5iq3Epl3oMqMOOGKkUaackasXjUYBkahlhKNTucsIrM0QlW6Y4hGXBz
W1SItwVHfpcSwAMlGte5uN8ZP9i9FDqz6KQ3Jh4LyI4jhKsAm+GAwTksyERO1Jf/
2b7ZKE7vh7kZaA7hqy1Zn/O4LiDQULn6zLJS2oMyPd7Wv4YmbtQuM6MBctmTP50k
/RK7EJ38Q3XWPnmiXEb+EXp9uRb82Ooy+MlWGI4FSDoeLZTvIDI+CB6pRq+O4gt4
W/fe/v0VI6o8DEuhLku23ADQAse54eud8dYnoWm9xkPBYOTz6PXpFVxSYkbDTT8W
vgiVD0LX48jzXnqR0tWp//XCqg4FatMeR0sxJXpKgHr4HPpdKTUw+7F0fBwYXVjK
TvlL+uZqsmtxLyEY0kLU3orkL5YqjRFoUgyYkdQFdsgV6Awq4KxaCZED7iqbfmsZ
W+R7QsTT/pPWN4goan+RDOUog2TXpKPHHJ54ubwLKQSNq1eOzft6jw2LMvz+pX2y
G4K98jO1wCJPDCKQw9CTwgyjTdXXAMBKpHzyKQmAIK/P00KKUcgpxN9587UuqWBf
L9Ygu62IT2VsyDuZBfvX9+vd44Fhu80KNZA3Q/tZzXxfzxYnHh3hHxO6SoY6pZOb
Aj/GnfkDA6kfbz9fiMlipfn0wB95bfQXL47HvayUtsSF2nuwR3kKATFwODxy7wxw
OK+eYlf9R6E+iBnj6KIGSZOszUsRBxs04v9EK13c8l2Tk2pdZeRbVjrsXEKauLcr
u6qYfEo+KjD/3CYBBSOSgBLGQPNr8Jlm4UVHGnQwTMgbgw8h18DTrka94G+kLRmr
omI1m7onQrrHkKrNo3AjXB371uOiK0z+hHf7bEymjoEBbFspLnT3aOhHX+BYc7Oi
rPvxLzGVBwfdU3rSG8HKutxu8wH+iuCvel6rY4HOFAq1DoWd6A68JHia474gmUTV
e+G9U9XB4jhMJGo5+7Ob9NZ5aqBz9fxAcdNEc4DtETP9HNsn+NT1dMnBApJ2jTl3
3O3CzHEz4/Yv6C7k7EvZijeFwGnHUpqYA6tAHGKlXS4FV1uQ2toz5gr4HnCWBQuX
Sa4LtWqUe0EntYKuIqMLoMkY7Z42hcGnIdqqJj4O9bEfPif0wR+XGZZcEEo8OSsz
BL2a2ppluo4gPbAI8rtYTq5VMTuTb/YcHk8tVV+/xZ8hDdglolmvrzB5W778a08S
YSYlbgS/tKz/FdiUJDdsPzuD1KdoDJUNdXyx81nejrrfQ9WTDixIZKJpX7I3+LWi
joDqndroYsxcqGcuVOpLAlcwlw3LI5n0yAsXebLuLWqdlGcsHbt7QjlDlF+FnsdV
XK7K8HdR2pYpaspglpIWMAAonRi9nnGjwf/DWmxuQv3qMCAUQ97SicWVx8npL/E9
03J3waXWVOJD8KEGmieDyH4TPB8wiROtWRS65miB1aqNvSy9gP2qv2wzO0/wbz5v
9eCX1dybV/XWsaLY96qq3hdLrWsQaZyKGHrK6F/+FGUrnTaLB8HhhOhXiDh/zgpm
aZdCen8Kr9tvv9r4ETbsDAMhy9s9np1CgaoZiSqLT4GDO+e1RwFlmSwXlwSJlUoS
yXsOudP0g7RgOyZrG8qJSpC2rqJ2JFnNR/9xAY6xu0q5wchSNInP+wC2SCpr00qu
ZfH4jw9N1iQzqtMU7DtOV00MWmwN2wjs/fnsxZ9OmrNx02lkC+ly55ZBWJiJLG3E
hhHtaHiwUBH9NfUukYXqaliXdyUR8lC+In58eLBXZWRECFUJDrX2MqLjsCYDhk48
Dfp1iwWwpvMGgshQMyFoiaL4YZOEOFDOyh/yyg++Z+FydOxc3jkDxGQ6XN4Xtr6B
GjqEfIAtM2tlpWXkLAAIMI+Gi9ETluD8lp8MGOk88hpI2OD4ZchVKU2xxNgEPlEL
1/GvyIOxVHAbTc/pRRX8FMqPGPkJ5lJQgfDnAGk5Z8usJRnyjP77pxojEB8dAECN
MO7A55vL8BjLpq/X+CzK8HHfKx4qcmzFITy3gnOKjEKhy3ezzUKuKRWZIP6nPwyA
+8GGF9HROaqOkbmsZkxlAJGBJNl911l8bF1FeTl7UNMuIg9mu5qdW5EzpFJnjRkA
AP7Jw3f+UN53JDQYEd3az6vR0pbtMjx8cKIUtEJ4IlkALcgX/DQIiWQB59/YSfMF
fy/Eq7CBH8Yfy3QiGhuK+kDTYBMQ1tZMs4Oknd4L6AYOvcw/au0zNFXSRmxUm4vk
fl+3XdXw2UJi1XeUm+wdcPd5BXysrmNP/13AJxJICKLl4r8OXi+BHHXzczX2gT/a
SDqpPsWMI1Yjk7mKoC2+VOoPNrHI2R0QF1+fIvRDYSTwbxeeJGhqRZwmPx5YFGNA
rzrdXeZfCpZeVvgXR6pS3RU+0zjyX1+Ao0mm7tRnKZTRJrLb8BsdwCDgX7Nc3VP4
6ijqIb0gtcX9Yb4sNB/NTNkhTsPyztG4BT5vJzkGXrQWubvo8Pb6jnBlsPG5AyWS
6lIlM7+qB7oyjyaNG64UZTU2vqhmgZvs6kTT4CuzdkUEzZPA+QD6Z52ajWUf71j0
367diLA64MxtTHDTvHVppiE2QEr6zoqRZp447xK5oBpIWDRs8axtZnr//HMRwWgD
M32NvVqSyZX1WQ2wlcwK9afFgKGqO3BigKSO6eLXG+1A3y8dTS6AyFGiG+E6WF4m
5rnlA/9bVWU/8SFO/FahSLfLDQbWH2cBbqwxalXxHA4gPRra9jvyoE9INI2BymBx
4fEfRrmuWhl/1Kmrz6eDb+Xejk9lMhkuwQhLCti8vtqopQX6Oez96J/yenUKrmed
dPyTxZfg/Js5dhVYEsPP5+Er8IQ1LfG+giIJXo97Zczj21nueoGFUHuaqvKpIJvO
KSZ7v/0pE8ttsihCboXdX6D4w3KKdrzYUZL3eikxBG5tgLVRtOYn7e30G0XiFkh8
/CTOZyW5j8PEyYJv0qeLJorMi78x/jDeXWlF9BivEJzveFkfpGGt4MFBdXRKZshX
0v/zBl7cH8kuAttsTX76a+0eioADQ3xjzt5IVpAHjySxh5VJBJB7w5+axWony0t3
yBpTsPSLoWJkFiHMEXcWwzY64AJL9rNeUT6FZKMplcXzgPo1olJF1cNm5F4Y85vt
LfmXgEJsEmhYEjxZWz832PcTOG66IldYEuPuTNgCAWf540UedYJaitjkY3pIzqUa
N54iOyNPORtczIkvJNiPasEB6Hyce/wkSuDzYjzMQiKf6HYkL4Oc1AmaBlroBWg7
luRKxH0f7MikrCHYsIqGV0vEHOy90uX1L2+dKTVWyh/kcESFN6/uG5e08M4EO6fO
DY+QPL33uHBoY+zkuIMR5W6ciHo9J3YdDt/URhW25IxlfP7FpRJhLTBt/8JST9Zc
oqMs2EU9Xsi4H/7NjoHlA54ROXM1xa/rJYFmfEwmaj2buhQ9qDcAaStD1cE5/6n/
myiXTE81BX5tpVVC27hbz+vju9WLp5W/NB3DSQXg5jjlv/wYLTHDlgkUBaDttyQH
POIz3v0H/xO/Wkxw09lYR0g9xJgcUC8MC+mIYgu3BrKCIbprWLPR29o6IH5qryu5
oj3W718ra6uUDYT+POUn3tNJC1WlSISgG6mm1CyvoQIWtZ2T0nq+Dua/Tv/LpO9j
nyC7tPxrkbB52rDsa8Hg9KrA5J67D58TgLEO2SAYbCXoW4ojLBW3lzWqmbGRp8Zq
5ogUcJQl4Uj6MAVHnCeD/sJexwoUqQj0BDOEysZVefljyCFTbjuJaoFkKGeP4Abr
FjzBtiuViUcJrhmxue3HxSmLXAbKbyf1eTuAzfi+/zWYJtEj94LN1pdRLQ5AetFX
gNTFnGSOKsLlKPi2t0OkgdN8Km4pJCuOKyiM445cbEhgrMHGxLUO3/A1xfEGmax1
+nURtwkr0FIezm1P+MwKmW/FTX3k98BRKyF1scYpvTkQcx49ZJEuNTJJWG8lW2hJ
/RzIrLvMk23y3jMIBcLyH3UO4DFBi7cj8QBnYaEP3bB+sKynHzgkd40ZSX8VH418
oBZft06nmUZEdk8AaYlUBI0AEzqkpucIVfgNDV1tLBGoeNFFS3Ddnbb/7k+VjgZs
6N9VwOT+kairxp4lY4rK5/nynOYvEt4yTSECCjHqdRqXr8uhIWZ8TI7NKycB9IsM
abXKrp61tM8Pa+3ahzqNIXkvrInde1MeDp/dnQ2WrQLImi57LSIucth31SncWrpQ
IZjvG919oCquXMUSOG51r70w6hXWT/25s1toqPpyg1TUwUgnVGaiVorC+k22Xkrz
aQRWJmK31vM/LNEQDSXwjyEb7Bdh45ePCMApRGVHz0B8ztLzS7aVkn3xt1Zo74/i
JuXrn78FiVjLC9p+P8QHYlBn7bKuXrjwpiLNqA/QglLeV7ZIIVAAGOkYrvFX5ke8
72Al60mtLTouFAuCsZL8j9YaP0T9kwFJS5MbVoYaBLV4RwiUD2jV7FbvxTWEarMv
j1PQdtLworn/AdJE3ervFgU5kW+4LKTMoVMTLC1EEtrCnq8AFb/htxNiyTQTrIOv
2jNBZsgnz0IP8M7WREtnpUQ9NV3r+kB4c00FVByXxxxf2B0OIFRgDt3h3R575JsG
fIYI2Gc4Dz2okLbuKbyTibWTn3cKYUA7TnQwtjRB9FcWKHmT108isalw/NBq+EEX
0EPoX4YuYK1bQQbMscEkudgMjpMew/8LYRDMT8Yy7j5ve4Kgt/FcdX+YMBlROs7+
y4fjAH34vk04DTJjO53t2TjfuQdgm3UvHZTc4NxT15O9EjEpf1EpWArGfL4nSMk3
N5WmOry0cUqoJn0ssHXAKp+uynRl3B8SMiOCTFodn8VCSYICNpUq7XiyaY35hLTi
aqY1o33sWUVAa0DpaLv1lxrzgXzDY0Vs0LYUNmaS3si8dO2Vt0FUJQuXB6u1j66a
jF+kT1weX6tCHif6uT2ehOXvpxQUSB9Mc9xC1CHalQcU/2g0bc0rW6vDNWE+1THP
uvsJi0yPnx50zcUXTXVBy4FFeFDxa8MGnC33KvJAxQqaNYBH+FkbHDqiivg68jz1
MzmNa0DIRa5yPciOim0lpTiW4uakKhMP5S9mcg/IwSagsTLoTZOMWoIoW/G3lx7S
J0J/T70c8XPGHQ1cLdW63gwHyq9XKH4UkITYblpuIa9tMRuaLJA90WsTFMsgC3qI
UKODx6f2EkWbQavmjJaUpFsco+gWXo6W2dTzBa97R8hcQSbZbUjQEAa29JB9JCrm
NDgq6TNne6QYa8G/rpnjKOvelbBxTOO9O2TWvi6dHpPz/H+HtgI4zhk6lsQQBHIc
ahu6CndjZYil6OfxmgJJsVoP5ViYZTMx6HsmtQMVag5fbaO0QDaiwSv3Ywpjsv7O
qHmiO5uhWl5YfU2gNJdWLNX2rGTLmQsN7QJscq39zcS97EMrmiD6glA5QAmZbQ5w
a9EQhhQZwsUd1TIEBY4fdD8bcNzQVn0BBk7eGb6dAhqvOAyPYOAh4BnVuuXaonls
eFJ1pQYEFVFfNfekEkPX5ThNgxl7GTSm0hp12WSqa5b0XObBRQOsJHSrBvFggR2W
aQXuy2VEUv1sX+laKiTg48Y9V32iesBgQCQ5Fshgvq5Itni/srgvnbdMAnLT6wpB
RqeZhMwXfUuEXzs0eKbhnBZMDgMdSsUb1e/cEFTlO0Nno/iGtTydauNSgJBSR+k6
u1H3JEIubZu8c8PybGZob/TeUG9iPUw4iFmYbY+SezULiKCGSVICuQgxGwF2z7ku
vW0fKVUbEEbHZN91Ri7JLUwgxSjVKU+af1xNGdCgz2r5Id5pKvEBgklPnlvnQboW
uafQYfukSYqndbn0SQtHRTJEojfN7XprHxYtnjYxQ/niABsu4l2LBb8se8Zb2Pt0
/tkrNMaJxtvpnpO6mr6Pq/PKEvafWxi3kyaFDSX8Fdm4RCEOPa44anhYEvVDyT1Q
limmxqzfaEk8EP8ykEB+4xGafuj4sS+T7auYv9eN73+yOK9TDrYUWZlwuzOtV9cN
Rz4BFfgmnWyqM8NvaTVAmVEKc6npqLJVsj+IutzzQOGb9Z9M0P3UHgTbxxJ7qmsd
9OqxWpgqg+Qd+MmiO1lLrZHY4qDVTBJZpni/X/OQBZT04mt2e1TvBkH9q6LOtPoP
feXmYks8+4qXqTWqu0Tbo4tY2gv9+e7VQwd/ydvsnw77Z+bU3iOcoJOEix37wG9S
lkfUISR8q5lhpHQ3HCJChYGNqrR0zyPun/VLwn1l6Yyd8c7AZ2j94wSfxn9TU5mr
g76NkpWmNAYgJdaDO4o7Qf17cRd4vDJbDah5+3arN9Y3eCXNUUpbZOrGFvG6SwnM
omtVSogcV/bg2qEjmC0a2jlod/6d7srUnw4zWQWIdULvlP8oivcjyktPVu9L7hZW
lRp7jSM6VyBWzkBuZqdPdJECJaGEwh6qusutxt3Bw5ITR9LiNB6ojVScfCyC9zAy
4vPAZ78Z4jDvL4oWswGkPSTIJ90mG45wFbqpXGSJrg2ZJllXbR9h5NiJMETXwkix
fm+8iVJK/VzjONjOAorX2cNWl19MI/42HDh6oNlpYBIgg8s52Nx0BvuLl4Dva5nX
hQ0UYKie5PMZ6X65YSqNrSTADLZwXx5v6XR9EXmXgWRElv0n7GYfyQ/1DheKB128
firL9f0D4cjVvjdUChxRoZgNLm3e/7XvhWGWlqTgEjw=
`protect END_PROTECTED
