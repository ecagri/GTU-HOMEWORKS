`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iT2sMYRTPQxCWjBXJAa5UFNEqvH88i6UO2+3v5TGJLiYeabX2zXS84bF4g/P1b33
AbGhNBBO1E4rPv2b1rk2q18aUuhxpsf25PSahUOt+GqGl38Y38D4el1tB/62Yfay
yvoRoXVmV4deXclDS1Juwu1j2J6V8UWMz2DS0Qlx9/GSFK5ey0pvdPLlAj2YZmpx
qtjhJcl4KNCgBLc229qsZEP7FgUiCDohi82cJz5O38AN9xcoRtIfu9FOkxg6loTt
lwk4FVIgqcofq7Yut/fyiOhBtZns3vZWf2FTAfqKJj4bCXcmgUMFL5GqqUXRn7GD
ufp1wa8LRRs/1um6+478bdXD7gba17fdsIQ+WhOSnDSWOGYK5PjaxEbvuH78FvTb
GJQUh12Yuj6vavKgukJ4KtfTO0rXQXeMbybJZ7b1eDLilEr8bUYXtAgsNhzZvlSp
9nuz+IDfIg4mW9tRW17Z10XWz9oN2OLvxmXdxJ5PvwECpVC6lLccFNFePLu+rVaH
tdxfRlIMDwFNv11GO0cvJF97HBJti7M+hawE19bqx5rjY2JiVPpCVzCH6qpROB1J
Up9LpLvwGT7nAcpPKYcQsCTTPk1LAk0P7ltEKD5ZRSUjUKOSc6kyVRNuDMS/TFdC
lzgFJGDeg5CLRuhxSj49n9Lw3eppZuuhiHJ8RfBmJV9xrubt+i9FOLkmpB26sWHA
DLoi/D7ISA301U1UW0J9a8rxlTb/WP65OkT0gUB5ouFFg1cj0hQVaVsYFlqq1VxW
OV2qkEwfC+YvAwSsuq31DCo+u/a2FieSnlSyr10Ejto2Qgg5oDqW/QHgQEKUfTnD
FsupnpgCMGh8bKrWaYVArM7WHnWYVDzgvimLhXP58KXFcRLy95aP0nb7HYg5QC8V
efzWg8nvN3JG/8v9GFaGiJ3l3nQQSJDelE/9jgqBttedTFFYDu9rjgA+LQWJNtdI
FbsUOu4/ItXXIB+DzYH8NK9XVES78SwfKMRRkRrMk34ZZa1XCoMAbobd0DYQicAq
yMftarA6UrQKtA0Ee+ssNSFjOvMPAzbiGokGSTkV7DlcQ2wy44+fwAPiaoArxGok
dm9TM8PFiRNb7GDWFLNsbcUwlw423iAKzdZOoezJKvK4mvowW8IySZ2eFWr2BJXF
k3cnOPmoBN1RT+Y2ueg3CUOA9IlqmedGwFSDwAGd6bscHlG0HMNvKtInbdVkAs++
qTT8e9G6T2F76+30hrWxGf6j6ihfehCRZEFIVR4r3AOXDpJTrCcZSKl4zwGBcJ82
ymPEGzKd4hDvj8TSZj0bzKih716SsY1g4vQ7Gnw9e9oKPYtdpl65PU6m6reE4lkB
EkiBY8uycQ4Inh0NOZ0j7TXn3uAhGomF5mwz4+X/haTa/dZQRSsSqnDcAiIPqJjQ
l4fwC5WugD1iLKzSqfKyUafaYcaM1mubqwS7SlLBbxfJuFy011F0fzFiC7nSAYqa
DiIaTLMl5cTpjMmmF3G2XmsJDqCszn++4Im/PGxfSrVryFxQtBBnLk2F+0qXWfVj
5AeX2t5PZK2JcLtvjUEguWAEEmB4YhgSUaayL42r2/7N43WCnrGwC9dKHoZgVM7/
e24xPNbDAfXTiSgHYZ5rD5RZDeQrh3nMIwOK3UXhpEyz2WezADnjgOrRdVL6Gh+j
ZzYjUEuwlbYxLNpkafRBNnpMDrJh7+wGvyJY27W8L19FFHylAJz3YANOae2iIy1x
FxSX/ZfwiQiz3Ml0eJReoMTAK4PlWuJjb1ubg3nibenx1TgkArtYtW0B39TqUkEq
z7SHCaLJx5PRg7JxbMlHPXlPvlOhGmRUMl2szSt79OKANexYMdqrFFUcMjtanmXy
u3gaCXwQnXVkrqqmth74MscGjjL48s9t/2ohFgtXYK0VXCTvyYuD3eTgP6bssOri
WEQ9y9SgVKzYm3IAG2k+348npX9aKRu1kfgpID0dOYc/swgShXV9IRlg6iFmQr4J
ujUqnmGIjTF0DD2eBEcE3FzeAC1MVLe/tYo4/6fCBAKP5NR5lxg5fzEUjz7/sdvg
xzpGXa3ImJyfblrqTFt+C82mP4/p1zEHVKjUDgGnynr83NVai3lekQv3q6mEd45c
ItWNkpMuotn5EUGkUVJWi3EotlpSBN1FEbYg5RTAe6/MJkVKxPIc02QW0AOFgN8f
CiSrTl80We+9ahCrZlseGkd5fqOyC32elIrhxJu2wKg1tX6hfjYIg84yv7OP6Bl/
x0ikosBeFL3/kWmbp4SZvk5KwSVZl6X3Oc6R9j6FJ27r7McqI9Iku3oq9xms9Q9I
RdKJdd0nmOZqm01+xP46bxdiBrgL6XnSZ8qdiTc0ZSpVhGUgh4pYip29tN88ARwQ
KX7ZlfMnOQrzdeR6DFprM2G1FUEm2/l4LCJKoE6DhpjaY/FVpJVzW9kD+1MvYXrO
3Uz7h3DGCNML9J4PVUfAWYjDOU1HzdsgJF/8KdWrJStWz+eh7qlR7PMdww0lp9IH
2USbpxPjiBYMQ3UOJ/kOQ7r7684EjXSrJIhYBdbjlXJ6OxXHGJmUe3FholWtxYsa
Jeu1qP+0IkdZxnTu3V2I1HYYLAPtikpypF5uDYTg9wk=
`protect END_PROTECTED
