`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TjWwuGo/JgOmW7vuyHcFcGsh5Xfjty982Ayjh8pV822+lZLCQA2DOAzsOh30zu+C
C82ItwwwGTFUvrL7BZaeCu32zBWxD8eHKuW6uyIWNihYKjXXgkLR5SDNOCljGwUN
GLA6hNqUm27cGBN48xJTgMzOpnftZmydYup3JY96gLjzEiYiYEjYSoBjauT/kvB4
hlPNdTDJe0D9/7VMwhrNGHWNuhUYQNottBbSMr7ZveI0Nav+xeU4cRUgMYH5ZKlu
ewPVlaZV7e+9S5TKxRSL/NxJszXW0rhYEb4flEkOu0gf3FOQWLnmF9m2G+RrZ7xN
xw4OFWbKjvHhXxb3ux9/lI0/9fFDQ9tGlMTVqM16k3z4jXLHqboY/sNffKK4DXQ4
U00CFVSns+YoDvFg9Xia2kbD9jGCVakqkrVLgXVTEjB1kvZxkaR50+NGo9ZwE3gl
pOH9i/o8tMP2OmqG8u4PJNhf+YRT2F1Nufq+H3kd7qFlOtWo4vPsr0JSWQjvtutI
etmsjChM9F3bKcznqoXL3GEpv69WU+lHpQmrWThZW0l6nP1UjktBxaY1BgHllzDT
IxbGJCYpI0vQbeV9N5FkZAmADVA9a0Uv9QvZ6KdhSDENpIRZ4qCDndJZp7ZkP2H7
hAM99SkRq1enDEPoGWvIxKi6oXdq/QsfA6id9W/zbjK2eaIchVOxc7tGuz7tFBcr
6W9cQJWV9OtIpR23CodusxmEQ5X968RxSmGNMsSZKUKxoF71SgC6u0tFC9kHvPHD
O4skKl5c0JWhoDf6frQveZln6zg8iAsdw7ewLyjUUA9OWHc2swDhdUTXAj6FjSu0
`protect END_PROTECTED
