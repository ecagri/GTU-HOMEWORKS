`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6iPbcaTDoqoukvl16ruI1Xd6YksiHuvgkrxTKR5+LTrRsO0Codyn/HZdxO8690+v
FExMzp+OlwrG05WBI0ih48uilj3J8yyXV6pS5DWX5Q8vKXI1B2rWNz360xLBm39c
qACrGz7+TkV7dhrPAliRbDRO3yvLj5RcSuNRydLMZGjqoz4zkOSf/vPLGhhCf2yL
C7vpBwitkoJkI4hL1uY3sEq38eBKFcU1/nnj7QAqYVtcK9ZpN4aCUzys9auGxD9x
Q0WbRgF1KdY6lMv7jmQF7PNkNkja7GpG1tOZPAgFXnGqc4yCXNyviI495a8vOO6B
UYAqVzTbuxaOnulQ38GblH/W97MgkBueBsmTJ0lUpSzHsh92c7siP1oPbAwDvkwb
8e9uD/Grqj5If++e/1DvGw==
`protect END_PROTECTED
