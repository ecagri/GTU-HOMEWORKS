`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a5G0VRqR5iTi3xVBADY1XeKuTC/6SZOGFQi/OvH3cjgxAv/vRmh6Wf995cpy44Bk
JA9/psdDuMXYYkTHWqLoXa6++fROpx1nlYBZwFasb4WWlonWe1o4U0b1DbKF4B8z
f1xZ6g3hH8ADZXPeQy4T25VLGHd2v4QIYwAkqdoLLUh0yEs+8gZRAnjCn4Hme3lI
0xOz7MyRVK9sXkDf+B/+Rw==
`protect END_PROTECTED
