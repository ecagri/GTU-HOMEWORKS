`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sxti/LZqKdEbSYijUZ8Ps8DQwY6S6ImjgKVnxwLfXU/aexzEBcDgG24yl6slDOFa
JDtlM64bgPkN5fGlzUxwE7rLdIewgXnyE4d1TTnqua3Mpxrq8L4jwLrZEL2s7yjx
gAjqnOwJk9FpvOatlwb5WtTJQ2oLiZOQEI0BlvODceqtzh7AoyEoSqzj7/h/mtKQ
rTDAikggqe7dAry7LELcs7JZee+PCmhvOUyCgQs11YweE00MEZkt+IpYYjLFRDK5
BrVqShC2TQx6YC3kw2Pn5DH4KBnJPX0yJi8Wylljla56WkbKisC2ZbtKKhlPrSg+
sO5jNg2WHg/g8WkrXFiwxlEVy7FPwFFT0Kep+aweEZp3F52iLQV13yw6bPy86O7l
2tTxWqiPJB5E5iuq2acz6UTi7yRHESb1htXThD5Lzg5osYCT/04DhIeXcVCuyrOB
XiazbEb8zIQuVBwfKGLC54FhkOydiEEE8HjYdrhkl0bql4GJoA2olzPi4RyPNqpX
GjiFOWec/SzCfI0/ueTyKzNbfMnhEIWGn5rqADQAY1AAm6KKYEaNDwYEtDlB8dFm
0N/hYh11Yn6qsHVjf7hWqWuCoGwbIXEeS/qPGvkU4gXrlz3QwTvaW7fIleaVOhb3
I1qRJVOk6zv0LjsxLFZT2azIlPl4JuXVSgbJtzRiP8v3wl/4r6yIrfo6R5rOwn+O
9scswKQ61wnZs7763OXLtpdu2P3jXBVBV6V/Br9PYBr99oP1fgwMpr3t39hhQqIN
BekOFyhg1FEnO9l8BX7mRNY1emgUXCLb/6w6UxcFBPBHorWKR5aHSOiTEaT78Nn1
SFq3aKx+AKpBAAxIi8CEEteZny0tLYIbtRSGB+/fRgfPSy43BYbD3oCpKIwOho6x
5env4ofBNv5eirSMkUc/7h+qpQXW70kl32mA33SW588vuYFwP+HK/xk14Y2hTrQL
v7+/UNltkC5H7GVF4DoIXcRefa92jTw9dVCT+x3vguKTksaqRfqdjIS5fi3NpCpY
+b7DFJ6DiMsoGHDquu9lXtmqJLzl4K1tm2Zi41raWB5pTkE/fkTi7oZXGVr8D5Bo
nHLvPmvFzJLU/WQBl7eMig94Ru2TWbu5PJreGmVuG50OSkLH1vWzHos5TarEqTLO
9l4UFDpYxa7gGQItg3OuwP+vfAXWmEeW1RBsRGOitV8rk4EdTgsAvm7IQn++2mMj
v0bVyV4wI9OEjHEheuoAGUr/UEXziUOjgu21R+xU2CVnPa+YX4USJkiAOIdv1oca
aBlp0PcBTXP4B54O1RasiAppdGWscrEcda8VY8lSZ6ERKmTrwPmbLa30dRQlUjz2
pz0u3znTYswV4egLGc0qjZNRFvuTPP00VPgSoeLTf8B9LHsxO4rwwHnfPSTASjFD
FE/PbEyKeLFbVxRKxVMcfZ+OZwi0lMVSxb54fSJTBIctQBMryMWoRxjaF8nfaUlL
mn4ElfszDYoNoAzbiOQgDcG0X3wOgQoP5w4EGj4YculiroEplZ0RD0UOu7oMvaso
U6J73lYlKkZ+YJpgvEQtr63658vffnLtk+IrjBWVDF9fj1DIXmXJYJN0bjz2Jcbt
sxkijYmSwBA595/tNgew1s5yZckJVOpjayupMCJRG03UCnXXyFlhUNIWWVtU3Dig
HW3kjHYCB//+r0o5GJaDoLF7Xji/EX6YGcPFUZUuOPICThG5rLLsKQ7O1H4/FlMz
yrhJp5xBtDyw8o2k4jsePpbCKWMCQlwxo9NZqaDqOqTJYSG/DFRb4SbDI3F+nDUM
nObPdN8Jz3556dZ4DxwwJNekZjTeERX5/kH3FWzUbDdk56qmbpQNbsY4BH3HWo0O
5QubAXpQT16OnvksONtLI6cenUCbB1o7Cx52qppEcGnGNf3uX+R9m0TsIsSUC6UB
HMRNYhak5UYulerEo8iy6wg37hLRWUVyeG/dwwPsU7OBvf8/wkE63HxnDeZZ9OkF
dkwMek+xvhIc+9CgVl0uo9CV7VXu3RYZ9RhRhizJFzm7VKxIgkG11SMts4J8XyQ8
SIs/Z3Yi7bR9kIyQwHS3L9C3L4FdbWSa7Y5M56goT29Bw6m41u91MC+tg7GQhIIa
mzW7TKpM7huMC7QpyBNabcJ/V8s57PTyzTGgnxdfhQn25ZBPKL/Gsk0hm4nDj3MM
hUNA1PWoDjYmDW0cVdHlR/l6uSe/UHB9WHjKR9h0sLc=
`protect END_PROTECTED
