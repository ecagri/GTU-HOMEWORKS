`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tqcUz9AJkoxgLQUIT7SrbzxTMO4elpVqDaaoNlmQj20sRHngsLjon0HyCI5p+CNO
b0VijF3w4TO0Y+ZzfjWmHcS8isUtZFpXeUSqKdF0JtGUJiLYe8/6AftnBVC8Adi2
Xou4rNF14yCpcyTMDRhlhFNxwP+kifH2t79CviJ/mQk84xzydP1asQolNAf+SN5o
iojG6Cs+ssQ4ec+4AcztbAwKyxZUAU6QE0Z2E6PwFKa4njXExAnXv7Q8TlYRd45X
VoJpEZwjm/3heQPPristp+PthGcwIbn0SrXnqTwnMAXmwbD5+VmPl2Kxpr/cHQKW
8E45mVHXRin5nZ7rzxefetzYUBQAF6PT+n2YlStvGqcbN0zWoWX8xi320GLjfh+P
/UD84awmKHvk1cQWLSiET44dDe1vLIMPa5czD+C1KnwfrswY+2io0nDbf87p1CdG
dNHT0uth5EJN5+s3hKXccWq92QoS6cNzUblQVo98aal1PZKg+tuexACa5cm0CdWc
nHxtnifq+4+wAwEUKax7KhMAyNFN4s/IbZbtx/Qpaaral7Qfpzv5vtu6/PZcUojj
ZdHfNjUTQU6VdRP4dJQEJGZx/bcM4WSEq+5igeLZnEfWjsuQlTRpHVf0Ogq0kbp8
nL1k1PMLsjr9C5oNQ/LuTyHhgnK/8GregFPegh/FYuJKtb3azmcTwdueJSRTYObK
Tyq3oQxdJll3p9BW0HK3+kusUvmSDKWpCYZqbdMIp+TWviacvu140ebrKrXRkJuQ
I0u0Gvx8+SDK2ONlNPnA+wvfnXSjhpwnHq4Scnd7JxCDXtjZtma5SYJWpwh4kqI0
PZCH46zccZrFu+nb+OW17NNrQYUu5cGT7G2PChPFr0ZzxXCeATUNiZA+KXM7m4fT
cq38njW4qkLfwBMBM7udTjYOVe0m7wallVMCzFbvDJTqplbVusxUWBB3O7ViIIcy
cHpMVa20D1rgVYZTI8F692PytvomvpsNCfm+Q3XwEdi5EPLxAjRBqAb/F1b+O0AK
QxX98yRP31tpz8S2MN60CDeaC1SFn7qMVvCTFM0j54d9bYRZ16yqpgaSJGXe9Z1/
8Hp6HLADehevrLRRtcgmasHYlze0O/YqzVzxOE5vTFJp382rcnBuUzrAjMO1uWnB
f2l8ioaszvZoqS6vHjKuEw9xMfwA/7JBJyXVSeaBMibH7FsCTwzGySkOfjbEf6Pr
7klUL2WmmMZNRKBI7oCU5/Jz15oJoCEhDnU8Au49C7cBj8A55XA7RcubdUgbQtCP
LG8tK40pgIVG6L7Bj26UVaXLeO4D2GqeriYhMbXuUWFhuBl7yCEr4e1RCuMylVpu
QS0XLY8036zL05n7OH9nRpFZrLYNu1HlbfBJF9cp2CNfixAaXXzmWIji0n7gL3cc
Jcgcu9+uyn6drO7n2AX0zMgYVrqRP9Vhv+q7sZgLkrlEZJEbK0Ssrl+MZJwbs2WF
r7P9qh377hkVMBCYbeHlcc3gRyK88kpXnN4ZKGJLUFzVf+g8yiHzCiaiUtjpq276
9w7gy4LsjCRLsx3B+s4E9xTRjxLKa7p1xoQ2GHenZcfZUjL01vcsOMnUZSgZas1a
+W86nytv5X2NdgubcKEZOB9G93C6AsiJW1+wT94hYcLHBm6kPbIn1MBl3hP+5MbX
sLZk7fpDnbeBnb0gAcn5Ry/FQ9UePHEfS7Kbf0BT6rg=
`protect END_PROTECTED
