`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/2+VYM2xagKo9ZGKwRlh47wV4HOYcSo2tEn0+3i7oHHlZC9dXor1DKrrMCwxR2v0
V4riO2evvdnTQS2JT8xl9t4RAYSaUqD999Q2sOhPvQV7UPe6tApny4/rfGXiF+Tg
56jzCTDmTcYrigqHYwEV37JRB5u2CG/w6QWmUz+xIqE8j8UHjK+MxpvQoQdMK1ms
T8OHcgOoL6UMyASj8i9rYXsFYmHUxABvrr0O8Yfsr7d03qzea81q+ByH6rFOU+oW
1pwm336s1AuAV6PMFgRY349/lvtsM9/sm4Yn/l0sNGumJtxciqfkbMX2LWXyg73T
oyIa732MDeGGLLKqn/IqYKP/jJCsWvMPy4mQLrigueZYb6qxpFikExsRdiJlwNXe
jOlYhv2J28Of6DEN0XXYUhw4WRvcK6Z7kxnQdEK3afOKKLqBCqdeI9UJ+wapsLtK
pDgq9jXbRZDz8I8vSrMCHr2q9VtAcL2igtfAdy3a+tBnVNADwFgcR4WXQI/xtSgZ
RHweoAEpwHOU49zppsAIIfwY7paAN/jzH3e9pImI6wmaC/3gt7j3/TMWhb3/2Cy9
3cbLc8vy+n3YmmhMHV3kQNoH1XlICR5XMnUqtU797uO66oGYxZf88gGTp5EywUZd
V1i6jh+FATFrOlPq9DB6MJPkBTi+99npA1fkW+gZ8BV3QKPm4AnxbPFfEXEeE1qZ
4MKYXdVKQsWmZpdNd2O+G3VSCy6DVAl+BEmor4y7beMsdZ34YpCfHESKI3lCTJrr
SI2CvWAgRaJaJsOTgRR4ABb/7VmmuF7oA4l+TeMi+KJQnszfqspy6ZaZQKIegBJg
xxOvGzBJ3SFa+0bk2EOEbyHhr6ggWDU4nvdMm0SXQgVtGFkhb/LpuUN47KXnOCu8
dvJuHWWY5l8x85OWl/DE0CJdnX6R2WKyEjwt+ecBlIj5upC6c9j9IeIensXlPmsx
B6+kGTynw4TN0/TOduPiPTjCmRJbV0YCHM3jakbT/lP4LIUf7oqIvt0o3iiC+HhK
BkMZXpTQhLQlna2qeTDZqPd1QE429RDVb5iUmhyXpk9h82wliCTsijkL4qHhboWk
GVVWfpEgVjptw2Lx9+bAMMxmTKDApljUA2V7jFXlevRnyuN73B2jv//S+Q8lx+mx
iRCs4kFgPVVm9vuuF6YxMWuXTAh9hMy42XUIbk+9Ne08yhm8oJZidblq1VzkXABp
EuJhqRqF4LgfidY54ayWjtn8syI3HsyMXIxAbGS+dl5dtcWdNPc7X03vxu31OznB
6AC12tEysWc8z4CmdN7wnZ55Pc2PuVQBE8+jWE/q/di0/pyF6iBh4SjMqtSdlzdE
+SvW12QhY3znV8DYVgNX/DGQbTcDeMz1MK40jPKx+5jQu4uVjYDDBiPMa4aXbrFv
dzAxcrVQX98o71xbcr6jEqoWBSxFHKNGzQIJhginIt5xN9HmdeKIqpli9cwklrh5
obMb0vcD0jZzETphGogXmV+Weywns2X3wmlP0RmUSLyKAtzeMCzLoc4lPttPfxZa
RU4RpmGLYQjmFPXGt5eYspA1JEbildtj3yeCwMBpWwNOIc5wn9YsyHlyFHi5X+wW
`protect END_PROTECTED
