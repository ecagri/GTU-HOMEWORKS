`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uct4vRmTPNfJ/V/wORvaIs2Zyy/KDqgGu1BGD0zuFDxJ4uawep6xzQdN8GJqWgDx
ZNIKovR9VQCqodz5ohOCuntdi3lR8DxZEJ2/mlmxgH7jsAeh6NPbUe//IEVV4+Eb
+1hZ6B7d59CKeG2eTvEMP0/49cUFt3eWjX/5WD0hVsfsyrDlNXMdueAxvkp3kgRa
ToWJ6iT4p2stK8VyhupHH/zWd6nmxB/JAsemc0/qyn/37D91QEyC43pl2goOOJ8e
B/xgV8P3R+mx3qUXCVRliLGQ13rCaZQfAqLNDukCFDZ146LLvwXjQwn7Boqd/66/
nlgYzVY/kEtIKuqWRzrKB1LAa5evRZhnYuhGW6ssiL52OZ4Wu7UZby/bS1WQUliy
FAOF5IS2nG3gMdnntfxR7uKVtEOJvzueYTdDa1Q2adom89aeWXL8U3jquS5zBjMW
8IE2Q8sCmCkJ3znA3VVd9shm7uAIZ89gqbtb5ruxr2QGoieppykqmYps3ejKeOrb
hAKLW0K97zouxSae/CikBw6HGLac67A0XNRhPm/+XHmKIhMyaxuWR32lL6dcJZVW
093HS1CE3ZqxfReMhwoajE4Nr8H2G4ddDpSV5oZuvxguH3oYPJcdu2ac6ZIfsJKp
q8OtvKtX6weobxJEBYdQ+4BPeNqF7uk12+5EsUigHsNznTEixHXpw3PiojcXiqVl
euTOqfHLojIk9jUc7u3lk2mGGZjBewnLC67V6/1/v2hTtaDfiSpQ1Z5e9XabryIh
fQw9k6SOc0g8VZ+duhL10b8Z8vHreyMojkjvS4EW4eLQ+5PodN70XnDQ9sq4yO7H
ZLMGnbO5M2gHrT+AFP1K6wpsL0G3rB8xZPm0WhQb9+7LeWwb6mmCF1EaRlUXnL4X
cqL9YTdWnOEFrGJYkFzYLv2fYPSBzKqA0Pph+tRQI9sljmoj+Pvbk3VYQUw6tLAm
m6QVwgA1UYrY3bbYZ+awfW9m8x2f+WGVzjYuDmrpKW3NkjRUOZalzVPL0UhkkSia
/HVBW/lffdkUhQkxb/kffjWSqGQqqh1vh7iY74TiUbp1v3y0fhmF7SBW7EvemFXJ
70aJXxZolp3CINqoEu/T9Mqf/20N2DIftK9QXVe1pXnYnaPBdprmorSBAlDRVy/p
XG8hObH+KWpvHTxAE0wbwqAyINPcqzCMMmwWVBwOtU39LGHTrWb5YVUShpLmsGvU
q1Fp04Bn9T91SeqGJABJ2tA0XoLzUqtTQYG1aF8aUmmAVrkLTH44YXBGvf1qznNW
EwfHA49m3kpGZchIhWKIHl26G2W3/fypqqY1i9G8uEaTtaLCPVoiizD7zpGXJLF9
eVQNo3W5jxqROXNletm1Mg==
`protect END_PROTECTED
