`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SiDVETHATLf9YmZcwjLzQ0qlP7G1bXGuR0n3WL9wtIH+c35N0FgGwn5C4aAGEQOH
QLcEaJSs23wDOZ0FMa5wdw2ODGgF+AoeH9+PBwoSBn1OyFRzBiidbohSEFOhvDXg
Kqa/2F3WQnchQvDh/6lYp83YfhDjtc7BzgNN/KP6AHMiVW9qmyFNqVZTYhxr1PVN
dRsUl4oNje8bg/a6//71DVbsBPX5k01BqwXgX5PKn0bnhoiWNazRFOcWImePeubv
OIkFsth5Ga/8/iLl1HYl9NFoNAjZ4Yv5aOBslb7MrFfw0xK7nOk7karEUUlocu3d
+dOOM+jZGUOaKEp1vZPwzbwtomL4U0Q+21IPXgjUkUOw6CQGkp5CS1nTBSXnyC5a
M9DTMwDGIqJq1dCBOX+1cTSYo6U/XwopznFU5LGvTNFfUMbvFOyHBQSdSw9SdCWV
UYSsapknXrbHG4p/QhPRYGvCPGNediMOAC7+Geu+764TmQtTPy+PVo7xPkVDwwHH
84zbg+OhkyxHYzpbbRDN9KjwbXBL+FIgqZI7gAk/FHOQsdXjgGa5dwBY3rsGfz0A
`protect END_PROTECTED
