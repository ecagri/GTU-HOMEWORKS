`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JN6hNw7h9KEEKD0JGE/I1TUDoUEt4MAvbf2fMJttKuL806T+zeuA44H7C2khKL0P
zs2cMW839eGvNxpAQofOTiVl//iHw6c67JV/sK7/giZy/wVfRsW92pShpu1KSjtI
iSvmZFYipn4AeFbvPG7w3/6E7tCYWafzWGHTlifV/ne++skIDMO0e9wsCoiAl0xr
2vDInEIK0RmSsfKJSPV23FT2k6Wqzw3YThXRd5yk0UVMoKRpvxPl+HxleixzaNXn
01fZZK3KgzP3T8hITGUbOXvRfwnLqhecA/WLGuxPc0Kzcd74lt3so99Ic0Qu2alr
eAfFYMZBBobE1L7qS90IKp3KHpjhfzJTCqsTnhnjJB8hCOfuFTVAPMMsKTK2mWlV
FJFsBaXPa3sIs7Hz+RS8pFcmE4Tvti1BsTWuQlljXO3UsQzHWojb8DiSw47EfykL
oTNoCSWEfWJE9wyDW/nfUi6Xum8r6QQQYMHENVmMFySXYa49YoKuKdDtDrpBcpJo
Eqoc+VgO7vvaiJFoUDQCVU3jfSxjBceS4z6PrTe3KnlLiynr25pW6zk3DWcqL6Vw
xH0KlK/ASTr44e0dlaL0N8dso8UwfjIB9iZXHcY7Mhf33oXDr4bmgoEChltI+7Hw
fwPtKmXNrDhVPIKAMrkVS6oLohMpypYajbuJS0AZBnit1TGKgFaLMnxNdoY9azvx
MKLVrdvHC/sopOr3G7FFPC2CkUxLKFqpkJnBBslgmVPAzharAC7j2BgigT0CsfUJ
B1y5O+dnHZyDFLWCjVgztDL8BQ80NGswDsXJIM2KAIrQeDNsOz7g3HvF22wLk8el
k5lGuuQkSzFeoOXJTgdsnA==
`protect END_PROTECTED
