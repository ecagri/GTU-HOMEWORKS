`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kjb/R6HYrAsVsJ7DVyg1R2AF+22XzXcukWEjo5MK27egKC+KJrzcNliDFd6CeJ3U
igOScS76ouit0JJ4Q7MzhEgc0OuwgKDHzbmbRzM5HaQMD7GnSHIzVslioKKnbCwp
vP/luB1waTz3jr8NnaoVR1e2ggzh94TuvxJxs8By8mR94pD1qHCh6QO9cvw4zOkD
v0nxzRomhrk8iG0FYheHrCaj1yLnWdjy5gidsQrLkjy/KmoMvbS+wTXT3eMk+DnM
u3AUSDrkA9ETFN4RAmr3LZGaAsO6DczODBxasY36d6EfikUqFL159VdQPCR4yGgH
nLVlNZK8vG9h1R5t52Y3lDM7CBatt9d4mVBgQcmN5WetUjvEJ+2QMaqDt43U+a+L
95FXpWHKYFHSCGm8ImZOyarZb9k2mK0lxhdWReDyKDfIklySMMD6bzrTs2ifqKSr
4OtdNMwTp3oWwoaw1+WsaNRBs1QLR9ALfpj36oaXkuJIlnaPu6CDBr/rBFHG8D3V
W6upcUeM5DlyoOo7aRVFPp/3OfkOBKtdnMmgP37Mvbc3058Uj54gaoNvRxrwEwbq
HcdxLYssO7qMsHKp/PUm5UpDpdBW38ZgPQdbmLNomyaDwqbsztpha+gqHkylXD7/
dYFJ1DuAVd93TeIULSFCZlg6ja8NrijEhHShMq+6vYP21gKI798totvtx1c9+FiX
BSWWGJGgCd/cH2eSefLGQjZ1PAEKGUkKUzZMFrutCL+E2MYXh+WJFZ1/enttVyOk
V0WMr8UrPR8ZihLo1LSoIzGz+91Jjkj0zfSbdHK+qh93sZABO1oAcQlzXCCrXs3z
e5ptjDOPJATjCdYU9sRhWXiVOs/hQRMuSL/JrsKag6Z8Z7ycxlbPXtlu67sYnA6S
/Rj4R1fS3kalbliTTrr7ZzwXOsGiXDf/+22mJoeVcExQl78yi61OH9A6oz4J/00G
OWcSH3za5hsvh354s8HfgU4ZzCm93G5FFOfHlOImW2Q=
`protect END_PROTECTED
