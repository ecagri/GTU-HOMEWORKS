`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UtSUYx7gZtJOKYZ16MtaNWOG4WT34epmK3aS/uhF28WD15QXXnyy53KZY6SQwm4o
DNH8r3kSr49WxuK3W774irB5rE8zwaZopQcBHySZsQJvhPRaKPk1CPC4qq+UMft8
0MIIZ1EEm1spXRwdCW6VuckPor48HG6nd82cDM0w8aB0KSNb7PDnrcasg1sZWrgT
IVWKup9JO4k0KnRyecegR1DvLI+JBBOeb96vWTQs6vF8BVXnYIJgnSnNit2JtfN2
WLHGxreFEYj16sovxiztuoy4FgfeYguOC7xreUZV/DwCHcquxjw7pLoPwd2XrIN7
TIv/k2MRxvmzC3hXmn5uazQxRgHaJDBCIybsLIT6ekGlxOz1S0qUAob95pa9PWhq
Pca27mXTfK9tfaWNFWQ5y2obWDQCDIJyAUW3l/JZA12m+BiOgzhjkKR+fUnzWUbz
GFFLaqq9dAvmZonCn8e1Mya5cHbE3dExK+oyIYLNR20JNjIsDzGD/lkZ8II2du7r
DT3vBIU5n9rSAZoUIWQXqxbSlEoqrQkDOw9XJSNYAWNLEEu3W6t5t9k0zaEzr12D
GvdDBVYdL8TvX7vhLbG9OhENkxM3WEVf0MXaZI1WLYPCI3pK+kw4C6axKS9BJFPs
ZSLFDcIvC/C6L5bISAqEF+7CnbOyAANco/Ri7eSxn8/BioPmMHI1ty92BuygXLA1
aNuHWg9wilyNd8/QyJoA/SNOYrlOWvx4YNbU4XHvQ9SK6pU3Ph31nve27HGrDbd/
XdYBRJu5b5ASWDaa43naCIy3yqP0/dOmlvQLe7CL87Izb68h3pC4gkzSrLszYOex
SXc3r8mtsKLU8o4SNH23JdjFKP/UJpYVGdy1DtBwYYRrNyMo/JfyRzDsG04+n2oD
7WnmeqzWutKr4BCGSKzUmHUg6XJu3azHaLiUKCe56G1Fr3I0brotrOxa2miB7ilG
87UmcEeLsoQytFIQEgGMgdEcdMKksaQ9uTPdd23qr/OvgtxlloyVp6+s2CexCsqn
S2pxpkMlHaKIYNUxbwuxFMeI0Y1y+Ut3Bc6eBy3He2D6c3K71AKpqwcobxgN0U6M
eOrmnQkhdqgyPmN85X5cX/7+hvh0bkOWiz5/9JmxQGlWs++hAjuj7vG/qkpn+Iaj
rVDigw888QRxmcLy1mldsA9MlS1aWVQR7JphBTT5oGuhLC7r4/abYEEWvkfGpWAS
DEAAv+xdJvr/+f+OPdOieGzS3InH+WXByN8pGECN+sI=
`protect END_PROTECTED
