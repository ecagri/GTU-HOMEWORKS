`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AZQuisYSCTDQ5iN4x8abfy8wuUEj1j3yM9LDgu6ecu2rBB0HsVlFFb6q3w7bQ8nc
jnkQ4KtOhTThNy4Kk+cStHHC3CvBAsr89M9B2FTBViDSZPqMkrhfVf2ZYp/Gkfyk
15YX4+OnoI1kWnWkbjkp5bBURz7h4Bsqk0AWwW/k12+Xs5+JbHhW00dSJL0YK6R/
sX2bj4TMBTKITOXFGCbY/XnO1/LV0BadmBK6J5s4HP0zUzT8atL6ER8Bh7A9Gjx2
bHKNBEiqX3j41oEeSK8Vqzu+xwZzZsOKxf0dU7kuvP8t3dK3uwxSon00Ys7TlQXv
kT004paghIicIBLz0x8GGn9Rfp48DKzJxgm3MeodOqp1UuVukbvDbn7PZW/iC0AF
/2yMOsbeyryOHw23woMbDRJ7zvnfb0ls3Uk8OPP+N9NZfMLxMBOBTarCcVTmkn8W
53OezN6F+n8yw5VuUS/EXl+Butopb/XaZkVycuTOqsSy7T8KTYyqPb0TzJIyjQUL
T5LTEiEVEmKjA1QgPdWP/Lkp1cL26GhT+u7iTOyDH0JzhtO+jAcbXxwPI6EmK2rK
h/SZSYejjEwUQaDIIwG28dHtkcD1YTl5xKSlBY2RkFCSe6791/T7JfScdmgxHUqS
YDZkJq8vAw2YnWe4pqvebAJg2YkWlLiAN//yVztETNvf4bVThN5gUiH2dIHQ4Tiv
Nj8SaWeqDvkc0ncZZgrfP47S/FU0e6ZqIG91zJm2S7hbY2DQ4Azs3t6d4YQpp1ls
L5J0107HW6/rFzJcT/6dQbrI4DWlpIaL54tqCKqcvLjKXV2rxHygoPzhrOgz0Qir
4EHxJ6pZuF0RqsEyCaU4F6T9MGNTrYEpTGLdoe2njjxPB/wQwQO90oeaShlknVRN
QiIYxa4sBAw5f1+uo5oSutKT9bVp2+yn0BEp3k8wCNOgYAamVzMpO8hk1Rz+oy0K
n8PXkqXTntTwZT7tErFgEVVenzL3ywyCEiMnJ4IY0Iag6YawXSSMoTXmOy7dsQLB
do7KFlyf8WrQa0F42XiHLMfYty/LQzHNQitWQ0mqCPGQvfRlaMtEusRJgDJEvtUj
rmDUQ1HCKED7fVIHEVgMNh0GXbdY71+7Qeyn4eaXL/dKdrKkhBazekW7ciT98CJ7
7Hmc8fpaXQau/+G05OjgZ0Dl6PaQmBIAvnDsq5p66DFcz2YqKj1mO+gR2qAe1M6t
7KzzVd0PfH+A4Tcfk02T9BoPUnF3eKdu71mv4oFNTuPH00f8AL5RDiMuQOhvKFqN
bKkmc9e9SnBcwjsl3RoJjeWVDd6OEHENSTtUNmm8IN19N1njbrtIAPY6wzeaheyE
9oFTtLKuhDP6xyQNuzEYsbRP7hyNpgTNZrA0iN8jJDIcS9v3DYAJPvb4argfgLwH
Z+NHa0YXq1j19RVdGKpb0xTV/MCYBdd0qwvySxGVCxCmEM4VerTlDDiRFsde68zh
x+XyWVwUhIdiuO4Yr08KD5YKbIjDD67YUnXIM0p482mPtIYztBiqOEqA7Ogxi8D9
rsh4oKDL5OTNw3aNqi287+IgfNn3IcRmY+rxaz/gSnR1w1Su68dfydyLPMQUsbm8
kqRvKlurpl68hl/v8tYQCtjJjPTP58qb1hx4ni+K50dl+RWj4Glxt9ND0+pVkh8R
cYl0Gavptcf12s/DtNjnJenld+sIS1BMI6GWMEhKMURb9HOUrFj5ACMuw7gQqX7v
fob4uWK/MtDFzExiGSJFv9bLSK/fFAeia3LTEUWZL5I5JQDnYGGNo2V/+KqBMrKJ
wmAtSf1VP8VV0O9IV7NvPu26ndwUHgtAyJhLRMLPGuzKr4eUZCDcYhBAZP87r/Z2
FFra8+Ky+J3vkRNslS6tJKncDVYsLjuBasdfbs85wcJutM3zUYu3dtH3NLuuX6La
OTySuGLDAz8HEH1PI8atoxrMDZae9zHmp0T2AVa+WR44V0MWEwk78G/7aZJAa0zX
H5DLLdrlSMGiPis+hxoSl63VWGvplugvqG7ezT6w02FVYuviLrdRPZCRpV12/upI
1qdtsYkFhhlsPKig3hG9gav9gqsSxCcF7bqwCeGpcBBZOgE4OJcf/xD89q0eSKbA
6y38RFKPAR2engkM6VVsXMsj56sG4wwJQv0PFsxYmEHqxZTfmCcIwzxx/iZJeLiP
daYTz6Auz9qNdtdP9Z+uWUC6JQGsRAYoHO8HR9Y6APQvtVQdHZanSTIbA2J5sNv2
6U5kuFpI4uAN4RhpF31Xnl3ejv/8ga2Md0pUiJEG3gd0XhmABlWkv2wMa32SsTjL
5Bs4fqOM0jFRlFn7sY7NYT41UHLiLaC/1GDSA0eREMeBve5okFjiVTqqwA2MdB8q
K9AAlgcXKQ2j/11R8U4gHwXSPXDQnYtrfJ2BSH4mnUar+cYCEBHC7gCWJIh13XUL
nmHbiqJ6aje/l88DZzLqLeWJDfVWkhKWu0XR8MSKcEGqj7bMyqHerxM9wL1YXjH/
Gbnt38YuINbhcOLOcnEWvNpI+l7OBe35glzqvWypwy7F87REEy74WPJwu7+NGt4h
Ohc92LngP4dBUGcqpS0Wk07k9xxuyk2uiK94z8Xd5nX8oQH6iX7hHRn7YfaY830s
86/Jl9X0JSUfeT9aBkHE4nh0mMexWhgYW7x6CDI2nGxDZLHjHOYtZ3gnbIeJ03AU
Chj1y+oVySzPfv4VPw0XKPIhaDGyR3998bN8t12P3KXLs/syYUxGf0EIdIF2OcwE
XxGWdwal5IC3wAXL88JlXzdt5ueBR4185ctpuy7yuX6qjxf4qDt1GRXvdVMbMkqD
u4ZqFeM2UfdYEbqNsz9mQfs5Abu/Qr92rIzEO0tn1x1y/lYyNYsVa0WJy16rP4O8
AXwmhBz/y+5NTH9yAUd5VW0rLNpFcRPAbmSyd+W7DmEY4IHh3HfxZNPpkq3/dLAA
28r0EV+uSPO+uCyiBRuwWveZ+cSCC/JqHiPaW44DiMksy7I0IciQ5FnE2CwJSU9J
a88hLX3RiVXXI3FhNW2sUsdaxvA+YItvAaJG0w84/Ew=
`protect END_PROTECTED
