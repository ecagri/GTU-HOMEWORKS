`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G2Uz/FjiREMrKXlNUnE1TjiLHDcgEF5DPikVZkBRld35wGe1AnmkL+lKldKr0FFq
rsb56i5TtoNaHLATFqyebXf4inO1XmzJ2ZqOX9ihH5ktJ3JMhSftXP3iTv+lJrJp
ARk+tLGUFIOQnUDTYeKasbOqLHQfrUJEW5g0WmUCpRQ3k3DMH/gaxuYuhkc2M6l+
uv91/VCZwraIkHyeWSa8+P3wAlFoukzge+Hpcb2hw2uq0+Z3xYBEzTOeGy29S2Cv
eKCulN7l1KJRmNuJn6V7GAJ7r+eki6cHTg7eYPWCSYxTKhSumGtzuLn291+tBenS
dNb84yVa7aUhhBQ6yn2Yb4+OJ+Orz4st5z+f4ceU8gvKoYLW7pMRMKQ0h5l4joBl
TDLwWbiS1ALaXaw8HCM8Wz8F/+nBU6TJN6OD7RC23R2fOIeN2dzOj9exw2wuXP1y
wQb6r3tD0VN1MQIdRt2g4Tikrn7P2UXfArWzwAyIfORESkSGHANDOp++XxOq43oT
RZk00Bjl1Bgxr4Xv6XbuDB+P66P6HbUISS2ee/K8skvc5RpL3mqu6o5dJv8keyzm
gab2dXfPxTAwS+tBdQLf1go1u1NCiZbI3tSInjiUt1NOFurEZmUMtgmj2jLxpm4C
NsKENXIBiAJJsZzTaOTRX39bRgsvym5cKemsbeHvxTWsOHuZOhko18Wgww9KrGyb
8P+EV0RIywzkWPubab3Wy6XQa2N66dS4Da8Etphr+laxgiVph+OulnEjLA5Yb+57
au+qsbVAMZluNaV9m2eaLOxRlnJZsYlEQLjbd2sNru1JknrccPLIa1B9TJR833Q9
YqDsFocc03V432PzPmXKbJI2hefyodxImtYbCNhmaGB4kqaFBj7kCxf8DxU9DODA
tfSu9vVfsByZvwD58mxttuV7Sz9AnuFMeJBJJ9CwjJNdx/D8M55cgSvlSgC6AMue
RhUbFQxntpeEyL9RkvAf/9m9T1fcU4Y8+cjduaV/XOB0q8oLlTo4wgi7La81OBn8
n9r9CI8SEXcvh+JZJ0dgbiroLQyukjqH1ShVwEK1uGFAO4hTkbb90/u+X38rUAei
nYTpH0PnYdYKMrat+RobkzTIJ5N9zxSyfwbuxbYYvVU8YhxQalyWQwJMBO5I9yWJ
wcaJVQg12fKmehYpa46/Vq+LiBBZKAWq7Q0YcXOHg5nB9kyQk81NcXK9/eApNtRP
iyMo4h6jDrA/OK59JoKFbJxWiO4fdD2kMtBQoBULxtZv1qNFXJ1kCsVej4nDJREF
T8Kg8P/l86ODuLVuLWiDENpvpeDITI6QUQqmon6s7hxKudNo55ygRUvz4h2kVtml
FbEvDerhAoP2mLY4XXvFeoXoq08HAf7wj+A/F2YWjWsGcRDo18KO4RGc1CM6FvOo
fxu6hZ2LrXRmSS+5pLNRuXvwFwM3oIANx99bhpCGTx9F7tn9NC1Jo8u2hcALKGZH
rADD/TjGr2Q2ttUxcf0th+0OPXcITLwqmVO4b295BKy6DsNklhXmuo56qIsMIEm9
Pw1uxGXHhIS+11OzMGDjJjq1ZwK3NcDG9mqauiN0cqZBT78aBvLF7EHTEVZ0K3qz
NylQJ+4OVJsna3fKbCneyjAa+Io0fKnCh7JuYWNp3vpj/X74y0shWA/bLNy90Kt2
ElYQHNqgGe+ve840h1xle677CFJOgCeQZQQi6eUstVtF11GfX8SpHCB1wsfwSiM1
1wuYqKPuvfFepNIj2qdkJNkKFDJh5eXxRRwYdtkoKuuLgMK+8C0RFdrdUF1XDn7R
JSFTZaSWmR3kIwh8hsJ1PPRk/XXQiwd6p87KtHheGAq0Y6JUByszg97pbucFD/Z0
4VMsu4UbCIPiTYhWcsfjJnN1SDass0HkI7XFjXvMrsFtmg5NnuH5LrOuzNf/RaTq
BFUU0inFlUdst4xleRgWUN0vOG3U9XlzR2/Q3AOoefCYGPVBXjg+yeMpuGPsHi3b
XFsVRLxbdhfODukdcq26F0Atqy4bnN0kWxhb02rT1k/e138n2BXiLrc+Bh9SO/d+
vpuIKjGRSsn+4LuRThIpFAc4ud7M0MYVRDiGV3pp1S4VMxbYMJ+bGwRcyyScOr0Y
tKiBWxfg360l1ylitMtNeE3igTvs0/SM5fBWjJicCNq0V9HIo2iyZyBcnWRjpwt8
KVklalzYPYWV7BQo4MI+Wj7D6m1VkB81RQBxM6VFDuSSKgnrXHOKo+yPNcZoRek6
/alFN74k3odkbKBLN4v0NXLNDFsFZVWmRLd2nbUsDxM2yEuhyjKIlIHXVNQ0qlsY
+tjddm7V+VUde6p1voJuahNohGM+kv4aJjJqLAhAfthDpAKIX+KyTczw5P65Rd2C
shZumc/8ZGvJrRYJ5OEalaLoXJiYADu7oV9Xb0Kw6+Mt6GI5P4YiPXjrRs9xQm+0
s7q7zxk2FxrkCuLznvN17zOfBvFgD03vnGpNVQv0TPACqXml0zn1cVCYcI90V50v
Rc04+7cvulKsTTLaF8DjCWngfxVPwEUxqK9wtAmex3mW8u8kPFjCnvAQVYiyMQeR
gST68TMgTIF6aKfn4UJ2OcgqQuEJVPPuGB3LcQxgxOIaCaoEHA9KiVC9VHyqVxHg
K/BiBxqqVwBnRHpogqGpa09Mk7PKUO1w36R6y4pB4pGOH7M8tZt458krrcsfJwc0
PZzNXjqp7sDWFNX4mqtxp6okS5ACQKvj4BhU2uP/pk+pulx0E112li0JSEu+aIXB
fZYdsqUCeL3/Orzd80B4pddfJmP60jIyNI5yXZqh01/MR+rxdWZC9HDAhdty/fTZ
`protect END_PROTECTED
