`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
38FiiTMIgPQdbIEOv+syUvm7h1/A+qmdoSsVe04V1oBW4qf7ZXWZAEgWskdXKPDD
eVjGLxJoNTNlgtpW4+JuzuV9WsBYE/nPtS5oXcbQ8p8ajPetcRA/QFSXOOhZ1gux
mFS2PQ1ZI02V5T8A3Iy4VJYrv2qOgChE7xynvjivPK+27/AabZN+iTP6zIT2hSYr
zkkxps+Gj0XbvCYUXnhlzbKwcOEXuySPbB9Ji3IAT2doOuovZi1Co/RIE9oreCPn
tK2M1jGN6ZTm1mCyZ5SkAatxGpVG7Ij2Vw5KMxo0kik0Rd6ISKXuMepXVr0Gnp6k
/aA5ME76i4Ll1Q8tDnIa5Pqsfz9SKPua9G/ccKz75OFTCc10H6DeSJBKAn2CM9qq
2wS+fm41TFju7Ali6169cMNPjU75Xl5yD+QDFJh1HMZgiE0T2cCGZeGglgwF7Jfm
fdXLazSquErBcHn7o4Q3+4YXNNBbnfAWx/bY1Ix5o494uTYoT733vLTGvu0ifJ3I
KOH+RWAoiAvOkWOQPi6C9c06+2OCl7GjzW1cFBb/Y1z41ma9vYDc1neCXCuicRQi
D7kotTG/qfVCR0WLDZIP++sNZP0EMLlSxnZ7tVMPNCMRRMLUb2GVxkNrw9pPkUXv
KQ0WNedX3kUfEtD1H+x1ywwLhDfUt6nmbsrMMUzfaiRL20ZmQkr+Cxa0ZWIm0lpx
xuA0IHYQ3+8aXAZFDXM4xvYXsAZjQJQuir25TkrsGleTchqRZWoqkJCYZy2sRe0A
cobZNdVoSaSRQtmO3NYg7VoYZpNsZZGMDJm6EP4SRAKKoRFSt5LQPVFXuC8De2mY
NuaZkLAyroYCu3TaLQ9zI0n35xbBXrzToiTYQK4556hnOva+rAgJZM4BmEPvg/oM
0HlesN8pr/PEAroJe2TOWoQszILx7uB9mMWar4U8U32PJZhR1ax9YSUPkjh79Arl
w+yKHEEj5DVcyaQtL8eBNPBbW3ycMZZagpv0Ya2RXcMbH9UDC8g4eh+PpQIZcCjf
/O0wJ7kPj0AjfSyUW6u93ZMzuJ+QkcEZTljxkmXRSQV380fR+VnTpSVWvsHQZG44
8uaL+VPY6qdW+UyS2x1I5rcljW0arumCPZD9mCB3JCVENrYtFy18V1w4tlziyELD
xEJMjVvTnZ62YTXauaLBuzabIThWePceWLjOj6XXs5Xe+9Lk3TE53rM0Zb0pN3bd
/XroYIYJwAtSt1fuZJ/fICIGfskA+RsmTuu5qKZo1hLF+ZCbC6OMWdAdIUxjTK6M
EMxyjYKVFtO76I3hZdTJ+gJlvGLgwnMQ23d9EirC8Jb3ko8zoctNof0sNyCkxmyc
`protect END_PROTECTED
