`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MqpLKMxGfii7Rb1lCmFQ2JhnLPbSI4sGTRKoRPJ2jJgk+esG2dwQ1o5HZ6Q9iM35
dlBWC3fHPOT99Ar4Z4R37g/FbTewaV8C4vAYMatHg58rnGGZhkhodfJ5n8rDUF81
zlirn6MirYu5YchNF5z/8aEnDSCf/J+DnPej0/DwAVVpyv6OmRZ9R0uZYXGqwt55
j39KgwPxQ2xeflnOYCOVEMJnfUmRVbojLxbnfenwB/Nyjxi2jl9UHO+g+IYH0f2Y
Vax27S5D+eGmblFCHR+whW/136Rmt6fERwzBdkuZNxzijOmiC5VzcdyAZsvu3A0Y
IJtWN6bRKUL+Wn5TDXWSYj7gWOSlSbaswkN4hajlzz4Pb7COjcvtS6TqOjgyEYVL
LYMxGS4mZK+bd3R/lbEKWFUBJ8/w9Z6q8wlmEGHAy6mZeTBPATLmehfo5S0Z9mmP
89GV0XCoKgSGx8v02lk9mYpT+tDsz49QJ/LoFbpnxlI23IxxNuFd1D5H8+xJKlk7
kzQYl+1ilOGXPE0tLXW8K4udDAuqy93JsnQUL9WrsJnt8FWS6LzKVZ3IKn11t3H1
1KzTLXP4ZJG87TvBvJ9CZfURPmSQeJgDTBAPtcHfc3PQIF3MGEH1ijsUfOkD7SHY
xPwP/PDv9VM8/q3ssQ5s1G8B7oaNZBeI4/WCw2/VHzhg2qttzudS6+4hyx252ksb
tEeBPst6Iy0ztYMHuJ39WWsmV27mwhXKCc5HS29v5/NpOCn9Wa4DZY6wd+J3wQ5q
aaXw9FqAXPqEeWYd/KevVevL8BZgQG4jITMJo53GU7y+6TfVdKJiLVjEEQS+rBV8
LXT2ZzsA5ue7LaHxDGXJ4LMxdduUpzsrQ4+yb+w7LPqBTHMMjjvhiX/wbM8TuPnT
7hVHXpLMXa9rs4Ktf0yJxup40tIfAqY9kJ65HwIkg7ulgwofXsEWRJxwjlHMlkw6
wJu1hnYhPHiORHuH6OUAkmKqinzB58qlDSktw7WejKQMzPIBWF55+LtscB21Hh7j
EK/9vMY027/yVF7zEEM4SsjYdf3ie7m0W25Amr8Y28RHlNo+yb3R6M5FMeEuP+ye
Om+308C23qpgfuQLJN8Tg9zBtuctp2w1A7cITXV1IMlufoKVafi7DM6KMr5/1n6q
AwYe/ELzj/CtldKyCa0y2rfTRpHdvvwndJYYmfGSp5otVp1BSGJhTG2CGdFoftku
ba3DOzfgTUmt5vMzkB1TXBD+oC8B9CGL8yfQwrqswCOhpWGBoQVtnPluEwPRWlj6
nCUIoGonl95cPMKuNCUCSggYWifzQsWvCGdPMUHiRgQH0oyBKJoHXeFTQVz6YhS1
tToak+Q2V821oQWNN/uTjxLwgE2Ff2dhLem6w0hQ50rxOfCmC57E7U1Yj6p20KRq
FCcJd1thX9fSLV6lCKRAv0PoVdoVX4YidK5i6Qr/HAVqkBczIdpad1aZBBWjPtVy
aSfui/X9uLhwAffXdBINXDuKn+sYdQGH92xainCPGRYdy3ZlJEI3KlYkaEZDzVwf
y3An079rVywDmLWU5aNz62ZeQkSc+mLyk2aW+S6nsTuw4WDjiz75/VIH/hQ47cPZ
/Cen/TfZg2AsyDnYN/YWjtDDf8sb+7OC6kOn2R5NXLozf8cU8klBsUTrA3hirpaK
J3veQJl3HLxVVvE1s1CAq14h+z5WFkP1E4WjBzhL+bqj9yp/laXZPcZ5m6Ooa0l9
hWE9ZzAteuZo1HMEpKD8VrMQJrE5kZZxnCnEWEA98YWLl7w1mMR4DIRV3kvdoOcE
snkeOpHbJnW16eixcE/LIEDHn+7FwbSUQiMWL6YUqTo4kU0SHq1Xh1Irra3NNf27
4DoHzErkJdRvXR7xBPeHIAe1koXxAIFh248GUq55eaMksQpajL4XjvYS2MseeWu0
nncHFP8Yo0Wt/FZZ5X+b4jpmDsGvMIJHA+qcM8BvYPmnQqwknZaJ6t2rP+cEuLHY
5mAYFyb0a1d06SAj6pVzgvy092A0NHfWRFjQ41f8KRs4Q5c0VhXrJgKDK8XM1YK8
fFVyNurSdCXQPpU18vbwxUhsjfNJuYeaugwZjHiKEn9LF71Ufe5Bt6ov6s03x4zt
vdudlYopqNygykEAbrIO+UP4uy6zfLmSGPj0DeRV50SxceLiCdFT2tTevwbgR0A1
AgJhU0x5GW8xHvH3HZG08rqfM5sjUOIOSFkCUevw34anrfPpXI0/i/sBTWWqRYjk
cWp6UGn2GA/taurGbZJAXJTJrk7gQI1tOx529LO6XcCGr6AN694cVSakeOKn3cxA
z8t/rmhL/3yzQSPX2EAM4owxZFHjEabTldgCo6s68UrTn8Rq5LLj2MOuzo5Nap8b
8KcDkGfsjFVwq4dPR5a/b58U7DuJipR5iO8n63QZfVOvKCbYlvew9ewNgvVN9QM9
aT8qNiX0cLc5+CG2sq6IA+S5R01Mdn6zG5ylu1sACH4ZF+vchYSRKaaePDuBMoZU
3MFpDo6/P73XRpGu7ilaHOcvvYfTUTQrE/1gf9adkRIW2CBJoqySAvklgOQHz/2y
TsnAt+wOc9rxfXDOF3T2Rw9yL5MzluX/Usp1Yf4IHHRssmi8WHTRarqMA1fQDS3V
juhXw1kdc7OavqQTZgl/kV+pNwdMn1pQVVWaeKz4IADq5MUDoJQCGKeq5gAfftDz
EiXJ0dX1VS1g4QLCel7LxHaesYeTLOatKBH/w6kT97MWpcRZcus8VWZbJs32Qx+4
0ldYmPtK5wkEfatSFgTcUTtdGs32qPPfJbCORopo6DJcr/YixcSUXh9MfnpTvS1N
dtBEt1gjAVnlufzsoDd7FvwByp0cLDaLq92rc28cnzssw7G1ylg6f+4E4IzT4cey
Ki8Afx/og+Az9fFvwKZNLvmWHT3uI//PHXk0lb6AlkjQK7OTVDri+OZoK/S1YJKJ
kIGaKx5Tm71EnaU8Ulr9+A==
`protect END_PROTECTED
