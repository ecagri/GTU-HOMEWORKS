`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TtYBBqRrEqzIgNXb3mSA9h2wstxZsLqR6oBheFaPI8hKs1yc/xk2QXuPMc/VLRND
9BFD9LZ8BkvnABMlOg9kOMlB1u92+7YwR88jlan/UgtIfRpQFbKDzlgqpRA0JDMO
YRQWlvHynyCNV8530paE/2mZ/7tJsgryOuqdBaPLBZKqcsAQm4buB3IfkPhccH7l
//DowQZERjlzODx7zxn+u5IFDitirJPKnBT7UI7G5XNpfGW/xec0CkqiKq9E/LC+
sCbBq/4KXPMfD48JXQDAXMlkVvE5jesBYDOCNNCEGb/K75/N1chSpgiQK2mt5EIm
qE/6sjltkkxkQ9pPjJINBpyGHWW6oq/LoMfNT9eusKCv1czGqWYhb5qzra8PNl/2
tgz6QkWGjoGAL+zhpmgPlQPnIdC/SmaNhfbuaJmaImGPjO3aJ3Pds+1zwhkPFVAI
2t8XkFLWnDkMW/iUyg5rd9EaeePD2M3YPqfOxmZYTQGmVNklUw20PC0K8oEO8721
wW7vJPj6MSvOqFALQpYef3wlZwFZ+/kQCih/Dqf1cVy246wMzOgF2A9rdbL8x5pL
wcL6pUhzHNqF2sHRrNh2PMyLtQ0G8+Vz7VW7PrUwWERT9onXZA7rxjuqhOWEEGZe
JcGkGnnNOl0oE87m10MZM0Ur5CPfQnfQPNiF9Y9HWrtTfWoEv7LHm5Gs0ar5mo/Y
V0R7XgaVzMLjWV9MtU8eSLjup5k/rLspXYnFlZS42itSOnHeUQ2Gs/xduvUVM+iQ
MY85bYg0dxyxRnbFHRWj7s7ejBrbYO6mhFpsR2Wb4YTeUqB78hIEC2M2lUXB6VHQ
uj8d3xEQbJLwlUSCgUOXofjHZ4+51WlJdhY412FLToJbngyPxh9ZWyclEzupdZPw
QrKTzDdaBVaiqyKvIO+Ste5MUCIqX1LfA/lqrCd5FtlK5pNYymEG5oL+GkMkMPvF
K4bKSfeEfC08esgIPa4jaM2K9W7IlY53JCl9vXBk/gBgHqiQUSKSbOF9jXd5znGD
MPI7VGog+w3Jk9o+WzM9HkVJqAm6kCy5SGSITo0q8iS59mAu/Th8Kjj9NDNBn/EZ
CF8GGst6yodFhyKnPTII6KnQlz848Fl1DNCIOgZfl+5gp3BHrJzFqxEhoYWJCHEQ
3dJz4K17aNW8ZUKvYg10jmBAgRsJ4YdcHb80tJG3xF7qmMWJYfSGMZmmKueqDN/d
hg+ZgVf6cDlMlty+OYnt55v1hz5eTEL6O0Fjc4P+Feu21wkk7WxmlvJVVex6DwuP
v6C6iDY7BgFR58CpN+nXUlAC7nHdV3NTuHmWBrEg+DsfsG94vsJMxThgL+/GN1+1
tFXHNlZHRFN02Pmb7FqgZ0G3QPKSYBvVbr6NUz61gwwGpnufN/RUA09oiyV6t0X2
omOBdmGAKacRSko3jgUlgyx+jCylp567u/w+K8MN+UUatJ/jR7b+iKFsxdFhy0Xg
JtTxZgL5m0CgUXu5xJDuzzqKXo3uN6OVY4Dgmw3vpBykRcFr0CuibsvvlEqIVuLs
mWdmtk4J+JcXhQ5ISE3t6ep9rLGqa+cFHSjszGqAU7xs8DkYM7hNHC0ysQcWAFda
WBSdVg6UHR9dxgzTvOs5K3FVSFcWny/XxPXELIgj628=
`protect END_PROTECTED
