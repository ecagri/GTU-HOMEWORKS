`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
48EqtHHPSp0UxjEUhCUabRHN8jSxRtTy0zX7rl68GR+edu9T+2lWoKJw/Rl+OXiG
tmOHludFh3bkZ7XBrHD6H53MWPUSe9RAPn0V64FiK1Yo5GsABfg4vGRaLdcLLg/O
lyyXB+UsE5UAsyd4n3ZoBDjra9rfezmcalnhRKU8MWBxKhGeAtSY1yK20jZNK8DI
TvfLDAn3bapHVPEEM1jXB7x8YJKm1O42LAMX19N8pRkrdxsKuUaXIAmrm2cqi9UY
vXGufpEPX/TmdxB54tselYhXtku3dhjO/RAOvfuG1Fs7BSfn6RFM0tdjxlsm3PuY
da+4oQMhYMWy0S2tqP01MiFg/r+hNT7QxNxYbcHbuXGz2hhJ4d8+3Mq7uYCqt93e
xPWpuHdMlslgDmOPjq/KJT2p/QCmoNv0Tpgj//tuGRBR8NIlguGUL+qciOn4ICRO
oWNsTj3PenTHHt7vdOuZ7/tWsei3r62pgY2islirRrF+BMTwK8IX+P6f+TEfvQzk
siBb6xYqU3unsYZ8ruZfl6CPlHGeeVzwdSrwr6Figc3RSP6Dixu+f0etGBC71htr
qA0130WGrDQAQbPjvaJtc5xeFqxNjGRP/sKC9XM+6MErKnzwVonwzAzlzOBMJt24
FET63j3HRlcTH8IbCpa3n8NeaJ6g/nogRfEP1bQwweE3RB6cAvMZ6i0RFh60h4dv
gxs5Ri8j6+QPrOl5xoqi6vjnHbskXnW02AjW6YKb59sd/dyLc6/YXVUUhxiOS8P8
Af0LARd/3CS7yMtrNVRLzybs4vs+UDuvp1fDxqX/oIX6Pt/wbq67IIjJIAspU8Xy
FG4HEA78yRGl6XYsG0oXNEydQtO+LpqHKWIlRvDZkaTvUlOc8sNsJMhk8xTMhb3a
jLtcjQJkGjXzATEDi/5zjkz5B1xx8kK+vl12tIQlwQIuwJgd8mIYpi4GZTqQytKt
nKV9bBe55kFSaegA3DB2sOvONT7QC1fAKpSEOunhhWtQE2W+rrjCpkogaLeu2q7+
lkb1sk3aaVd5C6cm1Hcoj8x4RRyN49Yo28ugocyJ9BwvbuzNyx9r29+iS15XPKW9
4kbyjABy52s4Xqm4FVpODsJ68YQWzhBgPi49MBPOi93GKgMLY50heiywSMWzM8Ex
70qdtqlAY/VbBHBvAhryi1SV0ez0J00VED7pJkYtr3Sn7MH669cx+kQP2s/aXV05
7GR/OEhlStKdA9rfppnSm2vN0i9tBoPlLx1kgVRMMIyiEfQUH6F1+njBRX2QU86X
euaD0CJ9TiERSksUf02fkzgVMP+PTLIBu0DYgEJREtwB+7ofXfJoW9Mc+ge+ZlB0
7qby4sil0cxLNGv7MlQlrg6CaKyEn3kWL9llYrTwhT1z138AdkB3dApTmGDMMij4
6zRYzIz1z5IWw6ERumXtnj0reOzNRVfVeWI4H2/MQLQgSLqsEOBul12lNdgayRLa
`protect END_PROTECTED
