`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MMXOed7dlJi1XlvPE96rUCmGAl4JDhKvBFt4aGhHUylhBn0pRCnWHiFp8vW53cFg
QDXTPDP/yxDOhotTPQlBu7OvXyIPqpVJBhHV5+9NtMSMuSjMJTRrEqZbkoM64J3p
awJHGJ4x/ByL/BdsBRsM/qZL42+/lXowzkiCk4HIOgY10VL9IAeA/20QLWpjkUgJ
mOYpVD2FuDPO71HAbHuw1DHu3yoHy9wD6Amv0ZpplTaDKYRg16u11hvzPy/pGkCG
Sobxy+pmEQrs5L1/t07t5qh117YhgTfNthZjlfAYsFcwlK1RExOVOueGt9HeuiTx
ntdhYK4V0wwTvjwrouvnazKJLhOhFM1g5OPWrUQf2AErqqMAXiGTR//tZpwmiAx5
kt4Ds9tHSb+2KD2eJGDu9v3gF/q86fForly99e27jfYe9xEaleZ+cDXEt5Gj/03E
tjwy5NeByIgWVZVOeE5/myWnWZPjDVJ8ROeAz9AQEjNBCSGB5fQzSpi9X3hnIGpw
MPMuA1BxcVrseEKS2340nvNlQ5ftcvWQOV1plN3yrRyXJFFa9WdnxkRIGMD1ydSG
9OUb2uiVsE6hlG9X7vFg8/1wiKa7FZGMCXM+YQK6uq9dJDOA1x9p3R02ThRHXhsq
ON7+CUOFTObqRDRCOxE3YPL1jqfGnWMXRlkdsthanbNvojsS12j0Mu9gchHvhlJW
YeLlrhKk604P89JMlpTd3u8smbC2w76jaRSIxSdrZaF02QhY6SzbQC48sZO5vmhx
5QSIIh2gwiV3B6Rr9wnTMjt3kuNyDWLv6r6uM9BcNzOgxSRPNcHFbPGt8jcDVEcG
3gfErm9VMPf532IqtJzemmkcp+QUubKeezr73OqJMZ3v2QQYkU2gtCOdJZOpKG9k
0wt3S6/8AOvvIMtDnhUwn+JtU+OlSzNY9D/OqiGG/3JTDaB6uVQnsRAJj9hCx9Zn
4R/ruqawS3AHY0jfJGZLoKMvov3ldq6WpwJ8GNdquEzmtBakH5jsXiclhO5VQuwS
IkX3pHq6W1gtMC7SvJmkr5YIhuVudlUdgYnat3lYtua7Z/0OmLEZgpTKGWFuvsWa
XPK/zp9flitRFvDvki/fMo+z8gZVVndhTgmaa5UMnr5foEdfwVCG9nEV1+GtC9Nc
PEHkkazoUNhXclopduzdRC0IV81t4McvH0g04kScUuClO99gn7af339NW1pw7cMb
XsFJCPbm7bnmjl29zaekRv7+lMTVXMzC1gZIJbe6vURdok7bIU2C2Xvb1sr4bQJT
kAcJAColvWN8YsI1VjivLFnFg2Olh3cHC0/fkoppL2SBddnRBiFNvXpxbnmGD4bG
8Q6q+ozs43ffC6v0Q+NNfqIFZ7wxN/eG3zKwhLIDY1cdD6hMqInx0SJkZbozNbFL
oOlygxWAo1YcpwpUttxRZ0tzFIz4BpnOOf7yIC6RRQ4RL8sarHe25PmvE3AwZEtv
rEy60YYJDee3AfEFup9wqyj4JBsm9BazkRso81TkoBxnFH8otPbDfEU4z6/qCBOU
NQzN3eZOhpeqcX4EYX+PkCpM9sQCn9mfiBhP3mlwcsHcdmmDUgw9s03EoFt8+0bF
xnOJWhXXjCOiMvO9EW9qlXkDL8FkdlIjY9OvxPxJpfkCh0HeY4NTJrpyCTkv4+o6
SFYmq1VOgHY6boXSIrlrCMfTTcohQSwd5zjWHpXKyU1cHh/iU2s0jiR10UBZQ3OV
NT/64JOCfCJoXJX2qhqyS/5hxHka5LGva3YpsVqZ3iusM69RJX+dGJ5EopVX4LGF
lZHF6U80oya86q2emVYplv71RbotOGVqsDffA4zRlpqYVT+WllO8fyC0LwKKpBie
APw9ezTt+KBruAs18xOFG7PfxyHB2OJLm7yK8fgAjc+ior10JJ3AtZSTRjbZOyNS
w9/RGT9HYczdwNe2TuuJBznarvR02FjSvt0t0HVtQvQpITG04iROzvCVMB8a7rlV
Rqv5qJt958j/wIpS/JG777gidXi1p9LfP6kkDOZCfHDwQXy076mKl1vEA4/S4zIP
fx2HqMe64Z2QsXrVtv2J/wnj7wDsNS3rl1btsCD43HWgSBtZ91QQXOuXbWBZgpyp
lqmHfeGeRwE12IGI5DPRlfelXj/bWwSVnox9ZogVC+3SpyECQ0yjS5sgaEZNN4ui
Ah3IF86Saz+XsQC2tXj1Fq3OaLkhydKJNGNI9ocvd55xqQLBywBq1VyRcc8Xi8LB
flwWVxFieOqgay2zs31/a6wz25IepR0Q+vuy/YHgwB1IoPBPaTniGizwYGxE42QF
sQWyB1ulKtDkXH/oSdgP7fcSSX1sGChM10Etu+WRtK9m55i4TrAShW7Um9PWSJAi
sja+rVATW6tT+VxHy/FSaS340hpX6XsqB9/X0Wg045hQB9TKo4aWRsyP8yswxLW4
5GsbrFyElGkTUwfR33LrVDVKqX4KqE+y8G28cpWyYF9lpAKzp0zO94Z0VvvK7t6o
DwXoQZ/Mma1/AsjmdegfonTDWJeMbI8sFFX+R2bsZprQ7OMmM9dq0QmTicUB3ppi
30MrG1KETH6E9AmNQg16XYtt2T50QIu/PGRef5ZGtgbRcpDPz/O0P8z+O2Hz97MZ
pCo2nhlChq884M5cALNdpY+U87B1PfQ2OktGXEsRCQXTu05xgFDAqxRApRpvqyKa
7YfWSL2VdSY4elKET/f8j5sNgq/85w/MCBppYfe1fKjMGTavvJOU9GO53Bx6EkLJ
5sQGr5WTC/IVeG1bjYXtERG4IaSmX+UcRHXlv221OSsO/YLMoO4vdwYky05KdwUD
+Uv/9D7D0EeWUVAJ4k6BScNlJoDwDuYeLCd7D2LvluMQsVaHwfSXJGAhIamWLfti
TzKCsr4jYFIXBoTIrxh8I80AEWbEmngJIkYYv54VLU+sgedPSo51R3z0reynDUbo
8rcV1/sCBoMDLPjEjp94x+c/EtcB1ak9aPe42vtFk0tWLBnMsD/JU3bB3hY3Yse9
hHxV/dGEzcB/xyXNlYVYt3PfvPBOybNGa7Dvw/BQr3uUtym+8k5RKm2m5CeC22Sc
MI6oRdtrtdI2Q72qGCqJG+rljpQ4LFYYabgSa1nWqeHGl3JvmgLNd96eaPrTca3a
IA9yNYTslrN0avUZTPbImHu/9fVViM9rr+vuVWZu23RUyCCr9y0fLjqEcwZSELr0
wlX5Dl+2MvWGBnyCPWaELnoaWynGEiXGwjOA8JD5W8eyzcCSU0Z8P+TLNtRRZNk4
m/iKyohdjhP61oPMKWg4dWV8yH30M4+Hlm+2vL7i5P7UPSxguRMt28dmAd2PkqLJ
VRX1b8icvcnMQE/zL38T+MtTv5fZq+NVKHRkQxN8iyjT9GkRvdXIhS9+t4XXI5B+
Nk9V6x/RyJ9UxK2ArjKGuENjMDlaEYV0IL02Q/7o4Dxwzz/D4jH9/xirMhJ2A2OG
yjHmo0NkXwIQ0725dnjxgExmc08TfYt5nuYAA9RG6JwP31EKO+9W6vU3QTJCt7As
egQmuTCGjSPy3iVQlRgCtUNiBOCvDTRWIECkKI7M6mbTgPZZuyGqjKgp72vGeaCP
Iud2L6nlUlQKsrMGAmpRdkXMympnDeITGFZxZKoRg3JuBJ1VcLReAa5DKN2k8va+
xXxMYf1mHqUpCp2WG6Ks80psmNu938iHjSVbYzLrvQJAJ+/eMJQosWaYdU1HpJ28
C32ESaUOgZTI2Wye8JV6Zho18ftr1t2zXxuiccEkbmHLhXBttmDY9UWXC4rW6Uot
eKkkROjiCy/U9/KnyI+kxLr3ldGuD+PsDdCyR1ofmwa9mugrnIagjdp4y5oua7vL
NzDTeKD0Vcu7+MaMl2EIpyGViNWPLT2o0QqkDv6D5YeAKo/WuRWdyesDcFNrlogI
FVgQNXBuhhDrZB+4KyxIHdOpouzz17SPTNosfvqy6FIB133RjUOU0oxduZUim4SU
2vxx7oDtV89XWpIyTmjCH6nT1cU/JJ+y2PWO82qnPJ2cE9PYmv5alw0OX3dwFjGL
3Zo8PfIJCB1oAn2gshv4q05EvHDK4jPxm0JO48ItouJbnn8xTj142L/MU92l0pXU
KE6XSs9YmLRS+tkAjdLLbzpZv5wPvULBPS3FbcBYmb+uNzSzqCmt4bTTzoG30qLu
SbfAB77k+a9tbp/8MaXLzbBT1R1dSPYD6sQ5/PmbYI3az5nMcnaT8PVKyDcEQifA
MK8+gwBel8Lb581YC8Q5rK/XAftseQojzltBvRtWnYpa2tYPiG02KNGO99lnP0mX
NAt3mMgLtvTr6yDOJ8smyR4r67i57ddBTp/VYkFed1kl1Nb9oJ5jdwkwALbl/+AB
KMpyGC5UFKeBEt93RmOA7sNbYPWT7bK/8hMCHaq/9f3Yw/a1Sf/8vrE2PE75rxB6
7wKVURD9yErZkJJBzLphuGWgRlLyp4du1SKFugvOCUACkWIRHAWr8ZvdZ+ymxcB+
z97Y9YM65x3wEO3SN+SZGcvq/biZrCgNCLJ1sNM1UQYCIGVQlxOaRppbkqveBEda
wiUGYBQgdRS5K1MNeazfKA2z6hqUX+K2PE+9JycdKOTNRt08KZczzG73WLNCFcnd
ynyCNgx3bn/ZFD551l5GdsJ6MVh9n0++KY8mPBoLH/a1nOm5nb4t17Q7Pe18q8Pd
pfI3GJtlndo6Vr1J39SmbH61uD80VK8Uj0CPDNh+yvHuzAsDAXQEVyjorX5UV+qK
b+nlqIi18PrJ5omhqimvocz8B+gT8UTQulvsZailT40SZs1aIfFPYvL1DgXRDO0p
MRMrjSs9uDeettiUYvfGMGr5xBEEOEdZgM7UmzjYRWdjeRie88T7fOAcAFBkzt1D
k0M/iDNLl67EC2Vt8CRsUbF9LSTNUrsVLBj3joGB5q41o6Jp/CkaoH99GqZ/wlVK
MJrPKlT3zTP2gLXWQj+W9FyR5NKSozZN7zdwLfC5i/yD1In3YnpYwHPQIFziXjnk
fzrux0JYbLRbvyzibc87oBkMCVj5nG6SjaDPIYBCtjyVjo2jhAvZ9CiFwuCu8KLr
yhktPTeHA6gy4pd0VkZata8TkMB3RvolE+RyI+pmgATLxgy4DKL/jnBZIqmYHX3I
UMoK7g4MrMAbtN8j8CT4L2zklt710PIedZTvAgUJspBX+Lh4HzvEfj6qhLKp+ho8
GWTHe59IYK2lnEiLsRp30mqzWkB/aEJphVpP7gzjDsIfsE+AFUfxww+xtaJUkBds
/uTQ7cykhkxsIqpi+23yqrGxPsV6UQMahOm9ajdcUyI1Xjl737GWWO3i2USO3tTK
epo1KS4JY5qOBsyuthIpcY0t5FXHqNBQCgESbn8iJ17PgjM6ZfmtMgZCtDv40qQf
vRx0HRtAsAGVOLKfbU/Sk7EaGyZsW9sRebkrg+swmHo5n5UF1C3scLy2CS7WIliS
9H9ecTM4PA6XkxqJsP4aCScFlWixB+ur/piZhzCBFFLqubwuQaOwl/PWn2Bg+AOs
W92YFwbH0nO7xPdE8WC8Ix+Uq3+G2TLKTmMfsFzaPwRT/bkr4x5nIBNIZK+GoCBw
/kx2xMeCUe3tIT0mO/+n8Sr8MOW8LZWbKdfhpn8piWAioF5nSZUlodKtbw0Nb1UF
I6ATtKMqLt9T3mwnq1ziVkjGffXek3IfGSUf4mAZKL7yDBJ2wl5DKAErwbyZsvIy
Djr8fuqRgx8SdDSAGmx1ZwW9MLGZ1Z7s+dVDlmI7+A/AiNJjuq4aSzD5EXYd432J
eq/sWDyJ7b18keU7GWyky7MpssOwK3td60iEj3vcsY3qtOJ99pJt/maBsq0/aVQz
snG/UfUiiyDMfrXBljHCaHzI2gk2C6ZNFaNQPenGawY6OBc9EENbc6x9I8b9CVOo
qgCxZGPaGhpsLxYbdHizkUpoJJqlc73hC/28AKWKCdGLTXV0IaaCPqCM5SFMc1dQ
1ZY7sGpFwqiYaHzSlNaLkgFrXQELq9cxNRU2PgIT/DIE2ooe1tKllz0Q2VgOOYeq
fjOReTmMpPnzN/HJ9e+WGFqYcWr3kM8T9qa6hbn15ccEDxVKUUwTTqZIhGFm/b65
xB4RzP1wpVv6kpYYHm0hIhL+33NF2Yoy75iG6dVVj+E9PwXqOEUeVkgXIqpAh9C9
nMZ6TPpJx40xkueMeEfMJgBxSElzeIuPJbxk3UcFTiLQb6WLYEGCq4iImzgJ2c+S
Qcix4XK+AoFNTOjtGF53bZuFkmiQCNeoyGqcsvE8V1OTxvsYeVluYK7tRhAjqAlk
2A8gNtKaeHYpCmO99cTtE9Tu/DypXb3bimuW+JT6DXQoHu2xYR8F0M8/a/ILjOv5
0HwnUoGJeHbL+sBGkjWIP9KitCYsAB3dRkwg4XaF/2mGpRH6py13pXupyLdPVJVH
ONKTRe1X6/eGdVAHwyAwqo7j40wb1hbGKv1HpbnZCrmnh7SJxIcjmWrDNIJg3Tmi
IwFKF9YXVgAk5uYsqyzvPEClUnTXiBExJblXf5L62bTWQFyXio32tuWJ43QhI0/J
Z3Ph4zcIel3eZHG7BP9u4Amr9VQJkZMZdH1OcIYHp/WIuG05o0hZGYyg6npmc0eH
VmiSrUWfspka/ZvYuhyJfVPAWAjq8OQ0tMm4xCTq1KRAtSwCmDb+3NnAFcJ/+R87
eXin+ZeSvaP3MjwGuEMspCeTmgZom7SMVqu/EkM/lSgI/wrYu7M/kHeqeSIfeJni
invkNu1P63OGZ1TKZqI63rygaXHvURDRX1dFKx/hcjy8fP3y3CHdIqHMo3Xnj+4j
Z/RPZbnoNH4mb3emkh5eZ/poze2vq34wZVkRFqfKk+sfjPSamEjYgmf2tpdpxeqZ
DsXp56WN30h0nx8ThXSdOxHgtu6Igqe26QH8XfAbKr9+1k14fQTy2WS07jWer0d3
woCvg/X5Gy6IGRypxMjlwxljdiaFTO6lu7Xv6828blRbq810TUVy9UMG9uDV+jFY
a5ofQWuU+DzQ6kY1KgRuBg67z2ufdq7VoyIQvw6eUwYIpreZ+qiqN1G9lLDWBC2f
AAR+RZN1qckOeL4R81e2s7gq3bwHakj6pN0TfRXo8G5sjyA7F+uadpnrXyCZddRC
+P2D6KcpVDOuu1IxrPcDIf18f3G2s5G0DfcxYXMH8HJgPG9HrT2t3NzihVIAg2Wj
lLPC4np/Yl/dkeFgaRZXD4q9O7G1Kb6oSj41qo2ZostJoGZAuunGiKssokKRAgIT
md+Q4Gsk7OzvhJfz6RHsh1Xc4tWtaySum9RA+S64qzRTjWpCYgSDjm+EKEVeMsWe
rXKZ5ZLsPlSRNpCgxVDD2ducdAxSVR4u+jJS/eLZKbqf5XoenvCqOKvXEAObT5nT
/xMoCgikVM5pnDoHbaK9AmOI8fdwkhfcMNbXaaLdmlaGdhEu6gcLxKlbt8NT0AIS
qzsVssUF1t5pyOsf0JCwZ8TOfVpfPOWQy+lrQtZ7H09goloeQjgjmxLesPEiTz47
Ae3U+xh76pyF9jVXDL+ZhJnuaB0/4VJtzbQLsmECFUZ6WaFUoL4WzYnE7tDNJKB9
IWL1e7veSi8iPaES7Syq+rQ3TsP44q7Yw2IqblNnybperuQODt9JBsdKaxY8lcpX
P15DgBiMVtZMyE9u5s9mi0lNt+HaAEGCgyZP1mMcPIlBene64iGC8ywUIIjSMUzp
vmiNidoAiXIibain0LGHNJt2l+Swk9XBd0y1p5plS0jGpUee3jJxUaYJ5yiQuiQx
mKIMB9pNH3wm7+A0pFSYRi5+ecbHoaLrDlaGrdHfMeoRQ6YFA6lexL50FJwXSruE
Y3pRXetgZFXdfVyf5KiOo73cxg7oy6pqtb/3GhC4vMJ9KKYSS51h5jyFkvLdXtJN
BygfLrhp6ogY9DZ0cJi4vNCClzE2O6VRNm13CI+Pt6pd2yFRdkc2nmyEZDrGo7t8
21g7ksx1NzFLISogJQ5+35p59Iq3+yPWKt4ODpvO9DcIfYvmdSRmc2rn7UODAV98
C1YZFPX41ASkvve26KitpNnAudOVQkyiY4PoUVzlu78m2c1aWkA8Ye6aBxoITdR0
/HB3s5IS4/7aCOQeF4kUWuheda6SzYp1ShOu3UdLgwEp4AD28zUit0fq9pOHh03D
HCiEfDOJYHCIGLtgpDkCCKPIAogivj3NX8ZyB+rV4X1dS3CrASWkEWT/eCXKoqjb
WxLPpAlxf5jtzKdCY1/0XPMeMHPZuw7DN75j0n+FkG9UDMIzottlqddqI53bwgPJ
+zAdA0MaxEQ+Svj/lBE6bho52fOxLeHASzzsYO78rlKirW4vIk+kakV+Movmm0Y5
J0pcUyZ/bQf/ryybOHbrmB7BC8p3M//Z8rkHqhyw3vxZ2mdtuXo7GO+Ngo/9b0BI
ckhg1vUMwTt5lGS6nCy0DHL6hef8zNcLuFbZnAF28eTt3gsdhEVbskfF5vl1jr9p
MAuHLzVu68F2qq8uapoJSp/8Bh+AM2ivPQnLNijShBWPy9gPlEuKNMC76cBqC7Q/
xuY8+KEvmE6jklLjPHbgk9YifTFFy4870viV4zQIcDTCp8Ph2WYVG6wSeST0YRnj
Ds43KSLt55fbLbGw2Ig6t4Ovm5wKNjIN3CB7sP9dbofdFUZcoMhogTwAGIdrWmaU
TP+DfTCGvOUwqiABc0eVNT2N6HYKj5kRj17YgXQvyqPaIVVNEveIzzkju4g2HVfR
gwZMj5wz+dugAzZ/oAZgAlSzl0JkE3rDNDyT8ekxh5Gj9LdL7+jDJrCG5uA+ma8T
uZViwQt5tPxLsuEtekDa9Xuf9z9CXKK52Nr6N0M3vJ80ck+Mv+uhGrxkaktxqghd
kvW8uC7CBekh6XTD8/O3kv/FQu94+ZCLvBMzT/NY6sLIUGgt9evaq7K8/7CEVbuE
Qv+AcTLQ1Twk2CLWB9Wg8Vx1H5AuOglspxglo4MrHK5lVVL5hOnViJCGSBKf9KVs
BNXrKCMRBOfELE5YcQH5a1oeagMjr2vKMAeYKYBr5T2hUdp0QpkaUlimz4wb1gjp
ZIgchXjI9z1RVLbU0C8w79qfh3BbJukg+tPVAMtSDwhcuf+TT+XLKs1lRPObLDad
KFIcMOMaDyOmMtcCtf1OoFx3AFPxhqAX4Me+npL+RWG6zSU0qskW8DAvbAfeosNO
7f1dQ52nC+VLONDtIiEvkhNc3iLJ3LPk6AzQ+xVnhE48V3KIY5a7lt3x8L/4H0Ki
hD54imcWNf8HRM32HaI+N3EWVff3FioVBCVjyQJyGw7gaUQQR8iFJKHFNaq0cEu6
cElBxf+r5coH4NU4LzXGIBJ/7RK2Ehty5OTKhvGtKpIXfF4Pm/VDpxIIMT8Uu44C
GZgT9aXMpRXx1I8WyVANjWLLfZgpRrB9Xvl55SdTq2ctbPGgO5mgI4FX7Uj2RQGc
7gU4PrmaGuT23H3m+SliDLa4Okgd570STfdqujuySZlW+1wOj+zhQiOksLguXBXb
+2ZPLxpOwM1xWinHf8cTy9RK2UB7v1zVrbLhtuQ5SZMgvnWHxA6T5n4/jXAgVA6v
gT0tYNcMOx7qGbztjxP+mAJYS2887h44EWVI0wOpWJAJWptY0mJFcWHQ+S/7cF+a
R3dv+O1rTn+8od0T/bQ1mYAPwtkQQuOFpzgi/OxCQCZ62RA1fjfJk7F+ZPyYX4jp
zX7j+y8yCZwVmGVkQkyOchvGorRM83kh1evD7RMsIJr+t100uaWpzZfM+UfOpZ6C
nimFGZwNvuIG8nBKiuKYhMpzrEMl1iDyBaEAeI+R0t2EBBQ1TXdqnXIwh3Kt3QRQ
toJPJdpmFYE96q8owVklCki7K7TkzbDM102FGyBElZoHNsd7zFlHCECbgI5m05Ks
3XM70LGuBaSGtduArCDLifBk8Hx41IUK/v5ORs9KnlQuQcpS4baoLL+aeAzzx+Iy
zYZ+WYFM3MbEVPimqKTqT4QbL8sV43RDGjPeqFT94d5xcmkF/U9v6ApHDTAc/MEe
E0Xihqnrdj4JcwUeakkZKxsPcB3jEK43y/1hTXI/kfpN7lSTKP6+m1Ndg6qQ1Zbe
8iweQpB4KAij+hhbFkD2i49pSshCffe+OPuqIqX1Ckg+YdvtAR0nZ43MjywiD4hA
fOkDtbBwPziAHFbVuz2J92troa/9lodtezGtvY/pnqodXinQhM2Q9b7RwCGeqEIa
HLsPqckKc8tHQWDncE3yg41swylN+pL71u46SwCW5E+JpqI4Rzl6Qxf4xWU7PCNW
tPS4wiynhTsWvZ4mthtgSyigNfladAk6hHbaQiDWiYZ41N/VBjinr9M4y+pt0VPf
HVYQt0Gfj9EEzNbi5d3J2fEv8ZrhOyIoaa4vtrVOFALNB6uHJGiskbQkIIBi9i0I
YOhm5QgYqfPkJAlAYluICZfrVFCP9nrpf0Mz6Uw6+GNQ5Hh/8FNlDnHOaBI2Jk1L
PmCGlpwNEzr0zzpYXi3kg24XgnRJqYBsf/jspQCS6XAPP3rnhGRkBkggrEFj40+J
jh9VsknFbFeyYBJJ0ECUOeOslZpc9CDNnvAQUknK58HsZ7vOU8s9tSaGXIaetCOY
CkkveP/cyz+m81yg+fSeK+fiC+hcZCbTu+BwpSYAHGmYbsehw0ScZrEGXTlvaAUT
gDFYam+LoDVQS/yw9g2sGja9i9xd5pohrBpJRG6LMOIq2AcVlYIHKC6xwMCp+C9+
D7+Hg4ysGUDICyNbG83vUqf0abzPkk04yFT97++g7a+LVF8wC86wjF/XW3p23TyL
B57U+t1bCWg0Ae5N2HOJ4shyPsTdmrwgJcb5IxZmXwwAzRaO8VPwFYKsK0qLVVd4
aI/J7UJr91XYI4e5a+O8Qiej3dQmBYwM4DDfOgPiX99e4B9ncebzw2Q3QPdJTIpg
9HIwqRAw+Ed0GZB/pd+z/3aQMzoVDIoofTmqj2H4OxONev08sElJhtMD4FHbDztn
Nc9irGjHbn92of38BnrngO5UbWLArn6deY7Rl1uR+im9/32Ydj+Gf/T6p969p2/m
FbeWtiGNghkCEGLyMe6VJkG6/2xir4ox/867lkRgPymMeJskYgMZuOvLhjcrUqmv
6QtKIQUnaFYLgUjVng2NiOstcRZiNYxTM4VEr2fthdIa4S1VoHK0MPLFe3NbAkZe
uLP9TSv1fEn5lCHoHvHRy6xgrTKbftKFY/gDtDb4stIYp5tzz4cfRRcti9wPg9ul
7N0ptQf+2fS+7tKD6xUklt5qBeVTVjNUjDIMijwU2UI6o7b3NiDraBlnxDDnXC56
zCfLzuTfYECK0tF+LkbVmwyUZXqvmkGLVINyIdxaVSDM0Wcm/3Ifhq6u6st23+oV
x1wAkYuuEugmer+WSqBSnwc6WmqC2a/dNvFwmfaNdpCxnpAdl3g82A0Yoz7lmAQs
O1NkesxalpEXtnSaEo3cB5oyR3MXEbSyPnwB4kGCcvzpUBuiJbcuJH7b+NiRGZcv
dXvcUKAnKK/1ixYoFZzf02ZpTYnXd4NqrEiD4687HWu/8sIIy5otMxtYFHxNvWrt
8ZF6bFIpnHR5PCmW90EGV/hHfT4umGuoYrb9OzDQTH0uH9wMYLz0Ae9HQ/mGu+oU
+cDp4KFNiOeohKz77Xo/HqhTWBO2by6zfyOdhK0wgfCSx+/GdIAspbf1iLlf32pI
/j/XtEGtzNNvAf5HknlxwJF8b1qhqATykc3Sn+DhzWvjllVpXkMkmvZKB6sDVqyV
hfPRswnwz+Kl1Xy38SjJenwXet1s1+7kLOPs45mGBoREbKmGA9XlsJrutXmdv6DP
VjqeCicEjldRSOY1SNQAu67c27eEZpZn0jKEpXriWMJ+zo/Et40mJKKL5tNL5oI3
fGdoHTxn4QnXOgq6NM6VEvZcI1VjP0ejlbizQVs4R0e6Qar6elW1RaLRX/97ixov
G2pWyvmUdkuaVwWrdwxmJhCNNxYPs49mJHTBBitli2W3VQGhG3uoMaODN2LhMNpH
QNap+QxAjw2BBGV7yln9Wvh6l86tDTTYv40xA4Y/byfVE5hI7Fmp003ZASTdiqY/
oyITGVpyGLFaZe3fRgM8uiJ6lgqnPPmxkaWfDQWbo6gTLQoJxmlBs5GP5tNq2jS9
pd3WIaUb6VDOh/u+p5/kgZxAA/im05mQ6UA7yP+0w1o38oncW6BsuCYczDrPTeMo
XZXXoBCqU/hcdSgbQs9zll/O0xxOuVQqfwAknRW5VOLdLKwWXaqE3E0ShTIpYX9s
xDIDAJAetBRTUGWVM+tkf8q6Kr72Lb8v3UA+0akHZZRJ+81D3U9x9atlIDROAiJP
svSAL3DYf2FgFUza7GXkqIQsFepRFqcfRNCuokggJXwc4lkFwwGGeNuMBnx7/HCk
Y4wVEu+gCarogFlVU8P8oOU2GYRxH3lmMBTjFaTZz3w4MpDV0XPqbE1gAAmIY2eZ
nRq9EqFVRYSINK+r0SXlCRYtvZOTCr+ZVRFbOiS35L9aG/Yso8BqsJ88iANxrcf4
RaZXDcjSjd1Tf3lQA/NBYtlRClE/rL4MPfO9I4PnKOLocduHfjMLPZ0l+R7M5LWQ
RPSeBP6t1wQO+Ms1zD8gwgPENlSko0lC+ANxNHifZ2FEt71e71s2UIE0/CYCNEBf
IB/vrJMvvhf/ebiBNBjd7LQk0fj/db3Mo6J/vTZ762hdN8ZlY5lDeE3020lgSZ2Z
csa4g8vFu+RpJxa54rW6EasX0On9al3t7iWjVbjYkfFn1YZDY9/D0DMfVrUCo93o
P31ou1OqRLtLFeOP5/QHDLI4zZ9Bue1M63euo0uGelRl9LzqU6oQ324Kl0vj+AkN
uymaoGRtzG0ZxHzHEeOxPOzjSgHmQ5yNp6N/Dt3orI5Hu3tq/ozauM6WUGf0kE/S
v0HUACQvnEPr/Nr0lLLVmMde0sELK96CMlHDQd2+113ztD/NVlqaNT6x0G6aLXm2
KGFR0dGCtYxne4bD7uPfjb99saB8rCcH61e0lThe86SmmjNTwUnQVZ07nhh9RckE
p2aNsSuDKfPOSXbbfkrvfcrhrudV5nXIOVFhae5KWWKnNlnzfo3oSkq1W5OOrKXH
SaEc3U6/a9waINbRB+6O9zmOglzc3AVuVEcIomTKpA/THC5XhihtLGxeWf9E4xsh
dZV+kBtZeTYxzqWJSFao0GKxP5IoNj7UTYWIbCRBESugTMcFWw++z3IPgHdo1VXO
wRHh93j8fElNvGF/F9BH6g9VusaAnXbdBtBfScusoVavdg4g9jR60pY9SgPGjHzE
kqG1tAoCIeEZRlxAvCTAQxrrL+s42/+CX8ipM6Qdh+WKEbCkLMfqQ/dHZguZ34Sn
W6Epn8yx89DlFn3XFnhmDBlLsFIDFzV6LfzDmTol2INZCWI8wssPJT7CZv3rq4Vo
nq1UR2Z9gqKwJKWSJ6yEtaO19O0ZOa0h9j38CNXr55UdA/oCR2SC7/qnRx0JBDxJ
Xmgj+M/rrN/H/Ii99kPrg3Z1Sr/IPQh9m0zJfZskUxmPrxkv3J2dZtQPV+7dIcMz
c3wQvKoLrFV8fdfcMYP81EWYSPgg021QWGOzNgVLf7sFQPPAHh9gMc8BeD0Ab4Sp
xIYl+oKjsBDKUYNPnp0kUAx78oD2XMFkU/gNysBe9gKzuItAcbCPtsngG0jyBy1Y
GLJJrhQKpiDh7XpsT8jIlBkkfAL/qf9cgjH/4KFRus1fUkNP3Gf/wSck6U97CCAJ
CbVXH1pOTKQD3avt+3AeNijuWjxZR87GkrrDz45pDR/FKdUdNAd5MMD7FwppLW7T
BESmA62JJrqS9ywiDMFEvi9JxDNJT/vZDr6LZvkQRhgrpNYusem+60v4Db26K1jp
420Kea8rertKzxg6fpmv0oLcNXHkvEMuyOPrqV9t5rvywpdgZ1NBkfi19utdj9th
j/PjBEKZLULZoa03hy4as/DG6t1ff6t2YM/w1C6nLLAoPHNctZWg5fov1OKeCp3e
jSOs457LNPMcGqIQwDom55t56p83Cf3nPwb+9g4BV7ueFv5UjSRCEDgZRegpCuGp
3gwItDEoZF/SdrkafGqFFfcVsh3s9gIeqQWysod5rhDf+G0WEbUVMS+F+aFNEf1p
qEG+3GIUE7/smQ0VWnwaok7n7vn8bOKVTKscOJR3yw66MEELdTnVd9BNGUuSXwPO
vvqHmiq/CJX/4Vt25/eswLXNF9DtEZMJPre1i2rYDR/Ck4Z1fQlNp3gOS2ogKa6o
hTjUm7OHzbqZv3DI6n2a1TP5E2ruONbs61ggSRTT1UbNykA4IT59ME6wwB2133dh
TT3qdeDIHD5nRa3oMc5E4aFpvTfuvfoZvhtOSGJUumhqjlLsktoVjujOXqE/PeHu
E4wzMYxPJDE7cHQxlFFa+8VEi3xNXNJi9/692S6L++/H1oEl447FuXO7B7PY0Ylx
4Mu+du/xo+mpPAZcvDT/CFwQtfCxJvVTDydadA85Y6Hit4MYeJbu1L3/W21vRWdc
RUHWYWeQnmlYucK5T+loJBSx3N5PVfA+ZSY8Omsj1WeOxpXP0PY5JDLboG5uJnGd
Fscxgy1Mw+ZNHGJgB072+6Gwumv/H/wyeGPGvgpPDCCEc+oD/3TM6VOub8p6EF6u
e7FuMk2G0IOnmkLER32e+yyPaWIj6JwxOJ9Ap+THlY+jAe2l/S8huik/prYJOnuW
U5oR49pO64/7DAF2QUaKaFG2JPrXLJizR3zYDiernEhqxCVRzn/HRrS7oZyQQdZA
9x6FJGOemSkoA+f6iIo6PcxQh1OjUV93yYFlH9vO/neu91qU8PF6lDJ2waaJPMAI
3QQfASANop/V1xfQnZ//iS9C0cmdIldchYZDVBPhbctw55AFvCrKSLVYbfKSkuFV
tmsj1ds8eqwVqHSgxzF8xuiiQuFJVRj/GmnKgJuIGwNKWlfPZy7GiMRWe5OdUa4y
fV49UBIUE9VSve+k//L30a2E8kSJRazhd3V53dvbw02I8nEtFQKkc9dbZpCDqVx+
di3jSjBDtxHFGAUDLANRxcEyso+VoWKFHfTCZCTHqrshSmcoVXzo/Su5KjX9UUUe
U16ckNAu83YIkKEbIC92yYfknn7By1RLw/+a60fUJGIo4HqhyMVZ2tvxKYLp2d1/
/UkHRG4+/BpwHgCPrpqWCNAS/5JY5Szh3dNA8W1Lf6O/FEJtMa33kIcZyZt7u6Wl
DqkN7BvK2ixCEvHnNO+DyaILcTgJCfzMKT3M8vTuGYwKUDFuaBlVIGhG3tYj95S2
WGKs3TQ5svTL3hWTIFLKcFbO3bawrvNmFNMidjdE+T5y48udjX6FcWX1vVaF/mxU
f0w6VeZsHvjg65BDrzEPWhGjiAU4pQSl5cXJXfgSBwaGpmfp7bE6YQFTdtcU2ZwM
MqHFnLMFgPtFzDsyUABLZb+zc/ZHW3NiCvLPI9jxWCnGLQn9HourrwcIWA38Yt3E
YfOPwsomDz2OilKCLw95pvJy7mnq99uAdy6DBgRVpLp0aF5R6RHaPV0Dhmbfk3FQ
dPFOFP2OUowe51ceZaS3NWe+0Shly6NVCjaSdKamMs68+g1qVV+NTqoktv+YqXp+
wC3LgGrtDk6YZZpHucIflEMehM4Y8BbUKud8O0+hgFZCHynL0rKy9wYoGxDzb9fX
PeW62VFpI0c+++4mMUs9W6z9+52aoh44pY/ynaQutnZml6o2uNlwVXCXaQqg2ByF
rwb7L8kdMauCEMRcGSKUOu2rNxRmhydBeuQP1JY56xy1O2xqgLc/apy+lrcqJJ9R
4ZxuliFXWgM3ZD337s9Vogqoh0p/D4JwXtxrKoTOXrabDcKZhDtmF0r6q00TVuMx
EW0+txnOvImPHyZW7Hjzd7eb1tTR8Rw4RPaWYd8/axFMH/tCw74mWVshwPDu8YIA
rKZZ507VDx2gKGihvOxxT2sfnWTNtm/qHp1X5G8NXU/W2FU49zFSCfz6g/A3SLXC
7vzaals+gwDaJHu8B9WVUUw65xPq8Veci8KY6VO+KMABQisH+wVKZ2GltKmZqH0l
NohCQOB/avLrwlJCetQyS1hoYGsv2jP90+2GiYROSvRWlFvEPEZUQqz9/rFmyL1H
SJKzG2FaW1rGuvbZ4DWD1IcWR3vortnlrRrva2Q23Y3trhBOEgxl+kwevoaH1tlK
JWDcCaxx+wYcCKMX/e3wet9SXZC3MLw3XUHuQxDsIag3P3kD3o6I3QwjJGu4tvFr
5Vm9514p/1RS2F0AaL9Kq0ROukfnwCAI1tNFjV+wzcGNCCTQLyYOxk/VeXy7oFOx
97y8MasA/Viqv0dn+U1gQJqFyjm8iQaSx1siA6C7lI5lVO3NjSRvdLZ+hDqHaCA9
c0P8pD7+5BtyG2UKEva3zzNEOcQaygV3GKaZ9KDMgkArbY4TIfSyDzcNVGmLl0PM
NMhmG4yqzSj+iybXs6Kj0jifvP07NaV4lW8Wwbj/6+mhZi7U/xsGOb+8cWFC3dmK
+egibOUMrowClLPthLAMUxsQWqtnuiDNWLpPi1Ikfu/8XyFucJcYJaYv52lRrghG
3wQtch+/dQUNIwRS6L/uE+sa31CTU1uUTFEHuPfLQKnkJyZ5ujGUotzw1WlszTRK
g30Gyaem+NS8is2KtK1DNRKWdekSCB4g215ry8T1qyxXv4cE4M9fL3fLZVwnUBuZ
xgGm4HPMwWnmnvmD0aSnq7jBgOc4fYTKdD4E9Ud7cNfwJvVmqwVlq7uCxx/pZ6O2
Bod3VtD93Qqsey4GtsAWSNZfwFh2y0TqY+vd4DIdwdWEfFkLLU7BnrbDg+NS1gAR
UjmdW++Us0jsUpct4ks/6lU1COqj1sCqJKsJHX/wWbCmGOd6bCRLQsgMNGsPnTjW
jEjSc1pXlBIQvdamVKq10zSzHlAP06Szr6twewyqCIKs3p40/e/Oe7N826iW02Ki
wg1Qfem9OY01mWy34+RSxAAtRhjcoQcAAN/XEVeHdyrUgyTtkCkDPO8uTWlwJiy9
Ga0j/8r8/K37MYq7FPgVkwYgGai/KN10T9/vgwrq6sBW8JQemtkvQY6BRC7jv89A
oR659+Xzag3TD9S69OFyPVjKX+Nd3KA+9gaYPb/KN09mvV5mlfIR/yPERicfseIV
zLpJKxqkBRWiZfC5ieNMiPJ3OvpnLFPWZNKMlPS4yaeXy4G6N9ze4ujKDouyjqk4
AN2eenV+zlXL2rnp0TO6X2mTkH8R9iz7lYIf/UCVoagtcXrm7kNapEpOfSykv9A3
s/uvuFPixbCTmpZjMnaRy71QmAeaJpqZveuJ4nolWjXSEqlWs7bjxNGNIRj+3Nr1
Ex+m/tYrthpJmvhvzVmKHhlKFi4D+lxkhQrOsj2QyJFdgTHOEc4bcfT3DRZ9Q1UN
c0+9ouraKuBkiPNmtAo7xMAz6i6IdThEXk4iwoxy+6JFXJFN39fGURS+GmJb6wKp
F0Jn8ZnFm1jvSX3Mcf5QyBloq/gqx9mQGHoYdzYtLJ5GnjCQkh92GZ5FrLU0GcbD
VLbayaB82xl9C8NP1WXju5oopt2zO7f5ubHU6VFRGLRgmqn80cYY/5vu/a1J3EdV
ErJJ6cB25MqcaH90IY/oKDuDyZZBFx+nADuSoR8O8UD6h/J6D6FEq1/bRLYw9xnc
3F3Yac+SwANRnN1IxYOPhX1KvJ2e+fOan8drtPQzUR3S+83niRUZUn5WTlCCVss6
ownV4eSu2kSHwYa1zsSCFnrwykATapKzAMns2/tN+C+ZIZ+UOVZUQr3W+NM2qy/0
Gag65vIU6w1ZH6Ok3o/N7RMthWTzfYa8bLHLrZ9Dqen14A8pnOnAlBoRLA8oXCTP
SbXQeiGZP/HEyCJGYu5gi9fdfL/m1t9NqDa+A6XKNtNuBq5UeV/Hxxca7Ii7YRCr
hcJsFK741ZWcV9mJoZW4aRTNFL30uoCambRfdsem8MLsFppOid/xnSwUhhaZJ1rX
uN9thvF2NXELGuBRC9VBgDARqL5SazbxAlpPMBa3O6BaQ63bKuAMzsRLKAVgqSR1
59BEjSabNflOSR4ZU3gu6nohE5/4xQyUgHkXK0WRpGUVLac1yTiq9ACnJCC7d4eR
X0f3aKHhwbLqBYFvhGC8uME7e3D1Byc9VO/gyVWwy75eA/gnxZE/Pu1VQGvS978I
eD8ownm/1H494LSbIboemqbdHQzM6pfDVyL5GSoWO9T0EOQ1zF4ePgO8oXRb+plb
PCabO/LWnhe6iqVF/r39ukHsAiKl9pWw1wVd+8ai7I7WSVoaa9ZlIPniFbWJXUsu
FoDUOhS4+LxUqz5ZZMraPlrvfkiDRR6bVp04x8SQN5iNCR5gae/KA9yyWsFfX5Vb
0Ix35rjEB8uJZkalXWJKnQS6BwrG+gIhzrchKHNVjOb2zpAkM1dikAUSo+VR4JCi
jcY16DGIHYtS+pJhE4/7CGJj1z4RJBagm9le9STWPJ777wKBm356M2jTqEMVRVWu
SaZNZShrnZoPV7RqUqP7skUHriFP5lvHXnT1+T829qq5JxDg/ZPVgqi7A0sIgup5
AHRaPem6MWg79KguuaEHGS31wucjgnpUqOsZJyWzfMXSwwczArgPfCVxgEaQSWOp
uSET1S2t8ZuU2yFMLUNR/iky3MoOwGaX+687K+EIo9cLsAFxUMIwIDUrbb5+hVIx
XO1X5k9emOl+I9P0XCyv3kwL+n9dFuoqIfWElvmkbS2+3nqG/7ANGW772tkY8Xw/
RC5tpM5/Pf3n2RRMfxPtMtX3btLpbVZHQknRQR58bpd7u+Y4CPfHpHTLHBf9oPx8
4KNQI6pC7CI9BLG6JKXhH5JzBAVT5cTTzXRg5B7F2JOYwPpaD0lPW80pMxAyPIUh
eZpGsn0XP5tDpgC5Z7q92zHUYOpy6+hxJzocALZTsUuJzM6icOQXoWsN9VNFO0e6
6mWysNwdIWZmYEErKWOXeJzEea7vrFj46kTWa5sz4gvrGlq5A3TPcEjuqLW8omaV
J3HFFTRh1hFPkE/LYjbNVWAaMtem6GbocWbX9S/rsDbEHQ/vDnuOMyweor1fd3OB
3kqtoidV8eECTENTnTiY7PAheakiLmXXetETuGEUA4qHtyzQ1ofZgkgOSxYH8OS5
Oc4txAg9LGuzaJcmHfKcuUcpdFi9DUWGXXRdE13YQbl+8D5vqjLHgCeCldVN8WEl
GG9A5aJNd2hMeOfzvOfSiZCvlYbfBuEl0aK5gFY472eSpQw6rX5VJJl08Co1SzBd
UQY3WpJyeW6daZ1wBbmVhohVPQwNtSUQbax/Xv4L4OpomsYdmgC9M7+5Nkg3Ekmk
aNGuaiXAwBR1yDzH5kTcVNR4mYjBtke09DGTS9UG48FVdPXPQ3bClW/YL35KQ55d
NoJL+MiAxvMcPqZ8qOh2JqHR3dAbLiLQLfOryKxxZJgvRF0X4NTYBwytJnHypOwr
cM0V/c4wvV2ApXIFx2iJXxecECFMBcZJegNSpmDFm1l2SSToswe/h80jyb7KrxmY
6PdjySjxJmWvx+jMlErXmRSXht7EujUvwWHwEQpDWmE/Mbjk4STHIDeFk9eI+nVG
tzp1OZCOJfQzujKhs8cCP4cZvii6c6pu60y7RG+rRRKl4Nv/MWRIlHEmRj9ONBVq
HCHWekWVl2ktmLyn4xQ9Z3XkJzr0DiVEmezlhFBZsT6xbmJzHJNdGuEYd8Gunkb1
W2QAniZ5g3ofdXOqUqPqL6wQQaNA5YBx0yRZQLQNejJxGAm/X/9nnxU9ujWxCCxP
JMaIadD7RGV3YtDMZYb0f9ZIEWzjCVj8936KON/3gJ356O8iLK77ZoWjN5oyekjC
gBcgo0K6hBxf8WA3QiuV7AG5uwLB7PT0Myjh0XgIXwY/pUf+k5fK26hWtw8WEJ/w
XxBEDhMqR2EJvdzjbfvyEsMeWYbMD6k8p0UAiGB49/RdvdpY4FwwtArJ31c+T9eF
MLQyMKDxFYjcMRccNQkUR7L9q78ROvy3ZS3Ie6IOywS1xC6WxmzVc5I0Wxx6PrXr
qjTH1x/Lq652qQdF0QCKO3sVvEZ08P+gMKfA4xH7LkBhxPsI7eEYcRneocWR+GTA
kz+wgKNtl0QcCVuQ2Xk5HBuZiGjF+PdA+npiHnGn1M/J4uCF3ekG9tIZUAH0jKk/
4XkY6bQmXAT6SXUtnEfxw35Zo/hw3R+OpMnOMutEv1D3NKxWAyexTi7SaGjh+jcF
RpF2gRjgka4dmEop8HCSTwuCY9uuffhWdGiYt91y3oXuMDsluijs6Sn2Vl03X1lZ
EaSBBdo7qVXmlHaholIuZykeMMmRd/67QjTPv0aVgPTcrcHs0VqsxmC6ajlzStHj
TLZqeKadRgEaIStuPyB4ptJKJQOcZDTMgzh9YFHOomRC6l1QNDJTFN6JVwb4DpJ4
scmQpYJfT7twsp5vNk2jAbFinQBgl8rTKSRQ+N4/1Ou/qtbjad37b67JGpHNYlkT
2z3vrfgs103cMfZDFchmn3pNxYbKufrSTjtfH33t5iP4cjgdxSmFPNzJYFZFrCmv
yweN6GApD89+dHBOOKfkvG2yRqB3PYB79Kp8H0GJx9rWONmAlntQbPWYAz+Dchiz
hY72qyBpfrlPwl2sh85qWQg5rodTxeaeBv68FEdo5DLP2Mv51wI1GJJQoEpiY8g4
LQrxtAFgmpxWUX83fdeQtujdU2ePsr91Rxe1kuefgnTH0V1AfbZhU+FoCDOEV3CF
GxLBI4ibGQMtd6A6VmJQoKSkU47TCxtY31FmZyLR4C2Lx2DYLjEarIOrcj6VOHR/
/guTUIFwPwYTHZ1X1f3FeC78COoKd/9EcQXxMcPaLr5QpDbdRcGMgFc+7HSQLTTy
TMYfmNN4MEPPVV8miMLVrfFSjWPicqU24fj/l6+sqziIDZ3AqLYdO0GvwLSDp2ah
/355uEzFvTjH+GdT/ANaUNCVzcqbE6OjF7MtOSx83R2ttZTY0y0UyBqDkzqsoxtb
6I1GXFk/auaNySnCNeTBxZJH0c/oPGGd3rb4dK7ZEGeHa3wPH6VlVqAQXe2FlrRD
JWTZBUUe7Ymk+cQ8FrS/w/5hErnj7iBfsKVzhjUK61yc6H8TjlxyFC8JGdxcbrF1
P8V7iCpZV74IGZ8lzSecPk4xsDZvp1+SZ6f6zZ97hWgclld5+fVvGYhZ8tgJcbT8
DjklB7TW+puPDqfqPlT3BBx4oWBwquEjun2BmBi6Sgig5xd7ekdGSoAuMI9NAmVU
jcBvidi9e894Laq07y/4jYtBaAgL+EmLSNapT1S5ijSIHBvFr+J7sfrIjCP/pvb5
UwTSr5CHVNnokd5ImJDJ9F8YWnWRgPYaCaFDLfqk9Ek7PwnSTXB35qHl/yJhOYTh
QyANKyL7++5GiJOy8ltBIrXua+L3bZcSk97gRvF4vcNgc8mifvVulwmtUSnjdC1C
4pE8Z6pCWsmdRNIEUoqd5fFdoBJyS7nPZUMX+ArE/4pn/kLrHzW4e9jfqsc8XA0D
t0e5IolXBp9qTmcl6R1t71R3u7esI8dSlxW93buWDlvZB4ZEXdOOXeo1a3RPOlfu
h1nXC1LiKvu7SP1rzpAoz/4yOPAArgo6OcHFQWVZ355s5GdaDw/2EAd5++SGcxAL
kE07gT671W+P9+x8D3dFMngcUYsB2ORVn16neLJyH7KvM99tgxrjI48ltUGxoOPZ
twoFHB1DQfiSbFdOLFU0A6a/JsV+iGf5yztq+8qThjIBQ4D2N+v88YZ0d0zYY0NE
xQk39s0D/GlwaPXef0tkNEeeNAi9We4QQP6W0UbkPQLy3lXtaMoN3IOtp+oHh0Oa
gazbL12llud9Iu38TDCZ+tT55zXGVTXvQam23tAGUI0aBRHjqVeszhABA21Gba5c
LezUrG03GpWtQU6SsUxAUzaFnrZMJrUUetwbBogZB+7mixpk0WlwRD0Bx4+mLvua
3nYqJ8WmyWeoq/LNh7fVlKMWMPV2udTKMAYawpLG5Ch7cgg1czf3LQe4Su5dwMxT
uRRD9iqcDzYNSyiUEeQAlTG5RgW9DsdDGEOULac6skl92IbyfBzkMzM9KMY6vhkJ
VZUPB2hZSuNU/vZE4MKmz8uCfcseRyz5YxxtjV5J+F6xNATRmiZU4QxUfZ/8vToS
l44HZd8HhIv3sxY7IcavG9ZibcGHZNwHNB8Tx4W7Dre+PJ/V2ekIbKqpzv0gDSm4
4C4qyBb3+/MpA8a6t2hshTA32VjtayVCbBL5PkejOSiXq/YYdnOdbIKpd177G7Jn
WAWcC+n/HeP/55WyFkgPhF9KoluLpJfdXb8h75FAd3LOSi4NFO9Ts9sgiuBg5hY7
zwbmyEnCBmRMyzy4+f7eF7r2pfqh12f8okW1mMBNsVtJ5VNW+lW/sI16OWBqfpC4
IsqsQ6EfnMGJJzss5wMY5L8vjHVnI4nBV9JQYlmJcL4S76u1VHYwg0cuDhkGbrgE
bCXPBvjCKuC6slCprUNL4CsukVHGQyb1KQVdNO1Km7KWauFQCsrYYfFct2HyCoPJ
sVnenJgR/vKDF/MIu8Uc2iuMg8XsvTZQi1JxIkbzqmdIOLZcM5va/z9pxFBOk9R/
HONKsYNVfY9OlC4pyg5qhcCG944DmpfSWzKZdOhgp6F3RaY2TlFkQxBMZQoIfjAp
3WitVuJIkiVsBBlKzO3vLMD8Kdz3zwzaBeWRL3Vxfn/wyky0bhUO1Qb78wEVcjg0
OF5VMaJ1eMpsCmdZ/XZLxT6aW1zkow+CUtHu1G+ZAKjowvBEM2hCoK1RkQCLpLQO
aDpRbzf3rn/l1nUSDmlBc0Icb5uC/dGMNYLiEyGFA+7Ezm+q/lB9gjMO3+msObWq
ZAfSAby4iFzyCo4uBV2erHkCUpluQ8HOHVh6ZTv9hVAiVteBdcCsVl9KN1E65knG
C0o6b+FO/QtTGtEf3JMBEpCLWQv+7ZOhjJxHokHGcB/9UFOSQmZDiTHqTQxz3JUI
1WhX1KjCfqmVFKtjgR84z6PeKIqj8InkHtDFTMg4BUzSY8ENgNvjAIJB9TkyzKvG
O/Z0w5w8U2JDdLtZuWpinEEz250W5l5VckID5sI3vrC8hoWLz07eEZJ+OTr++U1N
NCEi/IzmTCv6r6gBBKStSeVywRlpCHPLkpqTowIjSBTatsFiDPsr/u6oT1rQAlpe
liNWMJErN0fzqyxTr1i7fSFQXe7dgfx8Rvx58BilSyixTZCWLVM1FyUPw0MAPnzJ
HpHldfnN6gGiwbW4fI8GHeSDuWGF6Zg/G7T7BbnwrMrh+mT7a4mZ0FntNIx15rAV
8XT1lCVAw/mZX3/E4DoJHRXW0PeRoxXw8keWNZYOB941XXQqMlHDbqnorUiAFXmL
y0pdgE49MywbyrI/7GONd94HH8ZXnU7xE6dkLdRBhsFeqkMEZ11UKKi+vs5pOdkn
nVk7UT82H8836Ypr9t3HhvZJ/aYBtHQ4xvvsiiUNqJL15zALyidi5F6A4zgaTiQw
nsFAWSqij3TeUYKh9ITmmnr4DnXK/au0NR7YohVBOjW+rx2PIWp1U3qqtxazXlNJ
6nqvwbmWCkPI25TMS8KQQ3zJCZi3NYL8KhQ8lXL5HJpBSgMRbTylydYfiPTgH5AY
x/rFAXr7IpZmuWymb+51P0rJq41WgAunNiEGv7d67t06XQfTIF+fX5NkKApm9O3t
dcTJCNMZt2Hi3xF1jGb5IUuR67oukq5x9qx3SiwFx7YfUXaZDxuL15sRoluqVwjG
L8esN99Od++aOnDQxFfteb+3/dVRA6mtWwxX9CbbzGzkog9yzD9JMLGLuYNwCfN9
Nx0/Fahg02HeYDfi72aEcyOSz0YWnttWlVAdJIkgvKOzApibGlfSyGcZIdx33+Lc
UglNQZmtNudO4HRkXXHUMuex7u85iM0aXWuRCx9+uYS3KZQmqN2HW9f9gN022gth
/npd9J4Ea1ov+0axuufCilP5u49WYn1h3LpBOMNyeNiUqU5raea5NN0L3Pfj//6x
U4/zL5EYPdk1CWpN/DkFj+eJdWFcqQPNYLlkygaersRY2sb1+/toGLCw6fyr6kgf
7O0ZwTbYJu4be8JZzztOLFsJSCqK4kOkxuboQNxkU3/vB/zKOCPUI61PRItDTJoB
rI3XmVuaxhY8VgWl9hkx/W7aOcgw4qOob9AUrrlZj/1m5uaqzGytjuZ3pKbukE3m
+VI805zQuzKGSmGtwi7Obl3LpcOrEIDPrN9AlK5Nwy385RR1gyrN5DwyOBh+2Roq
KGK1lSpcf6mbhN9uOGNeCOhn/b4Okq+ysj4d17s8EVat7L3f9MDo/eG0mbaVtYZy
uK3UIAzB+QPg91D7jwcUeyLXYAx0iQIrZ7BiMJ89nAi6nGk04hwJh21VoH5GCQxF
BGI39a96i1+PnG8y2UHUUty3C6Qr9hqx/WoTiB9x/CyGAB0yRTUjDhiYJ34d9cAS
fjMfCDcgyMlaq1Fv+iM7jYRLGU3thbk5b4qiDdVLd66CcRD/I9aIKgTxRB+R78Yc
docoxGXozWw3qtkaUv8vGGIdwo6Ogf5B7Kj1u8bvQYgtledrehs70hO2XCPMTifp
OZJu2G+rHaqdMbU3laUqfpuDi3aqHDfZbkRyGX14yy/aESLa0cWcU2Yw3U7SDFOy
sutL0BOCSmMlCo4HgyPXvXfm7+CalwurOJQ08Re2lnnKsEAN3KBQablQq9tZuAXF
p1NUDw/sIZlcNHuMWkR61SO3SBQNBMdudXEUhtV6G3lESucsJZmHyaTkzZ2nJnlT
X/w2Xx+PCnZXx/a4Iwkgbhu3OsY0XmoRPuhFRxnREdVGrnZFKq1wrCmwdywK1aNe
z/ITcP3aRKUnq2IBFlmZPhggkhh0HKJ9nYf2Na0EXpaXezo3ZItdsHCPcAbBiBMS
QQsuUB/maLT9y80v1WwEcqcXXkJ2aeC0K3J6FpR07gBL4Cmv+irZyJ191kqmKyVz
K2aLc2s//9KFgN+dl7bQXFTxMa0ysPXsUJ0SUbDGNRCizPUtJaFq2doSDC4FMZ2S
UnTSBCyW18NATO2mofn10Ucndk2SoNS7PjMg8La+lta3fVTA+1vEDN8eTCzIYbO1
5uDyijU61G93Hk8aNcyeoz/kUvSKstIFxeZrQby5X3LGWS3O+HP/RbaBnUGQHQMp
7xCKm1NFMQvlrB53RMbUJY6uHqJWHH4sZ4b2aLyUGLwgq2/4wG8GSlXsgX9U4GAQ
BopC+4hvKCY3xXjP1TjbkUYb6MpTuaQPCBoPxLlBt9Px+3zhrBtCJJN7kMl7M9x1
PEKxhRqUfWLTg7YSF8wAy4e2mFqxVB12OtWa2X1oBtWhHOboJAfl4rePfBtoBb4q
e3wuljPAEg2id3Fz8lcD+MaBK679r+kvZJy/kFqZj27lFNCTRhf93I6E5nentihc
EGVtxCRCvOm1KnmVnzbj1EiJ64BhnuRTWQQnpe8w6+OUBQVncHWJvY2sWW7r7VUY
CQsRAJUhm40i9p7R/8Rn9uT+EqMenAjoAimHYdjMoVKnRjJExXJjsj4Lh24RUxMA
LFyWIRsq/1Z0SHxSzq5dtgYgs8FlGeWJwwGAzU33w15Cgj/smvsN0cA/YelhMlIR
XLSLyilj7mbdheVErbY22HrQ5NC7tvs65HXMWNcVRTAq89/U5LfK0/Y2h7ZUQsBy
uEV1MY6rJHa7HS71y7UdAw41G6M5q5VR2L0Gikw8lgDDNWDR157ChIHf2WPnYSLG
l5YsDR2p1V+Enfh9ac1y6HduqcZG1FZImLI3inU4vAvrPUWfU8G/9Ow7EAKDeqyp
9X9TSYy/3+Hm+pxkpxwRxY0sVH8ls0LAUfu6ULcPTiULWHAMUIH1EJGg9nKkfbzi
CV5E1raMMXz3IxAYQ0e95exS6L4+rVjOrIgqeLEM+0otBsVR93++hMKlSsevt6Pa
eQIyVEBzwjZahVXIWPr2IgebZ7Jj3OkEPnq1qTAYKpeWUWyQwQLprZjNqHMdwGrc
xUOMQ1ktkrUy0mg0zinIzi5Luhdp2C12MOQuoJDGwewgO4h7Sh6EqE0+8iwKlKdY
0f0AkHb6i3g+47zHn2ysdx/z9thIV8pAb/roav16kr0hlSSxjU5JSHOKGi5jxn+8
WZJo7SAK84cAvkd+663AO7PEZ6H4toGs1UAXGsfs0LmrknK91dLWHC8PbhvYua+r
OBVG/tAJvjvDzplAeJgoJnoPlmRYi4/CvAl072DhmpqVtJscBFnvjprwIrRobnvK
1EZr34mDKsO50YL653QllDsPULVRhBiaN5qAcp6EmgoYCjCC3RkOpRxLlFQIAiC+
+o+LR99lKuY830WqthL5Se0FhHyXMINiNYFtf7hqcKV4HtJG2oKBXvCWpkWIN6Pz
4ORKi7NW9w04+lXZXR4kARUzb4bdXvYTYJNjdAm8bs9V/Y76ZDJM85Xe3lUynxqk
utPRC9yeaqUdNEVIDzZWMvN02EgCIVTyWPe1XJujGnNe11zJMUw6iXHDN7Tn/G3m
86PsEfM4po0dFf1sFZ5u9M82Il5pAH9Cm/Bf2WflJD2UGbYFcgwOmKr4lhlzMVPb
54eVLAdAzuEI2Fnp1tCrYqciInf4seJ9W0O7TLMw/yeKOJN2Kkb63tn1utzwaLqS
6V/xD9DP+ZuD0RL8cuExqkNGak+RxUNte3gav9R2l9AxR80w1r1zfDndtcty1D1E
rELKpr8jK3trpDfTXPPsc3J3tw0GFqo7LaO5CJbYv0Wx2GnUhB3SBzmqoCCCy3FS
WOGO285syc/UPdhMxUuVgSobPrZmWhiuZDtqdBMOW2DkNqwNi2R19GKmrR0+YqY2
fCReNJ1OwCN4RhdUMCv6SUJMfyOiBgnCjTYnLm+qDovzYJZyPz3lFKjFQ5zQgK0z
+6iYSpek0mkTX2DNK88/YYlzV10QDsZrkdXV5aYkGmK6hHnFw/NnBfp+eCH617SW
88m9Sw2L5B53iDh+MKT+6lqQbkDaR5C6H8xsx0E8a+2WtZVQQUa5HVnxcGT+us1b
+JZLKAb2py4oQbOJq8bCu/baNNyXN8qziBJcdcw7IEjCUrXBVcOwejTYR3V2OCMf
58FEbVTkkMooskbxYcyPO+I4UXeV526zx8OiwVtrSG2BLOCULKCiBQ+yAjEJcxoH
2cqpIxatMebjbZKaMXNr1ZmWNVr1/GzBCjKNERQviLrDg7KkUsDMy6MYC5QuoEg7
9+dUjM5ARl2jXn57/NyfZCv5jHhYGll8S2o6XOwdQ8Wxc+mBDsCll9U8LD0j3nuR
NwHzb0uGvsdgFQZ2Zfw/gTmG6R12v0OyzYJ+0uO6zDoqmDZh2Sy7EjxYIc5RoBsb
FBHN3RQY5V21MQk6F8cMOJvdiQZ6vrLypni82r6ndrP1PquJr06YieJm2PYKW+7M
3H3uwZFu15oGFLtRqhSSIMv8Mg/d7WYo1Msnex3UVbaNgPPxFhoam+2jig9V87SK
Ef7FIxR/l98iu1M3TMjGjgvhYh8SCMC5h/gb/0ISc23R/alhKiUNWZDRq9XyFXZ7
QxYJlViKL9Elax5LxV2xCpeHgl6uu/b1pEDd5BsFzgUx+Z6kcAEAzvYSAJpIDffj
QbXl137PyL9kzWfP9OVz2MuGFw4ge5un/Tdaev4mUFa/zYO3gGCoGdkrJLmfUUGO
r3b+I07VColWvWIBYZFm8ZDRt5cMrIxzO5x6wQg028hC+MQo3Q5Os85P7FQ0bXXX
LAt6bHcAjQOS4b17WCaTk+LFDueLryYKsTUFr35T6katEeUpyMK2HPMBjNyKqTFe
9S1UqdVC/egw5QsNiY8P32qjdyKffC7HIeShDGKfwSDMuOeqMwCQwePUcXVBjjK9
uIC9Vz7KhIxFP5LvKsA+cW4lwIm+le9roUqrhx9JomQanDDmO+swY/aXjH9Ab21K
cJ38zrsOyIZxPp2dKKMrqjIXBmu36jmpaBvgGpHoFfXxKy+UKWsTOEZLTn8QZZJQ
Qru6AOkc1Tc8Kqd/gR93l8osJdbVyKwPDiwtuc2FMYg+S+uqNYRCwW7uDJdKeDE9
Idf/a/I5N47LreIvO8ZR8RgpFuyTbucx8WlswyZBumTVfn8gCONjF+M5p29pvhWw
A+3VwZcNh8HZgDigDQLDFzSXmLrcZyAxex5dy2cyKSta9uS2Ox9rJLtkKFPpHSTP
2WeEuSn8X3EtWkY916s2dsYAFUENxWc0Doaq9TKsAGoreR6xMD3skvhGlsFGa7it
QOWj6iwewKvwloCrdPHCtxpUgRubFxLEn1Xy59mn59a5rhlmCpZXZ+HYjjMWyrTd
hwsXT6LlH+LYHm6aoyakyDiz+JcgDNN1DbjM9mA923TIsPBfTk9MCnRKmf/aJeJX
rur5pyugRjrNNByWsuo/eCreYQ8ayBXFhlQlMU30e13w0HBPdjXKzYv9l2eWVWOA
x0/pCj0xYPsQ1fpdbh/SX6K+FdbBVOz/Mw3ffbtHZ/vGbhC+EoPtoAB2AvzjuhCv
zGqacnwCHdnfch10T8XUvN6RK0xU9YLqAKMlHjT1eJ+lu9sJAByERSopbTApoby7
SBpeqoXmwE8o/XVgx+Xj9aX2i0NI4SzvkG9BOzB4zKcWMZtlZ/JonOhewmcDWVg+
Ohw/Bc2rNuS7UojmTZjlHq5ytAXOJCBckpS+1HJlsdYbNONBbMwVpCrqens1hNvP
BR1qDzn5z9v6irsXC1TfeQzmy96Av7ShHwdo9lhOupM82FDQ6MlRqpYh7tT2m+Pw
XO48lR8LOZw+H0/gurxPrrkEl99YIek8OgxOKhtioEIpP+NV72/pRISom5Up4jPn
0yk+2ZgeC9VCnqV2mhDXEoRTSYKQQrp/bkMJcsixf08hjeGnbIQfdJlARNyLfHYI
qsA/J9lmQpkvICHw5R2+wtLd8zCfyBelzOwPqDGJFCwVVWviwlcTjEj5hBmDyS52
d5gMk2rIOYdUVfqhs6aDXf3UAa6nqovd0yf5nYweFN3OVkut4+Kb00GWNM8Mwhfz
ocXJI57mL6gBwkm+7DjqEaTQf4Rz3cXqz2I7x5Zf85ylmYzWth6RBGtT2NfrH126
GxHjMCPw24AkpqJ89eVebLTvkuu+gkwaZjHKcA0td+cBuiaAdUVnGGmgJlxwl4ks
B4PJEHVijYr0+rNxdAHZghOy5W385vgo83/7AtezMN3usfV8imfBlZG0Irj17lLa
XJqpKRHjU6/YPmcrrdgehNFpgpGiTZ+cHeP1XBjDRfkcepmDB2xaQNXmA3OenJvL
aviHdQxw8RGLhqwNSmb/+e+gcWBUPePpF0OLJNay5BANXbR1GZ8d9YWS2Dp19AuL
TScm7ZN4P69e81QqzfueLq7MZ8zDC6dY59NP6ZCWwJ8tqhXAtyuMh7XB39mkYd4b
h0bXaJ/5kYg9ESa0cVLzFE0V7XpIUQxU1Nt5Qg32TxCNK9OytzLFrvZZs72tbb0a
z8OvAKtyXzRuC/0h+8VVbcoZDJwtVdTq8pOHanod1Rw/Y9iqag/yhRWG+MjQbhXM
yG2otuyYpLQGrMU6ReEaCS+6vpZ4dhR9KpWIPx9uVievkGufhx6c6+CPl0plfg9O
gwIyF8s4aer9Glup03BheM+KjI45rM0B1hlB30eZoB2y+F3tALLCaD7LcXYzmt8z
x0Y6SXlo+wS+aeNgpQC/qOQksbgte8xsjMRtWMeZNoieSrkCm0IuXQd6Stvr1AuD
p/rPhAGoOHHYY5663tevTkVH27YO8zNw/UaENVvSKL2ZSxFiHVrU50RFKsJmz/CN
BDXz61HJmZdZ06spjBOndkyeP1qdcgXRBowq/62hV+mcwJC2MGrU8gzHbiES//EQ
Qe2aCkGU1Nut0h2TGuV+s/wkTu/Ej8TaQKlOmA2uP5apS1txZavFPwiU37uiBzCj
j0fQjsZF0Bd8PMnAr7pNrLqHv1kfa4oY4mragUYmb88bOUtQ7i+78W2x7HZ824Kz
dO6vAL97Iubxh5cLiiNCTjBMQ2jHmr2OmjmoWXiwzkhT5LH9tVvJZt8bB3jVK/kI
xZR6Uef1hiuJC5s2FhCRtmzVj0OB37jU87dtQ3/rIX5B95CgdYkR56PQd/tCVKHw
hhqGDwetzpROUEoOoJN+KgkA4eNJaD9DmboOocbe0mT79xIoW3KTqLVdkY4mfSpV
RaSFFlvxrNHi3Iw5Z+Je4YOIDkhu1PU7BayWhLOfNUQosmK2Cp4uQvK+niKCGThW
6vQlSpFTfTg4Y0lvfr1lHwX+k+RmzlAEx7lH+E0zstRN3O2ff+7nJcOk5Yq9lxhM
hM7HvBbuBQebib98ej0CQhiKm5wMpwB245wtaRcTS/jRhKPKw1l0baD8Ne7bEofr
Nh/yod/viw+OjH2GSZzJ2WqKC5GQ4Se5LXbJ1oLGoKOfxdOvIpToxO2I6RrejyGJ
KQPotc8S5Lrf5YlJ4vVCLA2S+NkmPCXplx7oUYphMVjagtaIDPuYmgDL5h5UtN0F
93wwTyIbx2OdPRf2dsteSHekplAattzUImBcgSR7JAwiHzjUQ9sQyI9PJC/8T5Si
Gkdb3N1woaN/C6PV0d57fnd497r26Ygo7RRdmb86NOLHEYA78bVZuOTXjGOps+NY
nQObcxuJMrqNMc9GEzGZt5VSHpDdJAFfsZo0fH8Obkf5o6bat3BM1OYheni42/k8
UUcOTsrDAoGyIh1dQvHqQJHK+fEmTpDS4S2wHKO+x8nDIbqn1i0WCP2m4QSoV5er
X3wZMYp3U0u45aWB+Y2DxdBjHoktUAQ/cZfcCAvEgT4OJYGecl81I+SgCPNzP6gB
JAEWKash7Mrun0msQXvzB0KrCJvzu+ZuuZIb+oQGruV2DuY+/hoBA56y4Q6aHdbq
yBi8l3iCrIS94hgjPEMh19mBN2A5AgLOrCHHA81vR2x2q/gp5rUqXcnEGP8G90mE
6lVAFIZkmvG8RwGYnxagTl4MePFZBqeoo9amB+s9F5nKpPVQ7NwDK5AENLCa7zV3
gKc1ztW8T7Dtylk1dSHdczd2JJ9pDSrkPSmm0UUPo30o4OkCJZB0/5IxjX4tYBWm
CXJ38BDCsEG1zDDJ4JYg+Bdk37bZuL6kiTgmR75xvg3o8H/vqdoLnBGsfSWxJ19B
6ChYnjpzj7OUX6AkxjL5Qt4UeFrrLzoDszrGUUxVC5BDuFqJDaNOx5yHWFm4Osv5
xz7Lf7h2N24S6cFj6uBNvjB0JeSBmzjNAlNB++V7n3FG4l87jogDNMLMURiSQCwf
cJWh7ssWQgohTPuk8qX9i5CwwBpU8sbbmuHRFhOKEo2ujLYJxwAZkPfVvOq7BW9i
viF2eMbARK/mIrmvcQx6FoNr3uilAkzPBC+X6819OwbEuEjiG6cEDEiPaM+XJDWl
GTucScXK5to4k60EYJ54tuCIvHQ6xlfIEsCZx+uwcG71aYk7TCBQqWv60CvnSNF+
UnX8/xSvPbYsn1z8lsGfRLnz0ot1lCLbc2RKZY6GuaURUXeWRahUb1EjmHcmCS3P
sllw12kQACETK6y8I9wiau1ESwdRjkU2G0PEO1Z164LvePS/6kE6z7VoyF3S2a7W
xlCMlRBVCED4owiyeHux0qNe7LQ1/trKpPQIV9/c5gE5beI07lZRAxgb/N3x5RQU
WeGHFZzDH4ac9RRN5Qre7HdjNOD4BobRy2JvrjgPJU0db5Kk2BWgF1zVQALempWB
iDU55LdcaviOsmp1EqPkG0CmQ5+NJXT6SJdBhAWRG77GHhC50yu4cGQFXEjh/zWx
6efsEshptjGa8hwCATIFK+KkVrkzjDsfxXhAat5mgCtyWf4/W+kHVYqhTKAbgs22
oW8Cy0A1K4rJUiZMjcFWbmkh+t/lvfTp7cP7W+rVSUZxvoSWMDECbFSNyutAx/cf
Bz88vAIUHv+IFgZjTsg8wwelmWV52/60+draxwWqk1IC0b2nJxlQkzL7rhnZby0V
/SlDBPi2qIf4YWId/oEKQyJReR6YlxyCmeBm4hD/GdkV3ZtUnGmIYRLg7eqKpE/J
N8SeHgerTBbZc692dGQ/RGK7gAi5P3EltR80yIdtujSTqOfe+d1kwHQSBfRzONpW
qAjvWpfopEeu6jLtucOzgwy5U0bNgC8gQChbBAtgcBF+118hw5xvTjfEW3JGhGBV
AhM8quOytkHUaOUQBtMs4NzTCEqexxbDaRHQzdFiTbaDY2c9XLD13k/gP17UaRqB
2+ldO1Vn0bhM1ZyUlVcfXSqRSqPrv0p9uZ9ZTOPKZuIGiFbBUV9+5BdiCeX8U4bX
CqA7KhC+cQAOz3GDghYHqLuIaQbztOb0A9yT2GKZB2+A5HooB/ujBISE0h+kefJv
l2hbkw8rPo7iMlZWCj36g06F32d/JJalITDIn2RkZZPZMsK87UDWldfjAxejbk1A
X139aVPQUJh1EkVc4wtu8dXhI4bDvicXQ06Iz/VYzrHA2XSGLBj4JzDDLwg2DhQL
6LhWDujfoPO8L8RQXRdyfWBVj80mAlv8q5kDqJnLoPWafGLKHgK24Sah/3+LRgwb
pMjD5lrt1/c3r3VM04W/TWcGwhdZDWne9o9p72euMDnUdElRPTvmI6bUEdgSbIbG
mg+O/KZLtKpnD+0tHaviqYePrOhVx8EtlalhB1O5GFhWbkoV/9ZNk5CRT5KPidrX
/VxzoHcZg3gxXA6Dat/ZyLOpHmSSPTZa2j6AG4DtuZPc8Ackzod0nUHOrgdzfgau
ss7lnhxl/poHilayrqKBUqW/9Nopuw3tYFbj+fw9PgyORsSuMUqosIFGqXab6QQ0
fcGQo01jkRf7D6+nlM0w2Zpoy9VHby9lkULaEED1ap8JPsudcIFhEsBZ+dujANkU
+ASWTNUyqRc0ehrZ2bAgcz2RjIf7tZPw4EJ3OhVtJhOA6yovaPve26g36IT8Un3B
Vtbvxlqs/i+HR/eVB9vdzSuLtKcuzyX0jP2n+5/dKNfZyhlyEea45aJGYaPaayqX
Pt19fzfRdHjwxnzXohuMhOYMiVZVxqT/IQy3gtb1XGKJ68CVkd/TVQpNtQmbvCkh
Bw1t/7jgyqTWWUkboBTob21Gh92vzOHdOnS87JX3tWdoaTVPiwv9blLkeW3BbNP2
qcRkw2W19Wn5oOuXs5ckJ/VJvKRmNA/0yGcw7SfkCS5OKsfov2GFsgXy39YK2qVq
a6rEQ7ryIZNcreilVkuZuGJ4uwyrRySsyhJsB4XPN3RQZ57kYUjHYZUt4dVSmyH/
SMXMT5VWrJlFPVNNMid+u7XnxUCShwJIKKIfANWH5WCo4gJYwZK87tygpsgdN0vv
H6dgN5z7269QGuBc/MHyTjSMz1eTNei1O+rsOaBC4N1YVTk3sHf6EaHeffkBXqXT
OjIDNiv/PzIhTgUD9uNtKsuGlN10zbq4/DnGcKBAJILjW2pvq6VHdDr3q8526299
dMtxRaPx9CzaU8IAx45s6jVJ7aJZ6F7GMie2k9Dy0I6swWwxgskfeKppjSgOAh2O
4AfAGi1DPxT7Zq+rhfZQmvOWRREsd/vUWMv7T0qmIewbR7SV16VUZ+P9I5awzdU7
TuNxIxF3n+fzG4TTHYj9f8CnSbOYMwg6OEeGY6VYW6UF/AaEFUdNwWD3kaLvBgAV
/i3657eRHBlfJ3ErPGNNN7cgyWyx7rYQRoURnqx0dduRiE2mQd8YHj4c/DAYVsvi
6mEGxI/88fuexrqDUW2kbm/ROH0s9zIxMu5vjPH6X0kT5gVZRRfC/SrXVNtxVnaD
uk0iKvhIA0IHI6qMSD+CShj81x7RftjQPDdpjn9cEdSO7vrAr0V9PqLOwD2jjRSn
p2um4SNUZoXbwZ3UHiFLRKIQ4nFcnc51ZsWKbmg4h4x9xVODoODy7Q7esErIr8Ty
bMyI12c1VUU/dNF+6mRqMLHrPkIzVw76Poxwu7zRTEXO2GbAazXBjHMR2mq1+889
96Fiaav1+GCHjfwtNVN33LQfVo6y9lbLNt6pLT6MoaagIUtNzt3bylC4x986z4/7
9b/meDKH7iYVGSdiZWE32TrqVybx0Chvl1zPJd55xrsyb8L2dkY9Cf2aW98Mwduy
fmnhJGtJGLxOFjY50inaORPnZkVi5QH6rzlEgp2MLDPyx2QeX//hvFWHV0AE0B0z
DYPv5c0TYxgNu/E+hVIFe3Lgp7hpn96c03Ixb9yIuRFuudgv0WGwPuL/ZPQmxZ63
FzOMfZgVX0W/h+J9XfkzzD1jNdpZCcY/u2PeGMx3LRxnQMREVnWX9l/YMpuVonAs
S4h+bg8SucbVQokWVrmO1ZXuUxlGJ9VgZBRyAYyO2ypOCQaVnwpDLjQ9SvI3oy9E
Qqj37jHnClVvNY414m1Cg1MyvTROcCj5asioZcDd98+6h1Z6HUWGdCr/ud6mk1/8
Mtu3YwZG40ruwn3lnOGShqIQzOJCHM00zgDoaJQvTzZ69kVRpUgMPJ/MCdKQPK2m
js68EfbUm4a7qXgQyrSo9Hvt47HknA4UcB56PDtA1ItTxJSfVDmlTJrWCv4AMlhB
05Et8aqAyaMS3ceFaXVibTIo+JpTWF50R61uq2ECL3EN7GlW78KsTudyaRMPDosI
onzDu2Rynhau6E7/XzvLBHNFAM5908lNMeXbjBp/VTV0CsvpZjeShaOrOisLev5B
C+uIvj1yrXKURtMr9thBwRcxnW/duMP5w6SxyTt1ZkVPSxJ6QoRqqc2lQ6NeySzF
OKoj3pWsEB9x1F7FKDipSbZgkBLHbInYeSciFU638D2CU3JiYjjv7yLOcfIYZhSf
0uybvPD6EHDe5RKTjxTEkjr9ENnLLVvbYWtsHtFq1UBunkkOBWVwh2G3Z3iXyFy6
RdbLeJ7+bJD/ZKSvyMXxrAEtXbB9jA3nKmBS4va+9b1R9SSJp4PHFijDtlV2xrY6
6K7LL4bag1azypp1vEOmn6yS7YEPIK7i5vXEmb3qgqmX8TaiLYh6BOktabf4Uzoe
uV0dw6pUBZmIOq1rg6dIaaM+TH2vaignilX1cO8L15tkZGgg6B867HbVukZWbfeZ
xI/sOFMhQc/8vwL7zBXiJQHMyDgNA0JSE9+MkLHNkFX7HHZ15Ximm7bzvfb9Pu/z
nCuUUtRrdbYJJAzyUzvHmLTiMB2z8Y6NJO0W3BNHWO5qeBSMTySblKbxBe0gF1fj
o9JLG4AE2agLcCS7uiRGsTFaTjQHrb7d2I9sZB1j5/eS8Q4Cifl2849JzL3xdYHQ
uO5J50Mw7QZpEHz80y2dQjJsfobPJ/R7Mk3CJ9U+bKHkdy6RREk0pJWHdq5ClgMW
C3A6HEHrEoq9NCJkQOH7cIWi+Nnbbu3YcsOlzVEPOHLPSRscDNJS7rJzodqbemvQ
OR9p/vsowh9n7vZ+kCiYZAsdTu6juRh70k1MKGb1LTSNDLm4eKwDVSCHwLHClR87
KV7WW2o8esQquYIDZgYkgUff5q2VCHI02DkjPMbyHMzeq6VwPxjd+I8yW0WkEijY
CIPnMS3yioYcECMtMAQ4kRjoEqCWCrvsoEq2o3hb3mBhaSlzLVtGFfEvCIQ/0Go+
eNCA+b8PkG8d8ho8JD4vZuHZqjjp9BfbEuhiXxbafM0ObWKSS6T7V3/mdDbXIA9m
vfwTJoiRzGEDZ/dIpAUhMXzZHk1k+k3dCmWw0ZKUNZerPIzIr598scqxTc+Tar3H
9bwoCgtxRVV3u8kfKBHbdjCEXiMx1G4xLlh4JgiAjwQz1jUsniNxLVsplqEmVdRf
V0raxcvewkLU+xguAF0rRaLtYGvUkqFZ0b6CaU/vfNbvr3rxZgKEYVVBqrfEV3Os
dAB6OANStRTkpVc68GFRDu3fWjQZTIIwqYWIJ4kZQFiA/102fQ+HMtx5jOx8D//N
MR09EjML1YtT2IYoNxtAV0dDLNPOpXXHW3ejqkNd6tVkW8kLEtkURBwyxzAQFPcr
W6BjADFaRAo066az0dnDI50YqmbqH5daIpKzOG4ML7Eh6pN2LnBwdtOo3twnWgFj
tLG9QPAtFjPDgOStm4Jf7i52uuoX+S/FC553c+AlzdzJeZe9V9e0CWWNGvNdXCfF
xoxaGQXOD4xk29/3C9gG2nR0VEisPtdz4Ngd0tLVW74v1V7Srv85qW7FJBajLeZq
5euOwg9oVevx63Xthd9IBQLuv3mYYQx8juVqonLHXByPzk9kYsJ7Gb3DUl+xWSUB
l7fpLCqQh/qUAvtM55EhdVQTI8ieqTmZwNujjgKQ1XWhxWVcP5Ff3tr46M1UYwFE
7ql/csfh0pTMTPwNoMB/83U+UH/MUhdo088jmDruJWhxFlQQl13fSVeXYz6y8Y+8
56a8uQKBtetrG2wYqo9BtYIOppXHUFAfue8s6G8qvYp36YWPPY4hE0EfeLjIFYco
H173kETDmpUgT76wfVs0BUtkti5PrgpUfdg8U9Ak5hIBdlAaPuvWRojv/4etOBhf
JjXZsVTlRsOXZ0uzTvYGyL+3Sm95kW5R01uBSTYzlW/t90hJ+0nFTa5fKwvXApCD
TIwB90k3f4ZNOQEwRNSVQnmuMNozDobI7xAnmCVsL7VdHUy77w3aXPFWOA55HENL
5boxxp67BGK+20hHXC4BE/bk+EQ4z+kMaoB+GvT9uIOfpV5IViGzl9S+D274oi0n
09KyaS3ezfBVL3jCeymXa/VAG7JVS+HcSK7MxG0uiW02jAY/jiTw056z2lSEjbG/
5qfDTj8HorojI23+HkX6LAa7yKbityTn6Q9hkPdrFqVnDp8ldP992eFCIhe8JDOf
rBOB8i/IbpGZhrX9fKq4QxwIZ3vfFfVDMOpZrgCmwlA+636UmV1EJzTvF6So3J3T
3WSc3uGdXQNgKOLtzbLv7+kAGkP7/zWzk7uZfg6z7a/jTxYmRqh01cYLjMazk7FT
czwtA6boVbSBO+0b4d/J+5Gb4p1xVwrwOyUqHfIHUf4McAwwlBrGD94GqhqgPLy5
Ol0n9nJqIr/UP9t0hI77uOrfPeAhBm4vX/I0vY4zunMpw3PVAsN3mJHnLszsTOR4
4RBp168iwB6SsSHAUgX55mRnGltCAXVIva/6OuShSi3YJCrcFSpBkRmr/v60ZTYo
ZVK2iWq+cNkq0M4fBcMPtpffiwr97GRpgK3f9aH+rljczz5caBJRK4vGzzlcCdOW
yibOomGjfAGwpmFgEayisg3QeCC0Yk++cwySeUQ/YRKJDHhQ5WYQTYqkGZv/FDkg
gqAe2J4qVNLaFyuU4C+emOL0diLtSKrDM1qWjcOzWcLgjSGm9YUrVYMeulKE2Z1g
ZLBqw+/F3JrSa0t0v/vkzBbl8YKRa6xf/8CnM05CxJ34YljXH1s/8ZODVtJIofWE
yEKTp/48jdETCzU4qgtcy4NZTPdDgWECd0j0D3C5o3eBbDn1cBHACuEHAwFg9QNS
i39uq9AhcviArEjjtF/6uqTJAuX3jTdaGJ1uDqwI6vSkGWoEL/sBDDKSHMR0CRdn
SRrB/pOkryRJ/trkeX7fz7t6tdRrnv23R4w9NXkr5ykrW5kiq8H8cLAHKdF3zZUp
celEUZ+2Hj49bJ/Ex9CYFqCjNmOiIPLMm54s2h3c5bhi0/YnaT9Ra9Y8refJ0Vql
tiq28mFIo15eori/BrsKjgENJboV+tvR/85ZOaKmyYQiYIN21+lxNVcHAZ3WDj3i
wlq06IqVmph3XblX2qJrOgQDPiSOo3NmBKOP2AOXAG6H9SfSbMYEZU+umw1vr5Nw
o5ny77fknw0tW8sENRmNZ1KlzaIxCHd22z7uHETB6WHPHaHYeJe0CSjYrYkSRodB
R7Ktx0GIgoU8YFHT5RwLR9V2mJpPBJ9mdWYE43DXOVhP0Fsq+hfSboMlpgjLPsl8
lHyJA4u0N87S3yjRVSPnM+6BONSbHxP3fqGMEYRSHhhczjGMzZ0sEOm17uGPVRHj
fKYLI6rNlVyVcmHDAbeExalRPzgjPAT1WLnRNnqhMzAMSx4c4oahpyZJMp+PL0H6
Dt5tXUQoxMVGPSoRkg+Gfl53hYHMBiPYzo9injDYw5Kbmw73EMioxKar/HBZ9iCT
ZSoK1Jd2AaqelHyhrDY/RwtU4JBK0Q/0ePSgjfjJLRz5htxytAwfU2VUq6hQbTKu
ETqa7LLtCAlt0LrUUQ/z7WDRR1fZmrie4GDovYYFKJoU+z8dW00QCZvtKQ4WTF3x
EItbX47rVrw5Eg811g2VyzDEZUfOGniBoCF6EIL4cg2jjfSLLnWOXShLsMbQ7GFN
5ZquKhKb6IwE6pk2aLzZDccTIcoqTmigPuhJnZW/j3/0xOngZeuzd8GPmQHrAd2/
h7EleixgX4c93PJSDRJI9bGw/SIybxbBzuMb+kN0FNenn/hep4yu1sRrBgOIOrRm
xrKLJQBU0lF4z3bQ2fwEEVFsvw4wo1z/xxPJJ3UfT1IbtXrRYy3I2qVEz/qmczJY
anAcXf//W8/5KXkj+mCbaEUcdSpKn0sEa/UMkH9lodJpWzNE9CyvtvdgaFigQsL2
3r/uT1WgOz2ntnctHydmEg0RZEIRybxS8RnwHRm+Jdt9rjo/sciBs3/0By2XFH5L
Ft5iSki8a/n7WGWSlItH+gXVghitSo3AnvQu9cu6eErLxkG7Qhipnqpb45E9uPbo
t9+0QDdx0Zli0k+/LzEiMsWaTSdsuQfPqyGtrgb4Y0NYasR/It4RrpvFZypAJeYm
IzZY/nRasQ/xTsKA0cKs4iolpF691ewHC+ISSzplZSOlARXrifCpaxGaom38No8S
zQi85ZQVF6GVDNVpDYrMpllLqZUkDCPFm1rH6pScIEVH7aZTd85HBQUHjEpR2QLU
M8/yhWy2hKXCHROY8qlrCdc1MVG6DWXOhxuXnt3eNPL1X+pRZ4mxpFi4XlCNwDAr
6YVCjQ9vbTXmSVYVrlO2963EjIrwHpxhtAKWJYYwQ3t8tsqb9PcgP4gLXMY3OBus
kpjL+6sXmKFuJSX7khMru3H8KjYoJ7n3d2L+k89d09aXISOQBu4fzLjD9EWT6kzq
0OKMEU5JGm1rGVgNEyhCPwFyuqIdOmr4KKXW4AbcSkhp7NBFammuKoVwKMapkvQ6
WjOLEQvCMLMy9gqQ1EqDs2W4OGxTr66sgshmNhVZK287eW/r4b/Rf7IuzKkTXw93
9IlzhJYQsGXwPMDMHYLE2Gwze2CUO1pu7HJRtpOnEW6Byd8o78Htvg0CdbglKg65
gd9eZ2LbrqUzO80r1bbjy0cGReAiI2XhO588fWrJR+KOeNRONR+Jhpvtw6nQOcdl
Ffn87Xjfskt69Awu6aj9Rfvm2AVAEGOeGbR2/J2KnNvi+ERhyuFRxcsIysKBgAAf
39GFBQViNlLIHbMWabdkjz6cjiSxLCVmISEvSc1jxVzUzomojpm/6Ns4V1rtTmy7
unyY7EZ4mqEBfsOD7ygV5Vq2LGsfyWgsArTd8PLkngWZ7LUfcGk82A9HrnFGEUW6
vwLH1VfSsSfep88FXhnPkR3ToNnfNZqZ8DeZLY0PE+hXF2DncXumMlMvEP989E89
IpFJ2BrZ/vIFgWJrCJLBRam1ErSnCuucAgeKpvTuGGoFZ4c3ec+gjAbx+4/O/NhE
HJKCpTy7jyQbHm4J1CD0gRRGnGV40BY/O2JFhQL/5Op/e5HGLw0rUALZjNMzOM7F
BP1Hb7+F1o0bkhe7f2LXojKRzRjHxzCzbpRpoYtfBL2le9exqDNZlE/fMZFOviAB
llBvhNvy3b2Jn7jEqNcq9NIjsFHL2S5CGPwhh3REzirMur8Hq3cRze/0Es0wHTMx
4seUJJ9RUwKjv/XjOS6N+lENC0yf3oafkThU6XqB6gFBL8Z7phT7QykQ4o4a+GUQ
5Fq75qYUcjJH1Wv3tFJzA/2n3SBrgU2IsrGHgzZsuFo7mZgEbLFD6ct7uNN/hpp2
I/4ss9AW9Miqdejm+RMYwQ+BEU+lDgmvZBs1tDCqCHfR5QqpZJKyA4MXEQBhzUKe
wCPlrZkwEPN4OVMw7xClPL3luVOf/seuoJd0UXgUKiVf/UkMvZK0PfIkebt1VkTN
Loi3+27SiKn5efwoFZKMeyYvp4Wd2/irTCwvcYfq6azeE4Efe32q+N49cVw8yW/K
yPVW2CK5KEsxGuOK/kJfZcOMf706uiCHn/nXGAYEW1Aqw2OinU/GgfR1jU+cxWMW
KjLTgtu+e2Md6gZp/CAPF+AH3E1j3bNzLm9XxrJ1odmOvqK29+6AFh3nPuUN/7Wm
Iq2YasFO+iu0Wf/TG+83jhnYsrv6CNO/Re3iNU1uR8uYypKUG86Ci0n6DlJGgHAD
mti3+mL2zPeVfT9kQLicGZjZ8zmzI/KcJpqEumR3ODejtwcNCvnEfqSseF06Xbmd
fRJ9aRR1cQhR/uwq7zkioiL24CNJiSxCiGyBSGuPLB7aq4yYw4NwQAIil8nrmeNz
b3l6cU01bdo91OXlTgGJmskhGvFCN5oCnneN/kchRHSUhQY/YnLgR1cfz6PVMZLS
9bx4HbZ7C6Pj4ycuqzccW/rGNe5gOv0hftWpmzCXuItgPAppkN32FMGPfup95yKv
NAeOjpc0T+A7KprEqfPi0zB6vB7NJPTawIRKTit6yMUjNCMjKQ2lt5XIARyhnft3
4duk2b75Nq1WjRSmFEUAHsk1XAIFnykvYS7Gc/9IZBsABHiA/XvVFEdcmm6I3vAM
ZpQHAQMu/11SlDA3mo4YTHsBZP0pg/W0kVC1xmPi+JaAclN7NoIPdekj/8KOKrrz
nxrwhP4XmTkIcK6p56JvV4nnFQkgAZWzYc/rKD/kK4MBRpmf4zzncg6eVMhd8BDb
B2LrmGT/CLvHSiIpI4asPzgRYPcsNl/QEsyweMwW/ijDLmk0Uf79pUIlTVVLd5J4
JiyH7ACf4qSJG81yih8ykbEfGyUyqtOQgtztsblDdFvz9qW9MUE4K7htnkGmq0wT
Y0o2OnOQmUi1JN82bQTkOuHVaDtLSH8C4hElvkiQQyZ3ccqzxlhGnMTJ95K2bID0
pc+QMSoVs2TqqDP0gn595VM42NlvoJNztBHlDgaHrHTybYK3bKVbzUpDCyKEvkNf
dNofG4YF8pY65Vi5ZJSGQFdw7dxEy2SGeNdKMR1yjVpWjrzMNUA3Tv2YUpVrTHGr
lR3GAZeDUtMoZPV+QDYXmcScDics7s9c0JlU9zQ0/GV9yBS3Wor+SLMz1un7kUkC
4tBq13nH1nJ71CRPIwT0Uig8zF8ZjFes27wRGjBAT1bx77m7eqcUabs/L2YSL3cF
v8nD74t4jHzXIo6/s4Aq0P/TpAORFfx+TIjXNCQITGv8hqiF2NH4NH9x7gJ65UjA
LMnYNLnBolUuARq8wYAMmQUo9Jn6mbP6RFaJhNlPz98trxI2LpmY4X8SkbkuA2wz
+TWsQB+5hfO2qLh1eZh0NZ5L5o2oct28INLj+DZw1y/QiJS8n64FXkd1abQ3iT0U
GdEbyVJjuwbjlsnnzcJHJ4fTNgDDsFcPbvaE16OM0nJJubDZoEcFYtFjJAMFLAtW
29T8LC1aTnPxCeLVZxIxubeZtV/Mg+xd1u9Be1q8AD2jLYiIwuO8ZUJ06AD9pPRL
BV6TgIPLY5rVUiWCQx6ZhLYCIUDcmJqShEo9FTMvtSmIgfy1LjSSErHKofk4OdT+
TgxdLxWQ2MAFsuDV+w7ADRmzSkvvt3yW2/mAhC6AEfxq7zXY3RwifATtw1lVTMMT
JEStI8EClM9sBRxAQrfJqNVdsyGSxCFNWP1BHb+bh1UYORSj3sGMG8zCAyovUEUp
dAazWRu3YhgyVAC6M3ZYFw99+pNgOW5xFF2p8UfJSEHOIigFgL2w9d03kLVlNV3u
e0PDuWyxYB8jH1undcVbR0dYwEMlLGRu8qcvRKTChGA6TuRNemGp6mgSeELYkdFj
gQ+8S/BZNzEkk6UL8wOXHdUsUlJdN7b+nm6cFre31uVfXdhnB6LYWVo55Dc0Jkj3
YLEA9XeRRJP4htj6sooqelPwr+pQrlJ7NrGJh4pBNyscLBMk7RZuq6WPp882AVd/
5n/mvtKNsQC7dtMA4MYvzB3/o9fDOsUJI5hAftbSTozt+nh5/uWupq+NWEBNxqgB
mbY1h1rLskwBeqDArYINbXluscpt9QCMt120pWQqli1ZvIj5jop+Og7XID0dQEyM
JXS7CIPl1A1GoCYg7bTfjvQxM1Q4spnx1b8WhdOQKj8gDuQgl4dMIVCLCxSJTOqQ
MKiJfq7Sosm1pWBGHGosyCDhLszbKIMp92NZT/cyggebeVq1yQRUiNSQexhMqTRt
JlxhzmZIGgoYLMTyofOMTetpTrUrlEBZL0ld+O+OAjlWgXN8ziehXXMgM6y/Dj+t
8UtuFBOKdFdUr74Yd6C03Zzr2Jsk06HChJZwTOm4vzw1UGBfdbi2fPMP0Uo5LWRd
XfKBxIvwHcYkmOaKekPnTXTCEQ3YLZ/AOfZzxAxj7hJTZuGWVtyE9DYxl2ag5WmL
zO+/VYkaAx3SNHAmPoG1JI2K9gUBxAwZeZHfQpGhRZi2iWwndMsIlc96ZhSV5uJ2
hVVQY9bJ6l7o3NaOzmZH/ti5IrVCxyx86rSHN88h+GNDSK0eE7Ou5LBdJQzMW+Hi
qG8Ll1RRNbayIQWk2yMsZoqC+Y93FetBkbMVacck/xazh5R7lMmV4iR+vT9cv2vp
LpbHVSnliEDv1oIYBfSwRrcDkYRwue0JaBBgTxpd7mTeFZCgg+g2tn+5Z1csSKCy
RTw9+ctV7OPExGA/q/YC8t84I30JxYeVbxtXjmjBkcjfOWmi/VzWJe7PztQZgwzj
G2bwK8fwGAm99n+WKM18BAf3CN3HIqBuPX0WnnJ98mObBtUseV8QE5a84fNvxUng
zM+xkKTnuSjj3r0fZ0da6597JsRwzeK5Cc/gB3dIkwjf0tMKlocNA+jGykYgrYJk
hiqeaW215fbypJmx2yTCYEGLq0AbMfsc6Kk3+b6+1/YyZyGycQNsGKy6/mFsLBrF
bYLHNmf9Z77Cfz3XRjsp/gY59gIb3+oXmYvhUb1ZU4+Pm5DR6SzekmA/c44Zq701
PFvnYk5FoOcM7kvGrlFW2SbtDqxBcGlq1gcUBdGjaFvKpgoWpKe2nixUN0mMm235
a30Fd9MOENxEG3LH4EdqGo4or5TK+/wVPh5/l7cbtgBXeBCxq6qoSDrI6jRzPAn3
rleZ9pHkujvyANx+1fsmzQq64DZGpEZxPobdih2h6P7FZYSHsJ0IUU4QjekLbZiG
QxxEgOoZngkszPAp1Ce/ioj/yws/DhyPbqspmq7KhKw7cJnuxghpNmBOSmunIBXJ
uHE+A//KWhXkBtdvKjPIrpSNBKwzt4TY6cLUANlZhFMUfPq0tQGVHJO8ENSHKaVr
vdefKMNIyiNuN4xDl3Nd0E3lut+PxITJAsZ/QGnt448VobgCuoa14VH0VDCw5g8x
dMK2BtPdWDRYQv5HQWHNuX2LUQ3GactqiRMzSikZOgXv9tI4nFUyu9Kec21S8s75
Raj0DZT1GBhaORgyzcX+2nWT+H7EBT4WK2Zus6hVVS4knax+6vxZcWPNeiGHub9Z
D8uUdthO02zwcnfmsrnCbC+Yggq7TBgU0ZXn2B4op8dNwDSj1K0xrTD1YV5XkPu4
lp+oKxu1tMuyuxh2pJcOknc551Zl8X7OwGY4Ti+hahFFrae9U1cYBrWh3pfiBWa2
92qG70WMcsXb67+7tcsDLmMuSuB/Evp9vveSAIzKROj4m0iX6m1lvLK+dXWZEPNN
ueuBXoK0fgaTPYpWqMz6Yu1KZ7DL8dWFbLTMuUZ3lnkxrKjEosK2HCtjavA0CT6S
OhTfVmxsbCiSYCiOrob86/5D8At1VkEqNz6GFg9o09QPfhLtegGAQgX83Kngwl7W
TIWukZAden8n6ohr1s8amk5xIVjuu4wVHOFiVDcRHtl2KRz3em5HmMmzoz25P7u/
NjELWha7FuaJEt2KyQN9FFEN+WIWUZw+Gx52mC+VO3+4s2ZwWIoZPXpu56pBDUOS
SHLcxdz8Ox02LPAo7IlOfTZXVuMjt9qZZVggtIMMcFEsEzhYFC4GPELlmqRurZxn
5ziIeQfsXnKsM3ZBl0oiGncJ1vRy7g7w4vyNxp7hKH0LSz2Eq5QQzNqjewbSE2vJ
ExVEGk95TeqiqYNABWZXSy9f0vLqqArRd3yCll3F/TXE2tQ9uhYfTeSUK6qfxdK9
UdNOlGvjSaQxABhX0dORwlRmv6MayFECEYNAlfTc7+ffXtXC/2tNC6ocpjhmUp11
+VrpRGsX6cN9ebqvg1TFtmF/0ijg6pk/08+0ljlfwlL9TkfoilJFFD4gPcPhdyD8
LVjcEl82X3GQBjndQuzR3uNkHZYBBYokonrdQ3V0ImC4pD7ZlBbqlW/lRYPq2B32
Q+IFS2OsgK89MJ4L4NgZmIgbMYd2k7I1djGk0s+PiETRccfAI5fGglV0UwYtoRyd
uEQ5k0lcJfK/fDRQ9hHYMiTrwbZBk/iokn3BkzEJOFEKt05pwooEBG77M2zAsvrb
sD2MGWDmK8Aa1xFBCPgoUTFHACrsvG+zVksCI8WQ5j4pACyEHzTCasjF6fpvYDmN
u0xj9mB6mTs95RlsEvLFp07XxxGIFCwn1B6vHCAXLzP2CwOW+i2u1Nfu6nc/CTd6
B+9PUflyMqL82HOLw1lVvyTYqkRVyfUsIzJ4JzYE9nml5qG8434sKj40KnJ7yYC0
XxIl580VFUOQl00C71iQFUmUaR9n6000oSkxZaHA/M7uQX7l25tCMWVmUh7cYv9r
7rcYpR7cuV10H5hAGdDRy0wzOAjZR4Yr4kNsj3Rt5v0T9SgML1w4Yd1MSQC/NeOT
xW1Zqy/YypTJipdnbdhQZZMQJ6kNDNDaZYrHmTHj9haUkNb4I59/wa+Xic/0alpm
eHtmNbGlBSJjhGHoycNzpaZiQKuDaNWzU1t+0Asep+VcO1A481wa+EXVMSjCCxQ2
YUzPjQ/EbjrSkoLMFSDajwE/nehbAUAJkgfGYrO0RX9/P1UA382krWONp8zxowWx
abz2beFgcwYuzvc8QZHPVc4bqAnECe4bjLul4LAE3lZoSvZTC5bl/0t/T5d8Ipky
x9kHYhq3XUlvmk4WMsYIyNg+Gyyr6zuZkHQBzMGfeWQo8dcGAR0ekqOZ9fFZCPD4
a0Jg13CPDXL8eX22a4sy4JxdjjeGMysCqH6egeYAkOdMYS5b4I1KIupBEZbY4nN+
9s89yFY26mzgiyXKeZ8a2UcTx93jnJpjEhz51f3UmQGUmU4LjrXrquIAErUqNjqg
Bm7gzks9vvfTIYdCDsy1uxWk4c29bfv+/O0ycVVdRkUQkR/0ko6d6+cFUNNK+3cV
Aa2ZuAhY83uQH4Mes2gb3ms+KqvDTGcgT99/jvs6F9vWSbqz/qoMpgXid9q7DQqo
ciUH0n5nI2VuoKJn04ujP+s6A/lohEB/PVAfE2SI95MjFV0tF8xRhY+hcLwO6rAh
lleYzHVwDVqVmlbS6C6IA7SYV8NvZd77CdmGhKeMk72P6DKWt8hD/tQ+sr/FUUkI
kNWaHA6W4b/ce25/hy3FB99gYFJIS9LSdUmGi1mfIJpej/14dQYmRGurvr1If0aS
cl/+7/EOyE8wL15V5AIKZ4D9NdZ9AramcpN/sgK41PLxYQQRZvnVViKhPaIyhLl8
cmsrSag7Vp9xwN44n3kU4HzIX9VeaDPWbvQ2R9EKOQpk4OXPJzRrD83QtnBtDo0+
wMhxH2qP255Lxfuk5f2IVjo2oljgeiqHfHVSG3yhujFaA4a/AW53mrWDb+Ns505K
JTQnkknEEhaREqvAjir9o2hOgPVf83neRp3bf3TzUxSB1VOZyeUGM+IaOSUL4v7i
5G6118HHiWr7uEJMPCRhJaftO5SrEZxZuwZFjw4Cinbngj1Jhrcd/ruET+UAeAmb
IsF6o4Vxm26NmFG26MiFhLXjd12qCf5pUY9OLHI7HJxta125c/eCdOchxfzJITY8
1lqPhfoU2cgWlZDaF3Vy5DPtUYaieKSt6Gi7EYDipFvaBHzOWmtX7q4CkQfRLczw
BnaGL6mKilUGRZ7aNm+BnfYOe+SGSz0NrWqfelSXTQOPKlZPD92qtf1iE5lI7CGm
vkpg0g5+HBwi3Sg6ousFIqzaFWxegjRjvt6ws8WHS4Y931dDr/rWa5BAyAibWBdd
ivOeo3T/VI4AU+k2sex/qCZgHQMTvLnbBbBKFQgRgHryJpUSDD35NLDIyRegi8Ij
ZN2BzC5rbuGUSybwrbFW+D5W0J9p6hTTmhYZHVrOSPoT8LwO4Z49Xi6sIy/i4qok
0ioGH27TOCGRyfx7DI/KJ9N0B0jLh3+EKoTfk+mBHzajdpMVq4pYAQisY8Tns2fw
elPBXjfxctXjWj/3Bbkx+N39AdX9z64BAV4Gjg2572u/HFf7lGccEQ7julR29JSI
YziQlL6HvldqhUDLT88bUY75zL7MnLpKpDKIJgdQI0ViR8lSHnC3VK1OATKh4XD0
GTiRtBB8Hr/3b69kiM5qGWC3S3XI+kW2fdce0dKxPZM6CE2eM0YCEaijmBXokGxH
vZPoWZhBabOVlCsyLW5qiOqxli8MkRi/nJP5bgim7Pp0nLAffrYZxhlWd5dS7cPf
ovwpxoFjJQOszfKqzOzE+xKvQc7igCFd4Lh9gAVkjfuy9PhIS2KxJU1Q7g5UPnDb
/IVrajn82oZ9gKrHBLReoMRF0F2eiI5U/1eImuakVD0TY7876UAWMCPCzxp3m8jH
2HYYd5EPHFtfVNCzRoBvTW/HFpvy5taByNO7eBgz1hLJS6V1ZlJekBL78Skjxda7
vlF/0uGuOYZlORRGpfnXuTEyc9e49eTPXBXTUCrN0TUxWDLEeIZdbcAlThwT8LfI
/9ngkvXJJjo/TqC2mkHqUep03n1QPKWgXv8S3b2No+3UqoWt1MWw5YKHJv8aINBo
2sP3mRowNe4gudLdUeEOHDLvJZXJutY4Glp9NQlB3oukhl3CASfUlubqFYhqDY1M
eZHY8YyF88E65Df3gFuCg05VbluXXMJz4K2IBBTpg1veHvne14NRi3RWBlYRKm8Z
d30kVRwo1MzWPU6r04A+k3ounSi5UdzgIiQJMNCWO9vMDoj/Xw4qzQ3EhcFmGgDC
TSeyWC7DXQeLcDeCqICgYtJvLgZ/YjdpHIA9CS4f3GCagv4Y+U5IGncT/9NvuZWK
PBU17jY0RjfyAV59sMGoUSuffdGEx2q07EIkQg8rVOHEKyoVxHNvm/lUoXZ5O1Lz
2SOhBZkPCI00lZwKKhoJowiP+TFswupcehlm+pvi2GoIVrBi5ruHa9M+oBuFgFeF
+cmr+xM6QBhWDVmJDASj1e1MW+u9ZIP/G5hC1IbnooV7KeCzN7W2a1ewJ6zDbepD
i6PcaTh0lZW24DMEwFo9yYaWerGLYvj85udnSjN8i63ISOrU5G3bvmGy2byV6qws
0IhXbDo/nkbGX3u94DOTvw0gql5CH4oUulnGDPj1y5PPeu3ijn/Sqv44j7uiRWOG
oT7Wmxu950ezvfPZBF8H3B2I9/+9qOK0/zo2uKDvHX/nrFO/mDgJPo6c9NzcwgZB
Qq3IBxooTKP88cgNVFZ9KKX7QzFbxxR4lq51QSEGram1mQWAxjZuBk2LMNej0h9a
hUu3oZxjXDQqC+arbLAGO7cBFWOBrOCDAgCbgreb2238UEQj4OeCQHQKt3Onr25y
YPiVsjwFCyq7HESfGJZgVPvmMPjN8f3vR/fiNtdpg3Or3zJFw6SPDBgKVPkjvEoj
GlvMHeMEFQbfC5W/8xVMUgFi/ohN4oxmY7dJ8An2BHX+58qkd4aOsFtNkfhO85tL
bMlZ0yMqC9Wrl3YDoekTlLRPXRKbQJj6r/Dq+UvJVVjMA1vTZ/pLUkNXcvY0XcfW
2cMejJ+6dTd+D9DssqOZVSNyGyjqS8cktxf01IQpkAFxPU2iy/STvpSQsLaTLw4c
IdAHvKRElRAySGBDt6MJrglbiimcIVYAc46WAfYKJbUfb7vRRe/XTlx4h4kII9Bf
45Xgm/tD4yDv/M0nd8rSBJdZwjtCelRX8fGZumLBhJc5AweTreVjhMmbmzzQpON0
GKZzdG2xqaPMF5269j5/lU/nKS1mNPzHiJNv77ILjEYd057jsK59Px0dlrBZ0/Dy
w09K3yulGjDTDdRRmzg8pTM3UbNVRwXnbRJ2QyA9txVi795L05/AZSPv2hvm0zdq
ZFHZWWk6v6U0te6ydUiDWVfb2SlW1Nc0WTSRcaaXTogWbSfa7Ubte23Jt0BPoTNw
A8r5JlOos1nETVeteRLULwO/xQ68+zvzvl2WaPgM+EHTXErlXOzTM8uLIiEX34Ij
p1ft2sANTlv7pY589jM9qzd60ihe5iN+e4voJ7pHFoA3iu5P4HNmxODGaesRRPrn
yFU/0pM0q2R0HtgWI3Wh6DZ87RHiNxXoBSmtel4XaE4EDucCgRCNAfknudT+3OF7
iSiTudjgmt0SgAnNHFukZYhXg1fXgq59YGIvXM1zRYIHgidSmw+t68mJwSjBvfIb
irME7FG2rnsd4r02Y8K1FBgS3GbVGCRzlrnFw/nuXveq1wee+IN2mB2lGtT2zHyn
Dq06CDZJsHgDD/+Td282dowuLufFlvUZRvAN1RE0yvvh2hBW8HMGq3NV2ulG3YaG
xaRPvHPkyn7W6Vr7GhT7HivtuJldHJxH6KHZ1q0ygr56iYwCMhkYb/kmOXr1wxVS
jy8gpguAQlPfSgZhKlXqS3Q85FYkK6JRQmXFM2GobfB4c9ODQ4Ys20HEm1LAWbfy
ewfvXu4yTQYezMOOZsU07ojrje7cYdvmXeBejXV1rFaKmiEfRWifs64+gcLNfdgX
q2vVo7Rc1TFT+4y57P8CzFzcWq/Ny/nGHi/BOj/iEborlLG5fhIny1d//u0pUgQ8
Mj28kjiZO5hdbxZVbHp5pd/Sx8q/jBGy1bdyuTHy5oXOn+MPfJZHQ431SEFSf4IX
7f7SANqHJC6vYyCRBeXnxGgY/07luRg0I/MWO+JdAFEyWZ+jIZz0tCactq2k8IuA
9gVX/2HxGsVPU9ChCf6XHSkOkG7ob4F+YQB/GxBa8defKLlCQzFKy2HQ1ul36kqm
Tp1qx5uV+GilMfNo1KMDaC8WqYhPQw90E1gNFfOSUNYVVSlOFQ/kIDgSiBonnpAQ
V7gtNs8HXuPu4Jyan86kzCAEZr4udvJh+aKh7vIHrii/xiPLUHIljWxJCFOaZl6k
ptvJyIro9RHzcw/x13db4EJhZumDjMIZ9h/pARgyK0RvUT5uutbi0ANpKSuC+Cqy
XWmXCdqk4b8cXfCXoz4+gXCPazl+N8PkeJF8VOu7z+4GrCWZas57plUjRwBKXm3K
1hsnHWfi1dSRPzSCxdk2rJuxRpxwO+x3qo4LvY/LSQXa2zpRtXcYvSSzNlPBa037
UzEBv918oPDSHlU5a5hOk+A5UFGrZbtg0L1ZIxGeqsQKUH7yjtNm+i43M5tkf+n3
mmDEuCzp3b/PXCEeMBq1jsPw3117A897anJiKjqCTph65fTBYSmdihtnnWqvBfNw
jiO51GdKatDeLuRClQ7W5CxVOPjYNXD9zLy7rznrfoPIx1jqFBfDd7aIq6Hrh74q
E8uwTVOVbE4j6OZHT8/tqAnwHLLKSkvXPZiaEz3/4AZs/YUwUgKCQrfIUJZS7GoN
Va39nId1mxIqZdrZDztxwdqFQHitI3a06s/pGoNotMi5cN+7/24iQOQQhL+Wq5HI
cvMSCqR5X/omG4xMmU+vnELB0WfhtgAOpeY/2X8h8nsTkFVL1TicseyWqacqBU03
KIY2no0kv34tjtaZd/yLiVKe6OFsYyvIQtUmj5memmW7mfMIWYFzdO3T1qvsESNc
xKikNM0ip0wsRfQEHNE8OlpB9wEC7lsgg4/TtnL12cDAo7XOOYNLhkjKZ6v8fQxQ
ZK83AJNqtiDJn1zjkEw544mv1bYjaRYA0y0LsAsSPGA0jgMuOnN6zjsKwpDOAS4F
qntK8j6Tzp9qDkJPWXUUaHc1OPsgJ2PIlMYLwICpnpwWrcdx6OVfDcQjOePtQz24
h+s7eMDSpYA/bdr+LBOzhf/t3PipnoVkPZG+vOm33dBNa7CehfkBHEaMlNUbRBX3
BXHHo4kMjU0kG7RWtfRbgkViLIUCNJmqG2vafzt40ALceR6hZP/cQ4WVMrJBENLn
nptIlY0W1Q2VBh4C38p3HQW0Vbd30bf8AJmdj2Re2lKakp3dbhAfa4aWCgxSlU/Q
cMGpsm8ngOSia2ZuS9VAHt2GTTEOFyIDGlfWb3DnWAtWEYNn61ChT69aTPUl72kt
VwuzQ+2cRwk5NLs/5eqVgfDxTHFhLg3iaSeViBz/IwwdhjUsx2EWlyWTxK3w6YwQ
ImxjERNoFnMZGxaOjFzkdFPxV16uFUGin/xSmusZSvzxOjUk4H6VQ8RhIVOZG+qc
ZTBUkZ4oskaN8x9iVhCH2pd/f4q1s7M8ZMy51N8J7/ECbPjBjFMsDexCR8lgQg/3
nDIQdLeKO0WXwaHF11iJL7rtUruZe8pfc4lkVvJFVtHC/K1b+vkKzWzS/y+JUgDz
/9Em74HnNq6PL6GzdzOcZxwesQxgDsXUHhvXcZuIH7M6QuqVISBUc76TCAOIpPxS
xuaWjgHwHrOvUX97mwS/vn+t7oIFJHOFw1ObRdU5zPJq/SmOkhGwhhUteMWpLxQw
qsgQ3qAZ4DFzYEVMQ7f2yUlZj4KxEr6uu9tKKerSmL8pF+WG3MiRsgkpYGlT0jEX
VpQLdPjUnLYxY9a9jvJOs6RPNX8rzwLG3nHr1r2JtLQXVoE3cQhuuL28LUpdLPFY
ONTAiyPOc09FXeXDHn9UA4SnXP18V4WjCtz28izIHkNX32qAZGr7+u23bGfAOnHI
xfpPE9dU97r2PnQMhpYPrDC6otuBoDqzxnRpNZ+m0RarZdIrIYrF7RGpTknj0QEG
oXFp+SLGVeKoXMZddHu1l6oitkcNdB55j/n7YEHYkZ8hoNZ37nCicQZu3nokba+k
V2StFv/+IBPBmtXnR4Xc+HjuBRTKymOHXxa8uaRLaA6P1LYYC1elDQmdRqzq53tv
BjBPVajTl8H39RnPU9H827yIAjdqFPijDHE3ZB1eo4dYmVAPCVCnbM1AU1pPU+JS
wf/5NvmEI/et3TFj83UXdEk+WXSYT2joLrDYbrD59WA2Fyq8AsWDa1XXBypkggyl
ogmjDZYTXiq2AdLLp4mv7q+8IYi1vnm1k3iGakxQRxLDOaKHvGhtiv3MTmovICw7
5Sutw5X5HfSY1gQk2cLeximGJQ2EghZcY8QMdijyzmiDFVo3BCU3Ltpe7CaMAuJP
/5XONIsCPBj8tTtpQ0pKt3cTVIvQmfYYNb9UBiLT3NvsIueNofk/tJ/b4hUWqHht
snSbp2ySSveTIYFlKcRDK1kUqSF+d3eQReCNL/oazfn6M0Mgxw/5a8ISGeUu7BLs
KstYMb00WzgrLjiltzm5+0sRtA/K64IoWhnxiSrPi+DjvuDnMe64aSZ5Cm60MMy2
fglqQBDHupVvV6jzVL2Bs2zV/w2u62MkufX1mkwIIwBDyTvpnIt2dm04KIKeEHMZ
Wv7RG0BZ4LSORl+bTQh0RpuG3+YedehgnDykXNQQeu+VTz1H+EGxnG7z6kPhZVgB
FQTiqSPGpBN8AhgumPXTGNuzw1z1SypxtZxKy9i6s2dBW4kw5jrO9VWIuZ0x+jIT
EESLj+7aDdXtHkfqZCJKs2dt+7eF7331l+cfrWi7GS3MfYpCCbhgMtYTcqSyoYtz
HkeUu9SiP5clJdULsFm0zxCIGO/cLyMKsdAfvuqPUsVotrcUwV0n11DZZDp7dzzh
EcL7yuYvktsgYSubUweQcm1zSB+h6mJ1JC93wwA6eIw6WhDT5XgUzhvQjBXs9Ma3
2+Dy9unYQpU6cF6G5Y1PwYY1jHhn4Ud0NigDEElSGXlr9xwvSjH+c0g1OH7wo5En
bph1I8JgM6pZNGPZmZj4R8Q9d8sRbmT5lzB0g/J93PCyBwfvKJlB2hxdeAZF6yi7
3dc4IJHOyB2UqdRiTsyACQMqcd8bLRQS6gEairTGkefLRJrVs6CXdC6vT0nGwQzh
5s5jI3Srw0H53SHxJdrVf68gXI131vE9EHhdGgcoeJK/K50DULyGUV411pKfD+js
qdXRDC57i2N/du4Mmc2H3At8fUdCTjZFCFI5rjxLmO/PDxeiG588YE5150hlJULj
doQwPMrVzRXgsHHqNPwZfY3l088Ig+5EERnUXcEQ9uTqs3o7qgPKzcn37Bnu3xrl
kmerDWl1dhREYwDdqfw36X3x1xX/A2UzsWtBZzJ9TZ45e4E3dQd7sZTe+WgsUwdb
P0VLRn6rxE/RI21gFOKjQeQpu8WZn1Q4BRBuS0jwHekFjP8vWyi3gkxuu41p5JbS
8BuI3JcglY5rJaK04+E66I8ovuly5rqh/Z9GPpnXyJvx0ry2J+tfAPwhCWXmJXb1
bO/qwUu+KhqpwVqGZXGPIKMNES16/UnntxiN4TRHQSgCtpB15lpwdO/vzQbRHIeD
j2ZNlYQCGgUxD7Q+FnJC6Lh8OUicWZvwVxEcSqYX4iH39XhhwjWucroDpQ4HjPC7
dTx5jKTpJ3/BgtnjkFi9y/uJ1Y8r23gDYiTpdadVTriES3n8R+NrET95MMFDsOZm
2qL7VU5VB659i7uB1A7jxQxGgE7c5L9+t80MgMDtR2B6wk78aSuH2RgaUJvi5aS0
su0LMgeHB5i5uJ5+70VcK7XHqe59SLk8AQsOV8qW6uuxAn1DaEpte8WStKJM1tno
RW4PmGKOEHBObz3KvAB5REz72xSPRU50NA/6UqVf2SxjlRKw+iUJaRAaJSxb2nkh
YZHPpLIW5YHJVaxOlYVfuPFEcPDHMZwv8YAcUjwQQ7gq11sx85D5KKWPUo9MIv1b
Z12Crbg0vqpUpvqzmFCcyco6BDY2+cIOOF7/DGbWB0fdX9Mf5zl2n6fLSe5+DyLw
2yGX1kaKYf4/B2v2oQh309uS6Fs4gQUMWYl2syEYLzgLkUSunFOim3PdGTVjr+wt
ULiHjZOKeYJXnH7gEzvTMeRmlTlv6Yjfg8BM3wS6IhKR6FsknT9ie+WE1HPsYf3H
Iipy4Jypv+pY26q0s2gP++40vApY3RzRsA8mxFwVaV8Rf+ipGVabpKNMqsV7ejCP
KtVlvM+ISzWFDeTr5Ejz6WPL/GnzaC3EfRoP7zagJH6NJSEp8FGNiwlxqXFKY0ml
+7AaPRHz/aDJDVxzyPAf/0uXuusx5W7SFJuoo5nCDKcRHTFyqJgroZ6LImKWBbvm
nrybhKHqMi0XRSozevqC9x9NhQdPWZzwTvFpJMmt5oLSwLrQ1wptyr+bAaXZjHwM
8Z9U9+Yng2ibO0KjJoRtbhqTraYXWioLesrT/fjv2CQmsN4aM/QtGiUGIKAvbPz9
e3BCer6diMqf/V3v2fVRJIiJ6c5A62EnQ5kPVT8JDfbP4OcbByj5PaWgc0zyTcf5
9GF9IHFskcj+uaMpphqo/XMTxcixOoIDrkgTqa/rJeJw3k/3NR8sV3GKPFL0y+oM
Kc7no2cDgpkL1HXtkKYfLXm3v1IsA/H9Ar9SGYYdKeO2P/KfzaSsxmfd6rK4KPR0
THIUPrSGoS/3KKqUyyQYFMiza/USCB/HuZxCE13viXQIfCblBTfWPnTSsfCL8Sw1
zzJ4PU07v0ZOTHxfrXD/I22NeGkEeExQDhrWqCgkmel6JrBzHRoPmqZ3vI0IAXcr
oj8QfUsMB/SpHo2MWXRmPym30bmrwT+evKYPywyc8l3GCnFrkszRzdWZzG8M7t37
iaXvd8TasOgpN12cIvVOsl5Pyfa3FE9hPfd08l23Bpczykm08dKljvnr3erzuVdb
L96I42OV9XL7ZH/JX8d+L3W4eNroPZvnmEN1Rbkzs68NsPIP2aB8UlFxaU2F6B2d
xC1dt2bbeosV5yUh67fBSrmVOQIIgzHCaiybQUGXfPnAMZJEXcVJvQwSmvorlNka
K5OuLugjMm0GN9jA+PiIExHEb6svHFIGbc4DjcbdjFmQYwFhgL09nw87E7jDwyw4
e+sqO0seGE51YmFzmPFzCXU/Ti5474h8YKB8fNJTKkOWYQLHxAeauTW4aQvq6IaF
7zMDw+auBZqBYcH8i75B8eI/XisOnJw2RJQv/PV4GFctm9z5Z8Glf4YCXDVE/P+0
7VbptAkeOwN+vZOuzmn80IRJCmmnDl/NI+Vy2Oc3BCJ5DbFbmzss84yBLIEwHGoB
zgZ1LjcZcn9TC6k5Zs8BPFqusVLK97SN+4hZzz+VvDeVpWKv/nMa8hLDGpIaPEzP
rHfXiwk7awlRvyd6zv85roxQ89KT/kACKz0jOm3F4N2Q5ErRC3b/OCcs0FiRo8Yd
ae9e+lSczWI2U9qrd2gCqd+ZI2gsVw5eW90miKXFKBhsN/WnLeNnSI9W0KQKVChY
PmY9EoYs2aIVbDZ6QhfStXOVudeIeGH4xDv2riltRw7JbXE1IYZNDFpH6rwbL17/
uogoFM2oSmY23vkrH9hGJ1nIcKUvWDtkjyIhObTG4wpwgxxCuWrJMEnzB9VPWY6E
DcqLxEhTbgbJe9Seg8C2sq8pJcJfAcBTVTcH1Cu9GLAMuwHxRIo7N1fxsQsqUBl/
B+1f0ixctSisSQ++sTa2bXW4SWT4DCflf/OgI/w28gsZN8aTTATB67iKB8a/3yq6
sTcOk4+ujXjZlH4l7rRY7EcLwtrR4lbAwCAIVrIcRQ5cbYiKHG6ezqZ85rdbmBmy
aA5hlxVbLdbc3WrbMYkL9W5il0TfoQn789ou57x7cPqdp21XTDgoqbAEnVNgQoEr
L5vZKJzOfRlAnADx/blL+yZsB0Odn3Ltzl7JkpGOi5gVpKMxZxu6ZC5+veYb4snO
+iyR+ufnGIlxZrqKrsVAWdp46HKKuaxOLjNDqRxGnsopbuKuwSC51B7IMJPuea8m
xQX02v7GGZeZPjuiTgOsTMVwfsIj3abZgq6RSECvbOgUaIr8wM6jUZUeBjyopErx
rlF1VFMO2XFCsiYxSqRyts94DY93tubLcnvmHjnnJoRXKwHhxsSB+30lKI/wPxWs
z/Cxsz23drQQpDZnudxpry6nGScp3w3mmN5u3bIzelfuf14kX/LLEcFfnhxT0bWm
3BvJH/54dqFZTtlTZZhRli/nwo2zAKqk3RnLWR8aD4iY+m+owlKjTqthRjBvwM/X
DdjrCXfEW+Qw30G1W6p8OCKp3rsV0USgbfRBL3KJZVUBRSeQmCuJD7hmIEuRN51L
pqD4IrIEYtXmNcieOPZjqkoEVqw+mb4zKXLdSR6a2sv3EaClPGAhLsAF+De5/UCL
sN5N6ZHFCQrPmDXTvo66ju9TMoCaSWiiuL+jMCF/GqBdvEpZ49//bwUaN1w2MIeY
SJ4RITU8JCPdTW8np5VZ81YfNWopAT2Jy2vpVpjHhG5i82aA56nyaK7npaRbUqiI
1KrBCjQ5YE9GA/JU/1lsniytBZ/KdZqlo50oTTDoVEHzRWyfwpmQw2C6WNRxfhxB
/Ketk1e/u6/ntKuoRWF6XRvySoG8UY1mbV4NDbdMQlgd35pV97wsduMpFTl2k7Tf
ZGP2XLeGoOB39L8xZgV3mhXkkmXFjx2LxR8A87+zn9g/nP8gp10inHVbLvsMVol3
xYXQAeOcQVstykcpU1TxOZdEECopIi+GMrCjXhjqjImNmQGRiqjeK3ET07WadS01
K7FfnX3O3vk6umOZZisMtPlLyO52t07SMIM6fPmJ7M8u1ax/D21RYD5RhZBeLJLf
X2x+NWq1XovH4Ljj+XmkuYb+Rq5Nhe80YrDtcWmzeIc6H/UWOk6AuLEZuLGUgdgC
w0kqfmv3oYo+fjrIbgLMSbO72Z7YGYKCa6LbxWcxa1dnDToB6zabo24Y2G5jIEKW
BBH9AOQryOZbvunz/nZCazLcjw9HzV4JOC82wXGzHz3BEZJA9vGrkpnNdbtN5RAf
2NB5JveE2z/qHoSWnMnOkWuSKceCZKho+76hLr4EbKEE5uBAbGK7HAq+cDgZDgbU
/4eZUKxP4e29UdhTLH8dYWk7xsR+UIdGHyQW4qt73EsObSl7ZTqivTHkQdyZYZ9r
IPX2VMPcOjQnpwSbOHFus0CF93vW/KRUVST4xsMuzyM58EcbBZ8AXhN1zN9bY1ts
OT37U7Cd0LoV0i3V/6hC2v33kS+4ApksWepwxbXtsxN8gvTU+DPngjmBQ/YkgKo8
KNetNldK78Dmf3Lpj7E+V4QX/CUVNTwPStLlJHxCQ19kCLOAUeZs6cKNj81HxIdQ
VZl1owHIwvmJ6FuS8qy7aa9U0JFXL2VrKJ4ZC01eOJ7SosjfD6o4iAkuYH+Q/u5s
a/PgG/NiMjHqJ+8zTeLLYjNmXhkWQ5wlfikejGodEieIdOk1A8xr84hJq/t6mnry
2cryC6OOiiVr34V7DHnadmhMOFZlTH5hqoQSHiRjKcd3R1+pzVw+e/9teZIlyCBg
DFWHJjC+/xHI4Yp5zz4C1M2mZ/Eqa5OY3XQtRpSmwOP6IDjpCLNN5dTun6j8n2VV
IcxLNo7mnOJU0jJjmhjU6XdDXLuU9yd+1JAMOm5I7Iy2ysTyUVDZV8sgrmMklkuw
lchttYNISXZtXeUBYczPuTvx3XeQQo87iKai2H+cuXbCK8UpsXK3j1QaO/10nAC0
KdqaEI3L2jbFGBFPF48beqGC8ysDG1E6G4NoKzoTCA5ihU70VgtpQB0x5aus6AYz
PiqJZSthh6a6fNkhH3YZ5NfD14nZE549khO7E5gcP7+g+EDSAvncfuf4gkeMq96Z
ZF3P2HKrOkiB6SZnmEkuu5UA3ECH47XuJGUgZ+GMr5TFeDL4KkmeZFs0bgmdd+Wq
EOr30Z+D+9kaRBoAi02VZ9+wDO2eWc863oOWlEXtb5UjsTT1skDCDlHNMHl+FT+E
5XDhL/+39PcYhEegAaXLX0e/Cu47HU2sJzCEPzteQvWDz1D+J1AXMs+7vDoiCb1D
4a5aS07o3wDz7+LAZKyxE5H73wdfuPLmBOkN7DrMwKGA4uHcaFBkYat9qTcx3lt+
tERXWam4mKcN0P0kQY3M6u8oSqDoTltBLHCILo3it/Zol2E3d3gvzXdwCN9yt/mQ
L/u8PfQJZXM+RF7wQYb508Xrwxem/sVO1pZp012t82LSAEzYRi379ep17ct0DBI8
1yiTA7JJxtC1XZ0edR5hEzjqYRgd+/sdIZ3GforIy7SsFLDXKZnL1ebCDvwWNHgd
AJGVUUoGXRG+YscpdrWtK/1dYJR5Qg6ccy5z/GsHvQ8qJu9ktwlEkZmYPFOnAuVZ
Cn+yQdYce1fa7zyvhU1wCEhbevmGe0hg5Z6TGTzqQpGCcEPMMfQQXk4Z7W22sWmz
NyZgS08Wq+VD+6XjVEllqWYyY5jJKn1NWzvr0DKdgMyH1zpLu8T5UM1PFn1OpvDx
/RqkPwuZGk3zVmV+ryMZCDL5NpJX3eT/pAXtqhrHrEvN+HmjsW0mntOOc2e3irlX
PmLPP5bxikA04Gl6edHtk54PjW+0lpSQnWDvhbInIvcGUERdofpz8nyW/7KyE6Rd
p+jHYVt1UqQYdCYZ+gPUHo6eViaH5c/MGMHZEuF5geAUa6tJ/Jmpq9mbzaITKQQU
QqPgnYCivVpUqAsdNGPZCownseWUz3XTMXgSQ35eoE8s+MSv8wDKSPoIyoo1ydB7
VE+pUjQSC7njusMCQnGuAdcr0s0wyqu7d8hBzVtxCyV1a9LVczme4j4FKO0osiKK
gslXpcthmoNWh2tOlndSFHRgs4iPedtALa2L43bZ1/krTaQkeU+HFSWk2ZijtbVr
qvSpVGVnNB9WNNkXqsnq066eRTHuF70YQonBeY4GEf0Mgvw7uE2ctqTxgFQA/CIa
EXkXfEsBM2glkiyPsMggJ+YuU12AgmuSDndgMFw4Kla+IvW9IynZtzZqtFt22ZqC
t2rGKwoTyV7ko/BhpshI4K7My/sJxSkYsd1ICf2XXOgki7mMLbxrrkpgPkTQ2Qs9
pC1FDuz/ObLoH6jKH0Xv6xayDcEw3icT+T3Eur2aCad8qY6MaRGBSEUbpSARBwq0
PklERnYKDFZaYV1BAZfCHiLDTax1EXVRAJ37edcvF/hWgvp+TfJaUnAhr8lsUQou
BhoUED2dknXqj6EVMGnBatRPezO5ptahxjCtEnqme5FvqDixxklebTPKywsNhKO5
kCHPTbKjPMoTmqrhAsSLmdCjOF0e4yoiv0ISAn8xwc/R0QlJlU5X0oPyhkiXstLk
X9zHwrVGnTl7StZEdSzS18DZ8xktm4JxIlN+CUtjIYW+Gg0UBPSAn7tZBq1tvPKV
8Q0l5ZF51HvLnCW1RFrij7GvwLSrtqHZRYgkekfLA8z4coYneSmNWPP3kJc72KUo
LguNweV1qDOhLk3gxlRPz1ZyrPhw6hCTSPsREzMU+e6yXi//5xfwFNxs8lVzEQxB
2rJ8dRte5k1Ytbe2FkhGsaCPEM+hW1/tLlj9AgAZqhj9NfL6baqXNssP/2sc44OV
I+mFkhvfBWZKTwY/t/KGZqexvpQ6bzvnOVubDZqSNg7o3fxLbSxonaMbIR36EkPH
Q3OhV2Pe4rsnq/e0Bc7lLMKftU+dfVo5eEOus10aI1Fmedzf1D1LPAG/nKQSS9ye
WxvK5MtFGeuDRMSfQcDROqHN465jJ+qrLbVSnMm7Zy/5ZUfIUzzBgk9Bp8oeI/NC
7sBNcu2JgO2Fqb7SgEyg+mboboAG/Db+r3eQgs17PswrJEwYfF6n5L4pFm3e96pG
A1cdlgl0v8TEYiByC0/PLOnAHQV5fYvrHGFslupIh+xW3YRME5llUHufeHXGAo2T
HfvlM/posz5f4dnlt3vwsbtlauiNojKCabst0G0SE46w9HH4CdwOItt/mJxaON3S
/LWkfWcJ5NNwqYwVhOviFJlN1rePy2eE9m8+NeBuTj0i+OtFxdA94ESxfgiGkCry
sLpX7JBmwe21euAzM0Xkd1f5WIUiYUz3yRDS57XBjyoTId9b0QdtvDA8dkzrRWK1
GBJdjpBpiqyFjvZ9pqdwLHdBPRnopMFIpxphlORTdDNfrG2clhI0yknXFkfXwje+
j1BNapcEKQbnLM7wWhzZ+Fxq/4G+HGD8gPPburGgQiBhncBc2L4+AW2QXBC1ulPg
vitC0KtgOJoSLdGSxnsuKUU7MfFm6QBj0N5sV/1/t65rEqEit3ivFBy6ltFbVdBn
cEWF0P3p4u7ZZvHJZ/qehOnVzyK0z0SEr16nut35a/aBr1TnlUofMS6ZiLdM6Rry
15IVqtkZDbP+5hA9Tdl+rLzdzCKBOE2vxfnOH/otW5k+a4B7JkiUrGpDVexpBusB
4x6XdMbc7FN5n6vtcKTYthhcRcsXi4qMmPAK1gLY+cG2PLOFvIwYa29XzuaROYdX
Yucmu1xV+CWgVEPe8Izc8Ag71ZYaDoCByqfj3kndOX7B3O5mNwEafLgfqSTXwR5A
8hewrBVJ8go2pklEgC91w4bDqgwLgYkfjXbJD/rafrUq5zcziqRQ3Ync3qhWvm3o
9fKnuwGS27yO3BKA+7HkbMbRoZERzl758b1IczmH7wLWeyVItN/pCu8KSp+o2LTk
Wy5t19Rn+aXYTGGqvlBaiLOSBvglBlVJS9e5HHFlBBwd5Vo2FCrlBTUreMm9omwC
ETODW/RhnMJCCv6A4sqFlEuEe2Azob1oHPzETNwh+1GeU+uWuhNhKkQdh1RtZLmN
tBrK6lpI0YnnolBwQMKgGzZ1P2E2dhyRqepFOmxxyv8ksAB7f29H7wUWMHlshaNu
DVJElC1cmPFDbGxocHPsT96/ZEuuszolnPIig8+TmdTXPQ8c2zivgnegSizunwuv
52t6AwCa2+seTlYIp+i8GbQRros3UGZAt5rcXOp/p6+89f2tQlaSnazTkNdW9n00
oop5pQ6YinmK2WWrHbz11y8LwhJ4X7pnI7hSAQWdTg/Ie1cDTMpq2+KbIsZuIfNk
2dHmDV1+RpiehifTSfA9f/XE0MUDI10NXVEAlzXXmepReYZVoOcr153HkIz2Om4t
jQk0+TEE9aTRprcK8POSAtnRDMBxKpMnwlDpfhL1DWzyXGD6Wc3Z2cERHYqQjpK0
L77hPwwEO1NoliqYjTkNict/aJ3+vkVTjf8oIBy+zkJQGCXJI6QrQ6PGu6lDXC2F
0DQhtpYxkkAdv6xJuEeqxadOqdZuaShz9x0i5/jt77O6POvX2nDEeDdwDcIP7MoI
/nhJNd9xVT+9uOgZh0Ya2mMRCWm1d3rUvERiQpm/CSP20jz8lEqQGvXvuFrOyzb6
x8MN4dbWP2Z6TkDZnb6NHW/0IxyVjMtIrV5/K6Rv/3XM+2y9z+UFbPbIb3za5Eu3
fy9txQ7Oy4un9Xs9sP7rP7JSfg/xSL7H7p1DQnFKYojjXZ7VRUWUND9vGfERG5Ka
7lWSWhdGMxX5LAI9iUBk1Jg4kcxl7pePFFQj9H5ocXWd5yEd9Tp+Yj0fVMjanvWt
SB2mqYWr7y9CkhGht/cVYzKYNzcB6sVYkNb2r77s24uLSRf29avbTaneEqCTQd8i
MtYSpy+HgPUBGx6eRfE5TvSdvgTKNPknvE1tBMBKrj4x/P+/oz50IUUsLTGAxLJi
4/VjZQNoQePqJsbd+lgh1N/uPHKqisbWXAf25Wb1hFg08mRIy+i/dCN3tr1US0oy
cm43oqqC2EM4oL6IrpVljW4WN5Gq1UwTKBaiq/GTnH9+luKfw2e2E/jkTw3w4OAQ
GfTi2nZtaW8zfC2o6vfu6DxkUljylmpzQU5P7jh2KNQ1ThUq00TGxIwL14L4jcAs
+HdHv/4Yb4XCLVECJhIqGnus1jj6PiQMutk5H7AZh7ysDE/U2HlWJoQL0jHEQGbT
VYhFXfH2IPtoc/d15vhzubYr4v5grSh2bLk8s1iigUj3ALK91EFarCKJt4ajm7IF
eK/uWBq3xskJtLgg9uWSFqdySvKBAF0H9/VeCjYOglpAlONvp+tO1uwh2P/YxTO8
uZ3S2Trm37jXu8TLn/cUqhGjfwfFFU4eT49fX/4XYczcic9Flegr0/haB3EMZ1cV
tBmseg3empD4OqLEA/g6YrHMYpJ7qyi64ejzaYjaKHv13ig1iA2Ed7wrNAe7wVea
ClMZlUYvalZ4trORgYmCDUN46dXREAYvbY01xIW62oMpxPi9hdxPIAVPKIC8okRW
8xT/2EIKGy4/NSWaB4WKMutEnjrLd0HKC9z+Ajg1pRgVYeVV/Q+06SInN1XtS6Np
Qb/jL2jA9S7+H26j8+Yj+9IKF37H3J7xoE/nKv1DMEiApqf4noM8CzMtTQ3qZvND
ilIa+qmJQz9mW24LMYL/2L0zD6PtVLg0gouexzT7Xefjylvxzd6acGD3Xubel9VF
pE+F5VxXm1UQa5ikmk+g8+eldVyBY91t2y3AiSS2j6Se9nB/tml9KsXEcQV2cSyy
qXQukSAUICX+5O3l9qZHBzxG0i9K35UP5vAlsCvTEgGy7GDOpcJMP+sZkS8KQhJb
apQ8k5NK918pb+oizcl6gcN7G0DZEPY8aNhuwpDG7/DlOIVdbfji8zeXCajyU4N4
iTbwhgbDgDakDbiL9kfySQ1Y4auG7qNrwcka4cK60ZnS8aVjp01BHiRrvYafhRd+
yA+HdPKF/ygOk4F69c33ML+zpQlxW98SI39Y9u47PGXKcUHZ8df0LmeuZL0UenZS
T5IYJNi85QwhzOraUYJbDq09oDjEffLTqmCNZ/XWhuIDAXAsjzU7dk+Gxw39BS9E
0j7ClV7UfeK2l73dohqu3qRUdCYN4ajsuZosyfpHUoq/TEyp4GJgL4tZiSfLAxHr
nXv5SmgTUANF5ozm2apOF6ZE5hg4l+d+HFfYCcq3tTMszPJ1b/8+2MET2fhVvw5K
iCjiZElxHxbyN14cZFcSEE3adHN08iaJ0Vu3bCOSAoOqNOkQE6mEtp+u76j9L2a7
lbBBShlVrOHBl2MTFDPsn6HSHaOqAbukqzXWt7mYPytux4JuoMsC76MRIdAKnXwY
VahCb2KXpCo3bHwgg2kxaYRy8U6Q9UEvJY+UghGkBoK84qIoxCabpYitG/mCwjbR
f5Lp0a5wGRcd3os5tjUVGitXI09JJcXHkxfpjArx1ZoWYGBsFA2TvLrQIn1t+VF7
HBpL5GBW6LNchBhzmu6jeBHnWEu6s84JZ/zMz9hM6vszqEsfKb0KpQy3qY00M+CV
BvRtVuQyzwA09bFUqVby7iBOwmv0vdruU8Bq9ZgPktnx6SI7z6n+3X2tRYAAwDdI
ARrcwRBWb7nyZIJIelXeCZ8C041qELV9uDJmoaO0kFpgweRIssFw5yXMmpMw9ukX
yWE+zr43bkZSbgFf3VtaTCk5yVEqEcc9e8TGzsMWW9LLQ/TqlCFoT1T8VnMkT2ZH
3fLZxGiThvnS6cqzBCH+S0nCvJ+q2sRai7SrPfimekXq4UjNWfowdMEAx082+6Dx
K37qcD1JA3in2LDRRRC86mDyupQ3CMQ07AcJm4pyFjP7XhtSdMIPLjzUOajWMinl
Tecq9h+7Ui0FLsE2kzAhoj6cuyHajzsqjK6FZkCbj1rOUdaBhFnKzVWq6DcR8Cyt
AdNy3OPLwLAfnQD+J9UsPaS5i1AzJFshY+wc1alSIh81qbCLopbjdWegRU9DW9ux
+hlaozVFabErH0MEjLSFd6ULxbW63zVi7D0TrAaPi7gp7jlxdr+fLHWdVJN9wT1c
jr1QH7I4TVyv3NkRAY3tzTjSAnWo6vB9Nh+7mIPj28boRnq7+LQBagu/GkoCVmeN
VUMi/8uP6ftI4PEnpcps7W+sRaMfuwhXC+jxK3MEDtTUNNS+zkuFNB76Z1VSuzgi
wuW5WFZqcnlWZzDCgUdG7rxEFNW61ogDA1UoDuN0DACfdIHERU41awSEmGD/Oaaw
OqJ4svEL7bX/irzMQNsGrpxWMQj/sULw00nBjWGDghFpxIz7/BWooYTKFTPFJINu
90GnMJ2mj9h1TfF4/mEFreiwknIFkOOjOLMJAY1+ElXu78bhsMq5UeluhasGekDn
wG93QSFSJTp30U3JZTW4L/DbDykX9BJwI0YV/eQXwV5KcBzRIczvglUFDWerhDKZ
lv+X0TOw3Bm3fyoq9o8p+JThfasgd+C94soWGbssT0CLa+QzvlAubYY0gpc9KhEu
ebEwvz8K37P3KkTqnZJ3ezBakEtZNb6d6a8SlX8wfkD095OXfiZMwaRSZYCiQcIo
5CAzJJZBnIZJLA5hDNFeK0NdrxWczyKbdwG28SAVOjs6gEB+UpzMJd/ZFxcqVP2A
KHTYNZwI+67RLJyZZZ3efk4n7O/n3MD27rKs1UD9k3L3Z0+Ipj1SqdjqU8gLEmOx
QJ7WMIeCGoRfI+lGnn1aFwvwFLiw0F+QLnnYLepTAlQGfn8ahFOjHaZXqmYNH2Po
1p2umXgbwHTgr8KzH/J4v/0fE0l8Zl9ROJiM3jNeHXuAC69Py+UvrjsjxQnmS4eg
rNtfoHGpkxY8iNMp67wcSg4c69nAincz3mRVNSBSYDBmBZrIpqfNPW7FWHlyX/cw
fLD9i87VudFpDBbJlcZ8uta9BxATI4JW8ZYzr+vfCnAjLwWYqIpSbQl8li/tU3qv
sgi5DjS3t3dq4b6Iyu38ZsShw9dv6uX3lIG6tyTeSpVdywBfuXYJg8O0KhPV6pja
BcPvCnnXeSzBqZAOdtSYqTHpj/a7GzUtGWFeHBdX3HTv4E27mCOQwg3b89yAb8i3
d1QfMLs51OzLoQfBtXDQbdRN3eZcuO4szraoefeIR2owPHHQZ/447uSBStxxkCv5
uxukH40A0qh1B21FM5aTSzQ/QOPtWZMsqvum1YCzyO/SlAcqpZ6qdHY7A8HQcReK
9iUQVIGZNg+jyqbERwuO/2Aa0QxCTWehVTEfSeOwn8cc9SP8vA5HHaj6aBzPCwk0
9wtPc1/2Wwb0t0gR1CuTzfJ1S+Qag3Si/Th4Xlc85mc2uLW6CjafzrBvvwcEZckT
IT+qIncovoNrQZo6/XjygmtU3L8p4sE+scr/fgjvqq8dQ9f/rs99JoDHSizwOCU0
PGzMd18g1EUhj1BomxCMk65WzS8RIa6ITx34n6+da6/ubxnD46u4NtILKP1vDv4g
ZZy1V10Nl49KjzPDClrjaeaOqxesUzEGIhw/ccdjSJWnGQVUDUNZVmeHdsnqo8tU
n0jmoupZgP5RXovRs9WAXGlG2HJnUczgcUG9HxACpF5dIruDRTzfRx+Zn0gDmKxG
IMWRte6IoQM1ypt9dP2y+zh7p/o722+ULxA8e+Wu7Q+rUz6E5OZmcrLjzCy/Hf0z
rVevKRQwv03PedvE78q4EOxAV0f5ObaWgwLL1ClcRofkobk7JhopcQjn4Mei+2bG
Mgj1PyFZa1eLrb8OVLE0c/aSBNC0HR+xAlspG8JoMf21dE4W8jNtOxBGeEaP2W5C
z8LofRnpPHNQZzQmXhbrhzOVvJme/Lhkro1qWPsWC5Ja9tI1AkT6xnyeG/97DvRK
Ap7W2R9uKxKZOp0RPERAdD0cnsfj/eG8+2luUeeyJeBRAGExdFqhwd81ojAvZMiz
CXosdaqMC0KU/x4G7NVF+yBMBAjVTLHqH3iMmltBtNMTCuG2cg5pTYr+WUqFXHNH
Pk3vbDzb22Kq/KeioKN9T2SvykhuaFQQZUd2oRUDvqHkVtjcFsxhYhYzp8reku/b
flKjRn2qDEuzArX61Rt+6Z3pO803GTjy11A6c9RHzjcUJuroIlWaNJwqVbNfrHWi
/rKoT13QUfhqnI3C1rv3TstSJLzKFtcSgpirOc5Ps8PhpCmzlWByPcj0A/oyVomb
+nlpgTBGBpHngywuN+o6hgrYoXAKFQJ9hgCYnqd2NZw1dg8PoExhinILEkhU65n8
8PGJtM2spEnu9Ty/qX+CcMq4qDIlOLoBg1SjsO2NbxrC7AdNl9gHwM23lCeRmD68
8kNou//YdFEZZH8g/OdDN2rykO+I10AgIBCguYJEGso6pMoH50vY6LbYEfoFeKot
ZLyWIWRltpl7Xh7wtlUkzQOHcbgZPkO1kInlU7dp+zxHtJWNJq90B89qWG6R6K9c
8gD2oATcRo15RobSST7osj6CBk//FXRsd1eyFGqcgYc4EYRMfZjuKvFlSQPoSo8u
2DtbHmstidhHYA3uscNbZ/QWwlT9oj3LsPqEpDYWVywFD7O55mOKWZVPFsK0mK7I
r2CDP1JyeuK3lm6/OQvtrmnV4Vgj6d9Uocus3yiC8kuh2zo3fqv73omaCPGcrzL7
aNbjLuYH6gcxQuO01qhLv6pAThcTonOb/i2+ZIR+GJbSs9WnTOEztSWlBFRdyEg9
tNLhPnSARlQRCzD3aUg1tJBx2fotXO+ccmfBPmeUZscH0no28GFSdBGkyCyXvZuR
A9VPcKLChsp4Njxaxw8agbTMcPEi5KngYNsvC4kRPqvPBIwL23lKc3ZDxvs8vslu
SMUXoOI+5pPWHfnxWF8PCPvi/d8PWO7nMzSqmC8HXmss0m8wVc8kzC8nqv+76qa6
uoOF7y9qEp127Yw3etZXUo1PmUCkMKGMEy6SH81SheScRBsL+xwqZjixuM5XE8wx
+AfoV6GSmvZwZT9gc+8S9M5Kgyf6FEJV8J3jtubJP/qJ011LPtlXCCovBFmuux7Z
Goi5GOtLyhb6f7lrhklpIfkJrjp7woCemeL2L9eOcl6xqRgqAkpvGtoqZrJlGepw
miArtSHad9xuQWI2dEXB8rCYKE1SAADu+rNeXUsduagQ1hW1/quYaLQ64um4/Ax3
/zgcnbBiZ07UCQARa6v2n6z7LuaWZYBJfEidnjeywas81ir3FtcryzGuUUwQ3jc5
mlq2GIUlOsqhCOWqZdaSqknWDdL5dyUJLvAY0bl/Ni72dsKQtZ5dVryTPV+g8vn9
Hi+QJMv6WueVZ+Wb8qbc5UMTVJu04OLygNSXuCZnss5NkSe6yqY2cWy+13Jof+/s
A1XNuUK9WCOzKzrBMG/MLS5DmHjacB7yJq7i0v8O6YxZRxCiJx3e7hJnxnRq+M2l
QLjL9LCw0RNdx1vu9cj+o3yINDj1tTF0EJ4F5v7NCSihtWNY85q7EHvbYcY+p2Ws
dki4QHYRGzYp9sVB178j35K4oUy1FkCRRCKl1e9vRKZDM8ifnzSXgA13+TabmsoH
VCvp90Ehpnv8MwJiWr21KYr/YkMrxrTUX9IQGxRB3+/AEtnKvTfBLl2SnQlwNj3r
rNdEt8yZEg8xuAQaHbgHUVz0KiMJnCpHz+/knHHoOr2Z+13e7fn0iHJj7t/NNwJF
pmw0cFcgXfIA+Z4wN0qPz4nwR77ItwmfljYruzWpyew+tO832fcXdmghyHXor/b+
QeG579SARxgIMCzlkSpSKHuTsP9PfWvVJc/xn6THtk7cfT14O5PF/I5VLd38dFUd
8wGW7MGiUW/9HPhViaoCePwabhzO4PrQnsdpI3yHMF6o2M/fr9JZ+nvZlFYKLDDY
qopNNABmMB2d3UqLtxxFQHcuBUwFx1WzXfLHoQyXYFKikHfj1pwZ5X4pEkubAniC
kEPGw6hNtRTf4B8Kc033+2NijwqcbTJPbpq3YO6mcQ/jkF/H7jGBTU/YOsA+rk67
6GC/uc/TFxaxrC3o/34QG0x458XedTjRSlxcfTS9bazvwBJSIdYXvPMFOX2qaV7c
fxvDv7Qh8o9HrDx5+BBH8BU5aztUwm6nUXf6CbBMgvMaUj8feiIy+Zt49lZzht8T
aSo45pbiYR6JX26qEuJF5nZ83ZGofFfXeRtYsOcHiwkuThGRep9/Sqip7Oxp80MY
VqxLzq92josxsWgf/3rLsIJngffuUD0JFpvnnWCs6BwexMcrRKMe9MZNw5lIAi/2
vb8k4anxhUeQ+EbR44sJNa1b3jNAwEYwgGTAtMRvx2fBxerG3JJ6ncOPVftVUWFZ
YSaJnR+Fm4DXBzvvXyTzDGYaIfe7xiVbiU0I2OseQnGMNkqQRTJTHPDC9xBsOqz+
8Hk0yCyGH3WguouzmjcQUcclCB/j1k4asM70zpiCHeAhg2MPDTsR73rTleMojPSW
KXNBXOOLSwoW8x/8KJkzQD9Vi/e02Cfas8Ct2HAkSjEu1tGpdKGYSkgpaoE5o2VC
5fvrCKiOd33HuYgBaLxkm2/05g3pf06YeR+QM2zj228IOKUXaJXPfFjJ2PH0iWVm
56bt1YkfSjYGPeItTfi+iyLZlY1btSG2ycbn2eoucKZ+IhQnN9oZAJmikGBCUelo
DytdKfrhS5GgFYdpOGMIUJeQvKgysQOc9YKBkP8DK5KNE652PNVxWleDYawByEXd
P8Ta5h3YNXUD8FmEAirNoeBnKM7TD7cPgKu6PIQ2p+TrLcaoZpnCAH/VjEjPwvZU
2BmRN4DZeIPVqswi+eOTEbSmZ3OoZDtaVSsGtk9gRuQZL07r2zdGDPZZZTOc+ccY
TBE1i+Em2VWP2zLKlpuizaR2t96R7L6cPbBqSQrmUvm/XybZwpbCUa4QQaP7De6U
q6+Q4L+SymQmpTcG4tRIy/a1GoBAYjrzM5HTdx+OJK2q46WvCC3iKp0hAzKpPOlB
pb4ZZzGXx5WzswnIGSMgubxErDbYFaXPqndp4BE4qv4jy2dax0XszPwNE2cMuWUi
NkHrJNvS+VyVbs5ziAge+S45Q1BVGu9H+Td05ntfmGiIocyK3GWKUrctvyEmOm72
LUEoRIs9nDO+nVbrL6NUKufenEG5ZAsGQ9BaDj0ypU/0LnsUC/4Ho5+cM0XoM2IW
xKHHGpbVaF70FdBDORvypVePpNjTCdta+Inf5qTa7dgyc2Wfc8cs3DNa/DyDhPvC
Nbi4q9TL4RDAhExVvNvtW0zK/dSS8tzkY1N8vYD9paNJ0hXqYq8lheBonr/UGDq9
IrO9Ik9d3+ItV8cIKijmG73H8kAmhzRqi0pMCTqWYQ2v1hIl63z1xH431V2Sl9LS
exhBDR8P5A9NtBB3Yh+4CwKs4wQU86aUDH0Ga3tgxDp+wgnJ+Fe3edn9Fopn8X9S
Uc3ZDzfXU2ySWisaOFcScpBLOnFSynjDMyBYsPN2dC5p9MktwZM3MyAQkLZ37EMG
EsR4MmBw5W8CGcvk0LIaE39UHItiaEkIXD9/NWjZSBQyEwc3NApy+6xgYYxEh/Ww
G52tTWKiZnZSbnd5+WZDAGXqL0AQtJdB/5I+HAt0+t78Hvmrj6RcHJO0FNw5IL85
BcoyuuGK6X3iQ0BPfWHyg2qHBmTw4J3SNPcfA0iWEHutx7Y506j9LivtiHH+r18v
8tkQ2lZcc3OvfD/Ewzz62N5a1CZi0QrN2UGvZ0HxRlDnQgswduT6VKqcOA0W4eGB
SJlSEiOXfpigB1BSZLZS7NUTX4ov0dINa33OgpQyeM7vfu6egETznDl1sjt3uNR7
e8dNODCpHXvxVm7zroQ5POWEbJZhj2jcmn1SK6LfRsxpyo9eoDiz9JFbS5GbmhuE
p4KhxXHUQe3Wku85+xriW9+vOuY0lbS2ihVTd8XuFLi9xTodtGU795j/PJWqMbOW
Z0NV+79NVmx2dxRrAC4cTBZi5apyrLUwGNZQxY0yOCpcaXgBb5oYEsODrMGnsP/a
lDTvQwqe0a1Pgx7tESG4od0KSBf2TF0GHlOXxaZweEyEIoHqA7ijBNX2OdCIRksW
t50VR8HLDdszc/hRM+bjyDIXfCb+zQCSqkXqQm2D5r+4JJXYDQyEHx3+sr7qdtXa
3jI+HXeW5MQ9TNlxsFuhW0ZyU5HzKle12W0wn3/qXL57ecaDgLDXyoXwNrve1Aqk
Y6Uef9uefr4a3kbZ3rdXx5ZciuDZztbENW1rqyVpVL1QfVOKAJznxI0lg//YTCDM
XUHVdgcc8T2gpjo6j/X3E9OdiVOgQSHT42mbplpD8rqCApGhM8fvp5GftZxHF4Qz
oedkDmTokn7Shnv3eiGAtJEFUglds+7qOHQ8PVdNXvcYCZFJyMwXv0nIAZybVk9q
Q++3tHocQBAMX9YBGpmcsC3+A3NcCxghJaQGKRaFmoV6YazYn03GiZNGqa2FLBte
IQ9XtkQNCtSNQPQ/BylXifwP/CHNITwxF2E3flMLUXprUBJ4QZDN5UzG28tE+jaE
1CAddGzXEcwLit6GuD50cpGoR5RGUZ5PIcTPu7fxQuFDe+6jFU2xF6H6Nh0nJI5K
6xLTwhjZxx7RWOxWgQWlnsoh3RIIpbPy/VpsvINR7dJr2eWiVBNNScyf1C9fPLOA
93SDTowGZjc8xWu0cCVcAQY9Q6atqSg6EHlZLpNBqFQeWpIS0I+MoMa5famol2SF
OKkotA+V1KgyTPfzqWhLAN/6FxQQ93HJSQGWp+hopqH47wdP0LxIFR+C6NQ13Ll0
qYpSEvsoyDIMzQIFWRQCZzYWaGmcQpY7KhQSkFa98RN0NbJszmRjtUUQyD3I+afG
Gyqy4O6U2La/LAtvCjyZNuRA7y6L468rRm4kA3vX+i1yEx8HupbE/BAzK8xBUJ5c
l3ZESS/A1l+06r84genqyGgiDAEyutKyJV7CSx/+IOU1sSWftazvNB8ESv0u3N16
MrMp6XdxRP/B8JmBv5y1Vqpp3cmfTFBXEpIhtpLqd34qKZ7ModvM/wRDnO7eZ93t
kHGt//r+QO0hrjJD8YsL08sHrm5gRDHqVWV4u1bLgm+8QYrI9iPjbqTFeUFIcFNM
tIhcQdD+Hckt+WbzBkM8tQi1O1gKO77l9msY5Hu/GYDLMBp+efqsae4IoDESMVqx
JV8LZvmWGBfh3c/pE/1NRl5zyPhRAO+xsTpv1iQkHaY0W7SJRM8vGiPLIt8n5Bup
dz9OM5OJ2PzIQHE9gGVNYo+xNjdzDfxGJdaII5GUx0r799YyjWXfiTGWtUge26fs
KHpeNgdvmrffcJ8opzZscbi7AfNGbL1p82iL5FvfdMwp0t8znKct/4i1K8yAX37Z
Dge2Sep5+YG45rOJJdowun01E6Y9QyEpoL7qohtmLbGckiQbOexB45Ifogy8Zw60
l+JYCv8SiPbd9FfjYETeT/FbnOWBdJswPYqT2wdWdTux2XEfVAJ5vKKJnM5ARfQj
XimoNPeywYDun2xRkKLoRCA0SVVNZgY9b3iqVeaqUtR7zW1MAZTopI28m0X571Vd
lLJyk0NBglZ4bHk012eEuR9TIAz8x6X2uIkKKsR23sDV7Zx10kiJrrYkrMssjFWy
0C0vTZ7TM327k8Ngtow5mCtmWh+lcX0g/JYVtn1dzj9XFxguN52MHGHeW87SG38M
59m/ykyerK/UzNDLktRyTWYrKqz9m6sscsztswMhwoAScRlQ+Iw0qnHTX9P4GztS
o1ID2Rcs9c1QJEGA2H0Y30aF8j745yfNlYFp1/tT07hhb1JI8bbKb50bpmrzVkG8
d2YzbaC3vgKeG30yVCMWaWa+dqvzdOhfO43SWKEcvPQhUDOTfEcYdVJTRJ1RGvV/
avTO/+P79oBo+RfsRS8dNH+yCwJ61jaZiMW0wdUW44035NKa2y0OQK7tPkKeqxSx
mvS+z4IlIzA52yL4hVXfD7kS7PMxf4I3gGXJKC0WRCNWI+Q0nd+0fAVg9Cu+8ueh
cC8WJaPc0lp2WQu9T6HrsJASyPGkoNLZndwZ54fgbBReQiNMQQvTKgZ5hsfSCnzb
p2qD/k2w5QhqXnRMVxCReAVBiEeFPPd6C7naMVH13Mh1D9ga6mTB5wQ3XBmMoaRW
ywQmup+zHiCuxIewYzdCxTA7nx0IwhcbqU9562do9Bq63vSO+RQC71QUAxEjiYQZ
MxZXFefUniDkcHFXHO0XNLY0DzNCV2kPAhIsAcXLq3vrIcDT0VTEaRKnLq04ivod
YsK+qytWXcTDiDD1FJ9NqTLo7csSWOQ5573niBt1PlXppdUEelUZ1q8p+lG76Tys
EH0a5pr9DZRf6yfuCcm3FisZCgnq6vo2qrY6A/RXCf4ecaYHSx6KixubNkI8rpay
/rKJPzR76I4Km7ojnC/KzPfNfq56w9QFLO3UeQ5RV4U51/YDlGQlOf7pQSlySZXQ
73ytC6pc9JAMlgEJ4mMThd5g8jcFUMXAlhRlckE74lNNaLtp2V2lORguwuFxBLPQ
8GF3wIB61AH6nO4wVEsdjXciDBFpHoWZnrKB6PTAprCqEme0+3QVL7kccMZCuInr
tOtGVcrGsh9y6vpOnAjbgk4XRmzpuANmCCQdvVIg3UnMmNLNe7BiUjPc5eUSDsMU
Lv4PfauydVu6cVoGdAsX7s/WLSvt9gCTtKUwR7ep+b0rR1kMGpiiejp+rgW6oz5N
YG1HlaG0IIDeadkk3fn3zfxmGyaozdimmpdGw5MbHeN1IrDiki2gGVTTFFHNpwaB
xDwZpGyFIB9NZkFT1ehtR+6DLvv2u4RH5e2gId5hhhrdU6vOhaBzw8vfOvcAueZS
j5MYoyY+vzPQgdZWfY8ybCXPiDn7oV/vKa5lYUfAShSvYQLiGlOyeAnCOdJc7a3X
41oMFBjJsT8R2OOTqpsKdgBTKnIvzIIqFm7EL1L9/5eg7x28ph1ooZpf0wHauP69
gfRu2IpnSoR3aDhRpH1+bu88zZHeXlBAvfvb9DQYjqMB9/akZz5+resQ90jhO03K
1BgxOpxOR2GJr8StcXeaALswlC9ABgZjczreu34ZtrJCCrRnN7Cri4AOmoWFuqcG
YDELQ9CRjAuuTR8zl3c+DEILg0D2hDSU6DHL8xS/NX/Vy0XgSPJG068MLZwmfTzd
fAoYu3egFxVk1H7pEI5yjmoThMphzSPKiMLVuSieJV+kjZ2Ha4P2cP88mHac4N8c
9fUgG3YNaMsDdVEoor+4GgET2flfa3AWMgrRW8aGwCK4FlmwilDg8h2DCZwrw2a1
SVAZepMSqDMoTfBih73JS0lm09d7dGpL15K6Ql0w40V7gdqJTlOu/90PZAmx9OX8
lctNYxkFcAxPNruvAn02zRvvmqbMLvuj8iry36FcevC85vUcEaF6Q/gTf2NbulzU
tTqG5Sd6oUnWC8VxCJMGRPcalVGGeYPZZ+AIMtSo50cwd3Dc//bNbClhqDZZv4nG
nMFoGcJUpwd8Cq86NHYLgEFPUjPE59R7J0KnwM5P5nIdmwIz3vSSVAb8Ux5LW8b8
zw1BqqKD3F6s9R28GjPLtd6gkPmEFDMhIhcG92Zem3P/FpHFcbsI/8qDgkjeN5G8
wXQWOyA5DUTeXH5pQeS3mAdxPQGVq8N/OYF+JCTDjFATdA1bbuZIVw6bKd2Ckla8
zZM20LO0VUZZellFwg/2IVoor3IAfa7gKnvLTyfdnxKSAX1tTo8oiUseVlDwE7X7
Lela2kx0WKXE9HRcktVoCGcj4WDuYxmp3nL25lOdk0MmAQfmtFz2uq9il839nWR9
Ogu+hXS3A2dIhoMtgWUdq6JHlml7rUUNaDFuuUozqQ1QHmhpMBl5zjv4TSaQz969
hk8yxuSwTB+EpO6iLZ83GK5n7G/1meTtV8YTfIP9ooCIfv01jrwQCnZUNL8K0diq
KLpNthes3jPZav7uuCIIuYXqFwLRJGF5k+LJMyLB3pWMg/d8PrH40hU/XZfnzxzg
fC+c1hQowH8OixJHg3oc+UwJafllCQsU0nkDcYwiW04rqxMXcZKzNvjDery1+NvV
M5Q5DNjTpApdR+hsTt+Boq4UyWpzt2QmDYB8ZEFqe7yIcrtNSaVZFlm3F2XBtD3o
HRNFeF+7zFyglvVjW7PkLCME4zRBBIEFxp2CfN4bGs6jaFHqriBUcQ15h3a7yGwl
Z5p1bfWy8OjYmZ0Pj/XDYvxDCYTcN1LK7aauQ0H0PHK1MxGJ2lmk6btEqnCZ/8fI
8/o03iUIXmJKBYQwIbfyYvrsv3a+ETeG5JBqyyRPYdxSzXzNmZcYlC2ZEKXP2mE7
99tAohsRLFtI04EMbBEAbjBgCCETw5fY6WCEOvN2sSQ7QcsRwY6nb2NNjgDEgXQF
ECjZCwSLVzaIGjcZGEGJYxST4FVqX2P6BkziwUm9YjxICamlCytVpGr4WHqPk1WD
ADFIz3P0HEafpDNmcZczQe8L85qYrcx5XhRUGT4GHw1xxutx4dNxR49/54UrdeEh
4FFvwVbPbYiAdNuKBIglDhOtoZL66kIg3FioUvh5O7SZ/V1llIx2TSH9YkHGQ7M4
QkvdFZjuLgtbokjNzYMpdYaAul59Z9TTa/jj0LEBK6L7J0nXGvSfc5P/I/NVf8M2
K2AGlRMdYhnQB17J5OatRI3605e2oeAjs9ORJ4B1OCtv4Lr+qJErZyuzmWkEAYxt
TlfamPQ1jB/X2slNMxx5EDGOt5U2i+PL5E/VtdjpOE2o67ZyA6fDHb9VroOcSUIu
vFsEx4OjfPkrljhFLrGzIZV+lYQkSGPbGvserfauMswfh+tfJKq6ooPka+F3ejdS
P7pIyIoQXjwq8sV1bbrrs0rxL7lxOMoKjdOUQhPYeLcyxUPL+geOzN1nKatEcQZG
jkOjXJxOrdBj/YHz7NXqJtS2u4llmc+efEwYafzbZ6mZ3c+7YkwpKkzUTvgi28NI
39P/IWEIbYgjk12W9pZUVXu3zMwsby6lcHdMKWzhMSisegvcfEUk4lysFc12T5LT
7tSy4mTpQzcEE3YCRb5r/24YgjKhhY4wQ6KFWuZ+Rzb2w7vIeOKRVkSZxqY6nyLK
uMTOeNvn30ad/L85T7CzyeYp5thAE8o3wPRAYcBLRTdR99TWdvQMusPzvyEcehcC
NB4m9Ef4G7bl1p+58mk68lhSMM/WjWqxljOyFjWRbxWttSYADEi2brZNwrDLOVdh
nUlgOzIWsiUsRVoic6i6xnrQEa9XxIkPe9n4Zgt4BZyixP6k7RtI/k9l3ghQCXBV
wZ9sq/T1gtNlsJojX1Ah9/J4oF/lkbr4LSamntB+HaLn97mMH8aNwjt+/NHUjy8s
D3tTqfwX3FsoJkraytv3duwm5lF/g9bMLnRKo9VbVQA3cdt/QaYTBMHd1oX/E+VF
b2I7Jc9FM+7Q318hrsImBWreYoEh8FxdtdJqFeEDk5JCHJxNKN/SIgSyoAXKSoG1
doyEOtFeSsF93a0T/z/Xz8KHXZfIfns1lUMW9ybMRvEyFYX4/LQDpL+x3jDTFuk5
uwp/2uPPBbp6KzcYhrd2u/LnqvJ87jORkc3Io9CJPgGCcOtF2c+5IG4vnHZ2LthV
OnJ90Vp9nvcgejS7b/xkqPYfTlAEY+pMn6UxRz4Xk1Y4JAlzIt8akqCLx8o4mjq1
tdt8V2KUn0aXmmg9WFRMYr+rcBmCBRav5mllSAArhIPIhtv5AaRkHeBolLln3lkm
Vm/FD1ecQkbSVTx8VtPJPs0SuI8kisiFmdUgWKtQaK+pPMcqWp4hVZGbxH9GtOoS
FE4WIeQ46wROhi2+kTkjfG0uCIFgVbnOG6MRvdYwnKBR01huZ9gSB676kWgXrypP
wvJat9hKeTMuXNogj4PNmyGPsAriz9a3I58GblUnQfFPPJhT7/CSrR6nOB815wBQ
M6s4P/xfxO+HYjyBBzK39V2X3QTgT4n56Owe5Z83bhY2DwfQ3YP5iGo/lYs/cmfQ
sMi6c5ihHwQ+iACdfODD7oMtdnXDmnLVSuZ0Z0TVhRZLjdqOQkvOwq9pA5nHvPCs
Fw1g7FXDFx7Ke1K4d+941SOvUznMPh+HYN6ECpSHug4qgXNlTr+nABBU/GuQAy1T
K9fDOgM2Z5lrecu1qdoPzvztpdBjgEDG3cKj4EW6nk5OO3su6r4Ofk6qbGrg14pK
MWTeR51/WudcOZW0T5yATIOX15vRMhfbxJB17K/OzqsaUeakF1q8ZbUQkzx9J18l
KGM8maXYd0cDxH9IEnRUyF/cwrFXnA+9JsLRRvoHm87B9y5HLpUXhAJnzvdluHbj
V1Sdyuc87fb8XHIFhmII6TmEpT+r24LeEry6iKuHqOkBRlfvUpE/CpWmPUgzO1V5
u+xFo0QWHkZRIUhTfMhCe5GRnqlpHQj8HOOUezI+E9UcBe7e0qKphSlVskqHIQqC
l1qIOvp7Bt9YcUftmY4xO6XGXQV6ZuAKOUtloB1ZUoUio/c80P46lEHkgLhlct5D
ALFF2R/r/YXM3FHQtf4FHctIWnA5GJOyjqHO2u/yyEnw8ZiFad6XhAW4gwKxxKjN
8L4h6T7VafI9l7hUX1+6J3/GDpxeXcpgKUSoDzaVKfM9tQX34OSBVzz59im1cB7o
+u8RHS77G9Y710U+IGkzLtby6ANLDzsLsZfM8mHR6viMlEifSeDQ0YLlTCskguSK
VANBS9nYkj9qoU3JDRb8iSKGos7LlFPJydgfBa1Z5+VhQmy9M+WvYv8EK2lA7CAD
kLb23ZRzR0uE3T+0XVFMJgBSQzDzV/qFOfByL5d5cVKYz2HPH8OoFQys0hPJSDSn
q2/iSqCce0hEJCSaLkeiPSvGjJE7A+RUcqt/7j4QZbTbUiDsMlNPNzKkn5C6SzXp
DpqJokP/dp5SKjNaQY94rjjm5Jvu++Qo7X6pQdWRUouVjSf/7AyINXDNFnH3qWlq
VVURuT4gyv/D45sE0hIXntz+0Ad0Nn5IL4/cPnACo+fUtwQijBKL2Xe75kCcYiRm
QjuutF3x0O/3dOCY9hlCT1INUnJwU9sZG4Cji+RLdAP1LPA5KbgH55+0k1FH+coo
UlMF0VlsAKpXmHDClMQ3NbV8HIr2qbExYCAvVqeVthFKaatMCN/48uycqJtBIqfZ
ijguDFxNV1IjspJVjaUVgpA+U5gzugW1NNl8KFKAexfH+eiezNYRhKX12jXyaI0H
OEhoF96iocDIADOxLBK4MCvOx8HZCOu0y9SjU3kdNggZ0GwylHqSDmEEuO3A/1fr
vuBScy/xiVPSPgoIhEnZ3wOhXcjP2W2XERUFLyMQmqnbjqEKxGR6L/WpfFLeSZEL
7dnRwHTpAHVf6adZlKWV42Nk5HKy7BZ6EVPOy55VHICg3vlifU/pmWcfIDnAHqoL
u5i+VPUhbuvIRQW2jTMJ2TwaXpFfECcUoRBjU4j4uuJElHGfvSYA6D/1GnTvKX21
ZYs3vPAh8Bsn1qrE0iTQQOySJaKE+R4yyUUUAKR9wF5Cn0dgmua4ELbdZEYqx3mG
xf65lDL9GxiAaqfiEfeO6p4D8Xs0Oso62MRdXwSy+HuoxLoIXP57C41qEkeHr8x2
H0IpPqCWfepPvAxQUx2wXpfRbmLSzssVMsh/VAJ7n2t7MzZbXG2yzIQioLdG4UXU
12bw7rFaUdaFGMAWjb+DgvE4i61BYSksSey9i+oBmY+yPK7O/tbi+jCqN5QWgT7k
JzzTY7Je5FlqWRZsgEEoX8kTxopstV+ntP79SNh32tm+hC3bDTlCkS05BgTDfPTs
TbbcYoKJ2URj4lqagCkNoQutXXnVmb0jcUILqBBFPflxVVLfhQP44Ffhc7TOA6rE
/Wg+n8QunXcHaXtX6ZrkcwbWJQ82cLxRjTraEYCqXgY=
`protect END_PROTECTED
