`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WsmumAD8NpmzDaMxBkzqZ7Z4wptN/Y4wd+MPca7ZpoSYu3m+qN+Ont3ZNl4aEsJD
4KAlQR4aTl+nWtsd/p/JL1R6npqRWMVGLeJKgmuNH8qFMWRZrAFwncU558U7G+yj
TmsatPmsf4PhJ50zqJHYod0HJ1O8qngA0l0p1oWad9oAvfqSeOxL6bOR4BpzAi8G
NyOvGe02z2ADhQ16Ne4pJgSUJc9IPDnccMLUF1UPsJQi5h7lmCzFeurdNAAspzQo
5MBRfOVNhylzl9emzePu55G8S9IGOIU9aKO08k3mPg6ItdnlDZHwKpQtMIawEYWX
zRq4x8x18+2hQGZqlnNfVfTq2CTMoZcEE0FfqNzY2Gl5R1AfD6h5bb6rxWDBgX0X
7sjysc0FMI3M/Rnu/C1nOE+o7DHSuNZph0+QdhQcOhkOQ4asYEHD900hSvMv6snF
zU9EwfvR0CPjxAMUMCnfwwNPi2SgJKy1nV2QFKwDmra5D5bTXj/XsF/f1bZB/Yaj
mIUXdN2XniOFS3bPY40HSPUAd67o6Vb3Xbocj82k0F/MjH/QDp1Y/e94LtWQCcJZ
8G844dvdtU4jzSr2v9ipAVRu2KrtTRrNWvOAY6DDlsWy1o0q0kSWmSHeMnR9kidV
12y4IHLuS/EQu1zSZzaZEptSnuCqbl6JOsVU2B4IpeUqWohsTVvC68+uUgup7HBX
ludnhmjgr7hNJXvZz99Lq8kWr4BpVn/4GT5ZbZBtBArGUHUYwR211+M+GWZ/4CXv
Dx0eqYYf4+rIvIlh2NT3huEu+Pnh/3Zsyo5eknmhkJ092kPWCVpQWtq0c/nRpSlI
n2VVGSZFvts95cAo9+zGHmM36Iqbqx9XBaeUrTygf6EJ2w/ab5fxF14ZMJXOt56B
UgxI/Ns6pAmOweaZF/eKa7slsbMk+ct5ndgeqVNiugmio1dfI8lBqEzgKDDW5FHq
PuyzW1Te6N/w/kpgQpDgzawjNujLljrvb3/Q1zjoGhkEMZgbu8UqumTNZNm6Sa5C
EH6hMU+92E2a0YtjUCMEJ8qkCckyvljNBdN8Sx7dDcFprHYrO0mcptclqoQ3QO0G
gJdbbfXxhtyhgnWugj/yQzOEMVhK2f7IYqH9PKYdFsPa5ESVIyRueB5KlG3xvKAA
nbL4HPW6TU+AMjStdDsrwieOWKHJ8hfMwDi9xKfsJnwuUA4nlOz2JNpqqICpwu5m
K06l/4ibdYtooNpiotSHe2odsRhIsVf/5WL/zzCvkFGgpHrJdWM4tI3aYFWJwW0v
TI3OR2gHlhteVlyL7OmkJUfopsMEKmvMQkzOcem6Fi1DEkoOx1P4/v0ELr//RDf3
sRevJfL1nGopaiQFLSQ+JTtcbtdrQiKBLuJkzH2lrUYVzmZqUpc8aOhQ5HQzhoWf
bAt50IARTJWr4R6gVSPNXp7avc93oXoPcdsUPd10T0Ylj35TUuCjenSfiVJfb+/0
Tg4iLk2vebFZu9wTX/gzbHOjbXIVp1ErKq5RI1FplYs22YOxePw8Nzh8sl73HrNj
hQPIZqQ1D6585rpp8STcHuhuRkLOnFGqjpMWfj654t4VBjwqPh2UhcQ21WNwGRxD
4OwwvwkzLOoe2seBmHPU1GpD26of9Am+sUQs0CwF+uDU/efOm3jSYPRvZbm5Zwsz
29j5M/KXtk4ErCjvUyPlBwkbNIg1ydWONqXq/BmdaeHDX68eh+AXOvtdJPb3ZvBM
7K7bC2URq/U+iRoaB19nUzmhayPuzo/HgUjCCcs0yTKqWuvhRqSKB5itfirRiqM4
g0AXDvr8NR/alf+1t2IzJJHHdN/+wg0yjs4bGXeBwUdo5bd0Q1bl1qDw27f4Moh7
tbrYJAsGMiweF5Y0MYnSzLJTUBzmylVO/Bd3//jIRFUBV8PxVts9VFrlDF8LT49q
2PKg8Wp9br0J9fgzt3cW+Pcz2VsYD6tqKc/IX/bHm4xszxBiiE9Fcws0LT03roGY
GOMJuW2JKGOFwQIl/RVYtRhmnMZKed5lfBOy7jFbYrVKNvf36eMQYnTVx2uLw8R9
B1/q0WKdch4w2WqxawahzBqXfP1GqiM6EBfHGtgpwuTsMtM9V54lHx+1fAnyPuq4
t+y/Kh7GQaLbwMLgWsQ6GPKoStIiYwrk0gQyltWStGmF7ga/61ovdK8z6IZhB51d
hSZ1u1jMDM4qoog8pSpU1JBH84ivgEuvroI8NiW3wb0qQ3gVCQ9gtfKKNh3rVCUX
FEAJ/KGmxiaJtd7xcdRcFLD/tsGAukUu8b3ty8gy2zTr+sfiHXYsbH12FDiQ0MqI
ttVyDAcrBfY5xx8yFN0BKXW/RSpqWo2UGAlas573efXqkFbL4unmjKglCSzCuxiU
/WboRGphZJERhBaMWNTpp9xqALSgwgNzM5TRp2RG8dLni7k9LEJw3RcYKYSbLUIM
FH/We05SILXwilVxWI1GA7MyOw1vvmr76W0iVDKaQa07+e6BZkB0V20bk8YJR2Xf
Sx8Gtxwznvxq3qiljBIWxQ42GYNuhuZ3N3HXdloIR9lErwm4BwNu2RnUz3iVZOVe
ibYKQJm9+TZUe6GtZNpm60EcUrYxiHAb1rSHNpZZFcqyAlU5p1XqzmfwWscXgNJt
uRLv/cghzJwK/aHuNRUypArLrnupJkp/MBfzTteXT9BempT48rgxEN6Kw9Qk3Opc
VSx0QWDAkUuks1jAcI9eAUP8YpJ4rdv5uW6Xi+ekHNrDUtNp2IIS+3jPoEzCEOfg
AiBX9OT9/0I22sQOJLLX+g240+s8MznPyxHFkELW7CvACAtZMLVOScBzEVlBOzhL
9jd7W2323a3+K7X8XkAjylf2VoiTwQC6BjPJ9lGw0n8KpdFMFEnFKnBd3UDNojed
Lk0eUFczCxiLayaDzaDH3siK1tsqzINOhzC04dV/Gi4St87XRMGK/NcmqTKNQ0tM
4fMhh5D9SFYCSn7sBNm9osU9Pcok4t16d1JgSTgsPNbvbCeUFEKGPa7iHbKrro/+
DdDea0Hiy8n5gxkFR5Vy89V2SLqi9Mz6+jrGTTjvYTbkGXOLFqdk4VKaL9bgl+0x
1frT1BMVIr5Hk9Ab5ZZox8XvmQfBl/Yf6SQomQWwuJt9rI1mdr/Ymz/7/6V3UktP
+jPLUh/4RvPd4kLGws4+1DNXazwjzNbWBB1B2pK8V+cAx9sd3yh8BO6EG5WmjpvK
VyWrZQildJWiNq3xT9o1UFS4IO2VASKzcWQtovG/yPZpt7WfGklJz4Q55kWXay9S
X+HHM0W6a6FSfqY5orjFt2ew8f5T9b0sdKTVTd3piipoRr9ypDrmsjp27JveM9D1
ACQB8tGJ8nx2d3gj3Ya8e1KpanE9SMpnA7MmU4iBv6a3PEyatZ9MaSp6uxEskAzb
BJvX9hRNNwG4gPaa+jk08P0XmhFxCAgVA1M6Cp/fAcqqYf2sP5mjQR5ztNZbKwE6
n83aXFKl6mzHd6+6tQ5AAaZkezDL5TVIY1QJVpvZvO+Wn4Crg+i5X6R7JcGD7LMX
2bQjuJgHybcnzt9LvvyzwR398NAgV5Vyyg1bUpm1QZDg/PmW4mGNHswqCDpAI+qM
lcIQbeNllUqczvqH9uRllzk5SriBvgvLOa68a8lyW7m5Asw9aH2oUO5hDBzajXba
+o4cOj9WEiikvOCCxzD0JyABNrJRdy9W6OTsIRAYXFctK94qwz+fWIPSfPxz6Ipc
Aw31Pna0P+RwMhnvPBrz7I3jNd0ZHiCEbOTAQrRSqgahzKfh1MfsEB8q3v/cF8+R
uy+4RZAXecDw5eml/WjZaM08XrfYuw6XkvEXB9XJia8//WBN2APCbi3x/JL5R+Wi
Q3MRUqlWojBSkPAk45smsG9PP+LDjJ0fF2PUSrgb1jJ8j4OzsoLsEaIs/nTKjnKn
VY9TMWAU6brh/hC6JV/B1FCcaVrzkM+lWX+vp5TEWrTF0aiMOZSJDyXWz9dpwooi
JF446/jSOm58H1IusrH84uHIPQOWDm+grODKGSAAsDga47w6z38f8Mu8i8ClZn/y
DLuTxfndif5E7FiEQzj87TtOKnJ40pg+Aj3xmtLJ0IQ1daTL8qvFOGdcIhuypSlJ
G7ODiftQjJX5789QyanJuR+UuJr2Jbb9f/Z7GjjSKd7d3VHg8zDbHCn5eI0mA2HM
Cjixh7p6v4+4xzQjrqsaPUHp3Zce2QBlzCYUMkV0f4r6xV/Z85IgRE/Ps3S65AmJ
oEyRMa8ZCAJunbhrCSjOrOtzfi3KDwz13A4N3zzcfuzmfOpfqA4ZcKCRYL1aQLjl
eS0f6coNx4G11LR0wj3n4v3wYr0ZCOzbUaEHv51DwdPlcQUX4U62X/hCJwM3/fuV
mrwHLh4XGDk7UsL0UljGRQa0np/6M6EfT/Lg7eyEixB9aecMXKtS62qg6LwhlEYg
27voAUcW1BSkos4WjrPP3MT8lDMM5x4mWe5BvJGXdEGZnF3wR41sswqIzVAOZI2O
ynBserQHqyq4r9JgqYuFC1QGNwywDCuyO6Xx4A3wxss5s1ogx4DrqV0BGUDNBzKD
VdpT9mQ98p3D6r5BdTaeIAbSTavP/rj/NgXIDtChKVPPoMrEfulj3L63eNd1XcBs
Y+PDwf1uze8cPn3+DjIhrw==
`protect END_PROTECTED
