`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BXjkf97f/79c4H2E7fpvI7T7Sd/SozmaDClFkyJm6JxbGCPHxKIHVlqooW3mUPlG
xCJU3URooPwwHersRUvQWsMV+uppRRPRFcduOzV2hfIRA8BRePS9P/bIer8kjAiy
oOvjhjN4WVFWOY6Y5OH0dnIPZaZJkDDMtFxHTEDjvRGYztoemDgbiK8bLwkz9cox
6y7jADKueXO1ulq6TA6g03+mNucjYO9svo9FVBdY3RNyVPQCSoZ8n9VVV5B6wWWR
CDgFOdjpx5pJtxnH7/QRAR8faKU5urODsPvHwBPbJ6nk8wHkmoAeS8fhrwyNAkGZ
Ht8cEeBdo3Z+yjMwqqQ67JVBEOUHGnTdCKQgaxOr7tv1CtqV46D05b2wFXD6/IVn
JTcSHsxfA74jl6IH1Ugnq//dB0l6gc1JFj1aBEfggkltJfojXgVD0i1PXbt1j/Tn
kPLYcDLLOa8nXYysqEFyjrsruVPRKwJGw0mo5KiqTI2jq5xIfn6ZpniaFaO1/VE3
TJs6C68GRGcLutDvox9n/losff2LoRAIBmK3KbFSQkQoUCpuOcvb5yIGKU4aXVBu
WMT5qHBcbbyq/C+wwTZWnzEmJ9JMfyGUFowvug0MtvgXR6DOU7KfzPn911hJtwcM
ZDMC81sCZqaLg0zv42GbTRi5TiCnZP8QlvLBrrrATXQwYfChdTRdCzi8oQ+MqAUu
vkT6ijOfdVPzffLnGw5WKQICVkkP6YZT1E6PrkY1gQhimkkSAjqBe6aZyxwVlgDe
YUwf7HmxT4UgvvWdAd4G5f9mck/lbTF8lZDOOhJCdjefYKA179DRXdfnc8udjaVc
frxyGovqk9ATeTTUzOCvk0n9GWx894Vn4ftQYj09QS/8LaMXMffAd/IjwKeRhScg
+pOc9C9v/Bhf1PdLj4c8RpgbBkvveO08EhLCfID0VaIvf8PryqKXkhlx2tC1jwMS
Kv8I+RcA/RoZCXYk2TVQrIn8rKUKIPeucw8qIxjOkVHFuPgzcyuVCc2xwLzJZb6i
pjVaO/rN7z7P4x8xziiqufSAuY/gTe9CO76Z8Wg8E5kPMN30latgatkTjPjZvA9J
hbQK4udlXJ+3kQh6LhGT3otMcy1bTFxpjBvdh6fAec3onJDGFowGGlUVJ7hf5N2l
cTNCjxafT/DpQj7e4eVtLc22rCdSlOr/imEgD5xRKFD4ssWTJ0ImXzmadx5Q3rYe
GmNeyB2OufkgTTY6vDvwLw==
`protect END_PROTECTED
