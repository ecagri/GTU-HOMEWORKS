`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8TqS4mMZSZWIyduveBA4r4oP+Y03pKSCOZGcn1llWXbZVuJX2QGcPP9Ixf4NGa7m
35BcwTWWE9bSf994KFCxfbRHs3jJDA1Wrs3cUcMgb3ZwykG6fLYqWKRFRZoXve8T
AjfzzZwUSjesL4EllRt4fWznOoVw4nlqm2KbLTD9YlUqYCcqd+ZXexcO7hsS0Drk
KLlGExbBuKDFH9a2UCoool/SBcAmgMkM9mWYej6JKglRBvO2VblwSq67sdlTlelQ
TgdPOk53YcSjhb+XqyB2DyUvpXXEL1uhvpULWUzOnzK4tAc7P/FqLebqiuF23CNN
AShPLOHFLq5VIROOoq0WuuEkQsJ14t1SfVnRIEsAR0TmyaGvBFv1RF/YsyBrOqrq
d3rj1w6oEM9k9AI7UkfmAqm0c3j85ceBz55OwZyX/WQfhb2ARtobb4mE+cOuV59h
BXxeIK7gbMCaT4UNAzZM2pN+cDRcBNCy49rSSkUR0wwYINx0XTkhKAk0bwiBUcs+
Ud/upULnTT3zuYxTosQZ3YFcRd+jayMqFJ+GRlnHLuAVSsz0CikQzm/B22fHNe8i
UOp6Oi2U2MLxVtwrpTXvdyqLDXzvnceiTkTdgCXtuR2Ikn1rn/Dap0rJR6pDHISC
bYk+4MvkVGaLIEr9CoY1+K22tVrhKBoATagKc5jZQg5ny41vH7G+tMGl2+nV4idt
+EOmERfgi4OTMFmvs/dnKVyMbiR5uO9p8bZJAwtgb3LpsngXwlRaiWSpBGIdhUG8
mytpudT1Iz47cC+Dp3sk4V0e9GJpd8z9XhGxxE6OlpsPGTlCg2W8CfJHVBfsWjq6
cjTFjrKOGvWLYmZ7LxVeh5BkQmLR4gVNIy3f00BmPgB6WzZcp4QfkHYjgsgWtmM9
Ce8CtXKBd4RAbwoaOer6TwRcM0kQMY5Dp8Y7GkVrwEeOhNVcHidyVAw5aQuSaTwO
Zn+tsBa8eh+Qox7hgWM822Nhp6B8EqyjcwVdZ86dcUyML2Vj2DfI1RU2fSgzwjeT
Zp4qVYwMwMnsJ1qD7c+kG5yKfxdq9RKe1skPLwqtPBJbzdfSA0EPqASryeyP83fz
2Gnx8OHdcERdhIhoFy1tYoWv1ukU70lmADEhkaPR8aW9GSEJn+PGMUOoxv+ozLns
mEseblkqf/o3VIv91bcjYdtNHlM7Gaqi6C4PfelN6qMW1kyQMlScjd7W30kz/71b
EOL4igP5yMKcVmIws2ElpoQ4ioyd58G3kyrojqzUm+/OrmXTsyOxl/yQQJ2XJWEQ
PREWEuG0aKu6Kzx8B8YxHP8heXIZe4ZkcG1CyTmHOC/tcN/F6vCez5WNcbfg7XMi
AF0qceP3Xdmi1QRhiRyGU8FmkKBE7CAXHBT4a72Sycrw6I0YTZ7cdUK6/4w5Il/b
i+KCKjANH2JYv/aCWPvqrdbTKokZw3dxKgLonxl4K2ThqGlfiX7H2EoxUk9Dwhmc
1Mp7ARPI1LcfceHTIo6cdrZzumcJ9Q7vQOy6u26/AzrYKOY0L0g/GpbVcUEOxVnj
f/R+X32Wvt8bqje7Rqe5HYjoPnykkHxzvZtKF45bgM94blzFJ5tZI7jtPPiuNF7F
41PmLK4EP4Oxg+eDY/kzfbl8qo5AvNpyhmt0VyhZe2aCHFTDywJbEZ+30pba0C/+
YBowISxOrl/1lTBwPMjWFmOVzniLgv3Mgsa6OMaSExBf7zgRlr2Q/uemlLHTdomJ
3CrsNOTKmR+dCXH5jHH7cqnQ+Chg9MOug6BV0YAWjOh12yMJOpDXxLRSKOrzK+lm
oE3YzB9SwkJZnYj/OMO5i3iX1Wx8+EHK1er+ljCGRqMpNdxZTqw2g+W72WL/4H+f
Z9ksa+1IsDlzCUKg9IdGrHqz5TTYwaMa6LIQenvd+vcawuEHj64lali9zlKEHftc
lbmbwIyUTTlU2moa7BVS2bdQCDx00kjBbhwpl1LSK3MsFMIrScA5zBAhsIw0z1e6
fHv+ZgaCwjMH1vHxsMqoFVbwzWASQt+5KYZTf1qo64JAPmrbfJmXgqb1Na1A65BB
rXn1BncAvv8eBJhPmT5XmaEAOuu60Ss3twHkxgYTNtt4NxMGuaDjxIeglPMEYKWb
BNTsBuOvqzc6fNTkqD/OxL4FF/oAeN6quPLYFv0/YxBaVptmOL9ERxsdZkht0o2f
pUfxp11xCNkzsKbpEOlWQUpYLrC+RvSLC4ZuvNXEe55l4SkdXi6/jKHpt03hoHSm
64zeDXNQVxl50bfBGzJ3AkvZRVv3hHPRO5/f5HmZGn62Enrhyl8VtmFUJHr0EoKm
u7x1ZYdXsjjixE4oUPoEhfwyUpINjXjnTt9dGH624jD4kfR1fhVTGMrtsh27PSFI
oLW5g+rIvDDRLaODa/WNjrwdQS9xqcCWS5LEKtH1SMXSkMQHXjfuUmE6bdlU858X
l7yQ93uUrJ1RjOP54fIUZ+EZJcis+63ZRzspvUlx9lCzSyHB9YB7qpzmdtQzBJPJ
PeBGNIBPTCGJ3RNpxjUC10jP6p1+YYOk2wVFNT5CxZHkVXr4af3tiJti9XCJo5YU
jWyx/GhYPaWFWTAeYVV+7Voioie14CGnhg7IaiRQwYCPoJMbMlEHEuyjefSvg7nx
3AgueMyX4zDgJX7ZBaPEp047EcWslSx4kF80Xu0tZxoy3PzAWgPASOVCKn/3s+pW
DI7j/iVj25OOhxA2HCgh3OdbZ+cgNXet2XL4XaaE1Cwqsv5fZKcSl2YpvJgz1aJl
xIBmmXNCmLDvpvTBQ3R6QkgJvruMc6rMmHMLDEKbQpb7MR6SOgiFP3y3HhoBRcsp
zvMUF0LuoVxXd/2cx4naLUnZHMoKVtwGpRQN3zX5iufd3k6qRG8Zj/pBA1xHhzRl
m5cMBmi9Yfl/xFNS5AHkrThDnIXNZNLnS0KlkVcCfttJEX2FakyYQCbLVNZgz9M4
QjnDkAkTRNXFX/zuwZr1wWYGP/UATFIwa1xfDW3hGXTI33sgMdH6Z8pFENvpHZpq
HvlRk+z+czimidqfp9/JVLkQMYGF/WHziAi/mhZw+MhGtlzfL2z2lIx4qdte5V7T
xomFmLrR9OJ1yPjuz14g3mUVe/iRgNCZAeqZ0/7WsDzooRrylDYNd+oCz4eJr0PH
8I9ljRMxSdFBLzgsXV4KhpvQmkteZ5rh9dewy0bCa54POzz/fiINQfk2hvekGdJI
hq6fHs3H46SBrikJrHGQ/4CGYMSV4SnZxGQaPNawVYq0vSpdjobKCDbdsYwNqY6H
NLqJVL9mjwa4Xd3r4ADaDGk/FnvquV66G+NO0gGIa50EeV6SecIs4W9O4MBm/nk7
0g8IKd3ZkRTLSSVo83ynRZF2OXiMzXfbBecYSJvUl5+qCFGkNruMkjsMPhztXHP8
dlqFMlkziUyZhy9RSQ20FG799Hck37IFeE6oXDC7dhMGcgaLJRbyts1701TWsnPc
Tp0s0mQ/luaM1dIxzHdxTdAGBBg7nmGVRFnm0z849WpcE8iBcvCkw39ChbVHlj1+
fRYirUsJ1Aynp5roTuhs+veRS8bq4bKIw+v+JMK81pu0JtL5omqmDE6h6ZyuyTOx
c+x7E68AumYgZr8b0MRkrfkotCYmWoZSJR09XnnS9NQ9CArlwJDRSYmpAO6HYndV
8CCRGEWxy0IGa3yuRGYDdWPw2JtCaA2RD8uK9pV5G3VawPlXW8lSygbPAZcH890m
zDurAIACbrcoBTZfmFnZk6qXH2nTWYswlnfuo+n+D3Ti6FE8/VLIyMnuZ+TjEJAF
WAJYMvT12REjy4B2Jn37NNSbgwU6HAcDg4FogdvGghX0Y2VHGwZVgHkp7N+0N9Ai
O7Iq3d3OLnSH+vg7Ufnm1vEVSyWtHrn9jcBz65t39KCIjpCdEJtfS+VJp0bBgJga
vLSrkiuvt0GWgrH+MU65ahs90SGKzmh3pAQCNWO28+y1VdVAXRld7OLzzMQOm/qN
j02Mp/GYk3ke18J3Gk56jmeArgwcmzLVM3GjYnnRyge+dCFaLYv9DJTXosnely0q
Vi0jkh/Q724+zymybbnB70sBZ06OMesMqGn+YGb8ovv9yaVtbkvD3OOqZuW8egtu
sEyroZF7f2IMtYbJgWOaASBHbqrA3fUZcOMSbf1Um5C1HPNymktYp3Y2119KPe7Q
JR/gp92uvsrPaodp4VmPSw1Emji9K/CAupFflm7a8GTzffo9Xt1iISrjSorbUZq3
f8Avjo/d2iX00LscGjqOG5wNhBUNMfGMOg4tdAHi6GNvla7P6J3iHIOqHQhFXk+9
7jZTtFn/d+gM0rnwG0f03HPz2C7OQREvLIP8IhQ7gLKZjRdguD15HMWetwTfHIif
hWhchXmnbn0pEhsTKZC+GbZNM7jF9RkdpZEyzaumTZZLZIXBlymSG7LF6nSEETte
2TOvO4nKLp5t5V/5zN1+6qfjzVY1IqjVF5tQ1ZKVAdwJYnhH0F/1k3QvJU0r78gk
XkAQm1PWs7W474vTYF1zBKZq6C1hdYpPdI8dpALTAAZw/eZDoXSaXDsVl5fTVK+J
ZL6uug06E3ES0MLHm3yjUj4dqRTlJ5eK9ZBKAmKPEY0aIHYoFbbDEcDuNI9MeLIG
OldHg4+WIiHjA02NUK4w30fLsTTTuLuTA9kakUD3SpbxpzLBBNb92P5/lmR5hfQB
uCnbTwc7SNbBj/65e+JPQkMLSSwe/WwnjLQ+j+kFkDR823SxKBWfPN6A8ZeRS8Te
BsdFxf0+giS7JlWa8+CHWhgu2H2O7C4vU2zDd7kMFwV0yh0jjEaN0OygsdqcRkIK
MHV9zKvnrDQ1xIACM1DNsXPrdesgqILeXKlZJE5Rt6PcibjnWtJwOVirjyIQfIRS
YPw/rjKYpRnpc9jC0gef0Y5ZcOZ+R6ffGiOVyzBCp1+GJBbgUz2UWXyULBSDj2aB
Flo18NyjH80Oq5wOigj0e0CH0RVS+TsgmHoRkQP6Xre0eQU8KfIQdbHzl+kxAunL
+JzjH7QBIaLbBWQjXrPQnF4SSeMw9To6Fl4rPVhEA/2FYNyrDUNMywblNy8RpUKe
CHrY4Eo6fiFkOPDNwpiqNrvNXbQtFVCOZLSMkL5L4N1HeeiF43fx3YW+MA6dXooG
Z2xgEr2oT6FOdYzgHW0ZfcaqBTx5SrDUJMWtqkKNaMbJyd6LaJfRt7pAUt0LTzsf
3eBvysGW327B7YJLrZPhXwVSv1zaCDfD2TMYXuOM1IQZVhutQMIucXtiqwkGPAHi
bqmZuIykJqEppoLsxFPgSl9aTtba2BR3U02Qh8At8GS2gwwTCkUqwIOy9uVGnX4z
78qTBTS6yZ5qvW8tbNTL/89KOWqYZaEAriQEKGUVU7XrH1gpD3wQoETJUZzwcpKY
trOEoj8X7VvU32aC9UsU5tf0560M9Rg4EQYb2UoSsCXBlJCv2e+GrNWFsnVoq56t
lOawILk8luypWmxUQggPKbtZYQrEPgPmz5K9+43GoQCCwEH9m6D+1dUSvlNFb/Ki
XQsWoop30Ve209Yy7a9ilFGN2URN9fMu+uIVxm8+y7Hd3KSvJbykIpo1sCT6V3ag
nNX8i8T3ca4GyAPv/w/3n7JAbmpsg2AABLh/BowJyV3SVbPp/0AvR4BFoL5Si7Fn
WkPyC5nmB6UMT0kaFfU4AvLu4yPDwKl/yhJEZ2axtY0EQ+TvPhTiDaBUT4mCHr+1
4YXalZgZo1yOy+bbl1ta/qQcFo51TC0ko2Tv+3r47ZVC1Wxif6/9IKVpSTYQbCQl
bhmHYZ+TqaAwDSHW8QzSdqTL5KtImigDaYGFaC3mfGw=
`protect END_PROTECTED
