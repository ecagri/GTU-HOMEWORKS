`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NcfPKvdVvFwJze7ZvXytt+W59RjDdwCBZ0tw8KVTfz52Re0no8HcCIxkM2E4cIDo
K5YRpZUUz8du0/nsho1ckc9v9OfHlwF59CQll5bMdRiPGcz29wkjENyFzj5kqgw8
77R6wcAUCXNKswqRxONUwVVRvVgJVWIAeHJA7LcFOmzuMXMHXkCdKUo9zxquMY8c
n45AabzR38+qENNhYsuYPATrhK0ABHzRrlZj0j5liSqXG7fzgDl+RaGCVQhsEsE4
JDzgjT7+NC+70hyf5+1Ghv49Vx7l5phi7ke0dYovq9jQBHFCwwWjwmjcIsnIUBd7
4rTUF4Cvb2HNxbXD+/LpmYmWE+KQXGcwTagL1yIJDKTHhesZEN61Lo9Reg+YrJ0i
6P2VISfCwkv66WSrVHzNn8itiGJDCX2zAsNo5bhxFKUWI0beSSqdnsiYJr3uzTgV
`protect END_PROTECTED
