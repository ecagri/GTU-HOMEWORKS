`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QfGQSYOSbRET3p9b0aQEPBFRpKayJy9AH+OpmaOqCa8G8yeewxLgGvY/NOjRI4uu
1u5HFw1v69O2AE5GP46bjdEsYAywGQEhifAjMpX9Y3/z/eBoiJePdD9rpxk5KfMZ
z0c/Vi9fuFoC7Oc8CJdB4LLr9ZnKPtJFzWPSzDWdITMGUft6VBiuQF2iH9nQ1w0q
jjMXd0itq1j9HyhiUY83kxszneAKy3xSVKrYD3YntmbD54xijxp+MR6HGZjQo4nN
QeAC7qP8CUZziNOIDJu18uPSUPAcuzSFYwl2GHjVS/NbcqFkCtGXQIHVsAainMEb
H69coQJh8Ly0CBwwBxju1I4HsS5IqPV87zeopMjI2Rt9DJNola9fT3GKzmx5xKWV
4HrTTOj4w2qsAmTR/Cma4YSnNa7urFhktKIvtEz1K0X9/+a0rrJ/P8ToWkrxO19s
Ni05Yflb2p81wxR86LQ44Q==
`protect END_PROTECTED
