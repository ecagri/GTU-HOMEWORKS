`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BeqQqMxtPwnZU3Poh9O7spHB9w40PhiR8j9T90xeZVcHDkQX4I0bmiXiAFmwQROL
hc1deJQCauI9R6IGlYy5+7BCcYMZjDIZlWAwfw6vkGAHFLevS4be6Jxgfxxc27s3
NfFOZxbmPbLP1VY1jcKC/ptGIMeWG9HG+s0rau+MtenF5VIFYEoUeBsF7hIdHKPw
mqeIeSpfCQUWj/tAEadKaVwt4BOIC7UBvxNSGnBd3Vj97ufdbJqzB3uMj7HzzXiT
KbXgtSfTx/V1teWaKLUWFmQBaB8z8/cvr1P2KDnNUFVoG3QtMN8mE7XqSTP2MRg7
2Bxs3JEaQZf0TKnOxn5angn3m3BvdkmHbToiaZ8y4ZteSqICAcBk/zLKvFdnI0v9
FEv+Xn6dLn52+97i9mxsyT1mOLCQsbgnmTdvJDYO7O/TxHLbVKDK5CbW7Ocwr7rm
d6hQxaqy0JNm+HlH6HTU6rjHNUGoY367ZMvvm0vCg5jHDfXU2X0vYAdLmGRteKd1
nO9prgTGrvb6mpVklVOX0//Xj0BfyZ6y1TIIQ04zDbNzg6uPY6H9kk/tSUl9gtY0
HMN4Lfi+AF/NFIT1kYLIrcFBov4D5Vg71T7yCM+ZfUysCAkHCv+TucrzQi+dukmv
EFeVQqK+lCUC2JK7O8n3ZZTxW+et0Pv2vegDFC1I1hrYH8uhC0Y4p7FQYBSDJJFk
hIO1KA8+1ln7Gv+b+u6XEElNnlQbnLcyntjlw7tfzryrpanXag5iTL4KtuVNwlDg
e8mqdVIpN7dbx1eLc4ANV8vvgkKdX9DN9pVLnHsP77w4x5khFTseZ0NacmjW+6Mk
5WyEAJOb6KNq4R+hNadHrgUipVMd8kjWsmCZyR1dJP1zFEQxUIqyV6ERqyddTAtN
e5A9DLLlJ5O7d/5iR/1M197io54U20tDnPAs5cqqjSdXGuuS87XcMDv56++/6xk9
QG8dbyB3R7pqXHi1o7tgSqG4+tENc+4f5VC2hVQPL15LxILBWu8D9uHu8YZINxk1
CT61vq/dkrG0ufmSZtNRv3aG2fmNLFS7VvZlJVVo8rczKGWgWGGxsNiNXn5VubgW
+C6rT/kjlSDSXu5w6pqaFyuUIhV+xFZd514sxCmKHhTNxdTS0z5Ib76iyc7FzJ6e
TdQYKeQURiR8RkFCrfmQ0hVNGZ17FXUEFqkXytFRHviSoamEiaQ1Sx1vjctfx+nA
SaYoCKwSteXmqAosc75D0Hn75HO4Bk1ipNrubq0MlxbTcg4z4AeDfCAM5aU5b0Un
OcH59RrN+6fNfxY+uSlmlhvbCr2EKa8Fn7F1cCeQShP5NFJc5u71tr6AZzBbKuWH
3enTchLj96Z7gmAf+1tCXfSYlvyt0JFJXkDEFJ4OOkbTH445HtGgl3SHMTr4rkm/
j2PydWrD5AiMZAXUuq6BVxFRAVU7rJIOFkWUWcLYmWrMqgj3SYpeSjjDQ929+RGx
UvfkaT0KfTMTIPx6qYXVPIGVQQ0iNgVw4hcTvNjzaYCd2nla+mQ7feyPEyQOc7jy
6KO0qVs7jB7oyp7Pn8bqu+l/6EouJ7YGp0Tl1VUCPRDisdE6d+CP2gyL7rcOTdwR
nrJ84D4vfjf/mD9RVUK5Ph8Mq866RfOq5Z+ofF4Cv30FdDunOiflRz9+yJieqGI8
8P4zKwnv9f7Y5s0l9b3+rcymXhxcZD/ddFraE3gWCbDy4nKW7RhKRgx9oupGQXIp
XLNkIaFsXWtXBGp5FHk//gEWeIVCm5bULOLrObFFzZUJYGsC1ojV3PKIz4ZMw3mh
aIJD/sx8ZPhkGZ7TtxI5valAQyjQFDufmU+RsvPQGuVdea1yUJJop+YZ3Hdu7rer
K27A0U+YTtyaFQL4GuRFSwBBgytSRxSXcFJShOywZmNLn0Kdp6t+bG7Sx0r183J7
OrXzpVRXq3w5a4FLsUfFf44s3LiejDrxN2oPQGjXyhzAfX0l1kNDiL4EB1yGeI5a
/RYmJ0FHLTmnZB9s7pJ96lEh1liuUh4cCfMWfwRBKgUNK850+L4+Hx9hNIV/xjTz
1ACVVvTojLllfpkpNzvToEAi+dXltOwHaRyPHJ7q/HnFNbpsD2/8X1obOmQE5S31
AQUVRalvyW395axYXVKXDJN1ztz5NuXklOwN719CzlRqvBh9P30vQ4GcsH0Ce3oZ
uLaQ7mAK68GCClNeUnBPaxx/hvBYiwrvDjgC+CU/yLUh3p/L4qEKUeT2985ynyO2
OAkaZBz9mFzc70lZfmpp3HVIXyCtdXCH5pM/6tc9wU6mpfvkNBro7Y/FvI3SG9uX
rIxM2FjMR27Cn628VJ/PGLm/PANwOQkoQTAYQSW7xu8q5Naq3j+z5Gf3eiJEmnCw
zcJzDp7BrG5+7F/HDvYicAbIMsKs3PUqJrNAkWr90mc6zl8ulcDBVEcJBXuB6JbC
`protect END_PROTECTED
