`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eo2O5xR1KDCxkgy1KNpUL5xFkK1GbYV/hLr/7k349m9Yin3Ka37qgE/iosOlLp3r
ROjge3HdpzhvEQFXwpkgF5NApClwwf7+Bh9vBBlUiNR1gyPxWMd9MBCrd9KGFHJd
XNoL1Qt9gEIjdFM149Y3meVLSFpcJlRAkeR+TAIB07jUkrubcI9lV6VYA+59KP01
KnXfvcH4raws/x87Y26fLD88+NC8BvGRDFwL19ZiovBq5lYsyZ4OBPqIAk9rsNpA
lXmmQoRHLdAnWhsN7OVzuS4EPnMVEdfBL5nvV20Iv3OmxMq3/bRHB+DQPWEZvK5T
l/v+mtIPyQkTJiC4tQjDUfRp8z3e+IMe2EJ3T+dUMsF21DyNktREoluMGOakTGrG
NpBs0eeoI7eqOBTE4yqWB9i2wiAmVnJ3ye5c/7LKExhJIxmo3nxxFEiHpbbdl/V9
CyDsbMzw2rvjoGJGH1lvE3HBztQigKlRrXX8qApCNMs/LWttDutXGe1tl/94LaUQ
0pZ1Q3cbBwynZR4hWH0uUSV29rnKzdyhsjjXK6J7w/BbQVqaQxDWHUSPJ/LIMq8y
j1qDOPZ2k719Suxjr8ujYNxkyiQjgw1nfZHczJplBNiJqjqOjQYp7qzaPDjg5Vvk
Rn6t2NKFxbvqMHDHUgTax4TzmrnxCS/LDYNTvJu8D2GARlD4+KmUFEI7vYgOK76k
ZKdz2sdug1f4/f27C3DaFDQOR+y/tHGstHJ5E9NWkVX+C4shbsWPPXGc94mCLoLG
15Zj5qlk6biXWr3FMV3teCjqgPn5+3Fr1XANxhfkAFq4eSHAY1WVszGs8sllfgOy
ML55sBOQXRMImW+os/P4X7LQuDTvBVtmAT4sP5gusAJfxJT/4hyZnDH4QPeQpkIR
/oqJa+OHU95IpN9dCjLpS1Th+F7FBSZQOuaEkx/DSfR9R8+Aabnn6qZ1jCfvzub4
EfJxicYZmZFdqXeChGpXVsx77IVDgt7gNTdLCcAwmxWtp2JyNbBsItuXYnV4d2Im
bYJhlUr1/4Javx+Pd4CGvSe9gFTIInuGFtjsmu2YZSKmuc5ouhF6McM1BrcMp6bW
bxmVwGW8yzeZZi/xM6M0BaK1x7L6fHH5gIrr8yOJJX07zvkqhilh+2TS/lFTlRMu
ceWiZ+RDZ8XaHmn+rVZ3CrV/7yK2H78Gi4mkKzZI9NeiCy0kNEgbk2juhhUHEvO3
wN+3He/XHTx+wY3SEy8WdMm5f4F0WBNeRVhbz6UBpJVqYL/Px+cwNeYP8+QFDhjT
G+/w3vUflOFbEEmwJrfWHx8eLeer21iFzCcI7HOunDpsIxuYOlnAibMw/gQKI2gg
N8nwQQDTDCBzSK9Cp2VZnTgzB1cGAEBQVDxdlB+7fbXDpL/ZG6WPHolOfXtUaUzH
ZJh0Nak97sts38Ii1iHCP1/AYMgUjnxHHiOflbTfn6JErTX/XE52PHR/GMN0Dszx
sDfkESavF0E6zXP957Qdke+8bYUajvGuS+HBkV+6W3Clx8alHM36a7m0WJ4Euy3l
6LLUqac+AkrJuHZfZehqeqT7eLTm6F4k9A+Ij8oawBe8BMs2FrpLzYrkfytwzm9f
mOfj7uh8tYG2Zr0PQoRZI3ii/rKgc/zGJZ9kaz/TxS4bq2fLdv0LVLyXHoexJ47G
7/OkAb7S98Fmy8PG7nzo64DjVo+2ctNV5UR9QGAPjiis7FYJ/QLWI/aEI203S2DH
/VU+gW5igBDd1JRmrrrIhmhDJWXdW5EIm2Aq9Zkij47bTp4cx+v4HYXB+NB/Vz01
ub/THOX7Pk2Udc2wBj5wv4UbN55YU96/lc1bzqr8YiJD4BjX5T66ojVIp1NLaPfv
gcMQJh/Gh1iVaFyTMCRI8OTLMJcmzc492bEKz2uXZBUHcloHxzYe5QPknTtDFvJ7
bWCgfo/qcPAGMgvgh2yDcW2e2nkL+xD7M+TZC//Ou1aPJRN/6bwPrB/2+D6cH6V5
2kCNod1kYiKDjeU2owRUumQGv/SY7gNfPZISkxe8F4zqSq/Z/yhn0W6cTEZH2g3+
jDvxG5pUsNEBKQRyOMuEcoZ217c9y0Ls3YAU7SLoZJ7c5f9XGcZ/5Lwm0ISGRyGB
DLT2hsg0wbgbkoOCEz26sN4hqdKuQYzXD4MGDb7t93be8VkzQ8c3UjyqECM0cUkR
bMO7MfDZVJ+EhtyS/qA0u9NxcgMD8HwrTkm1rvk/sWPEL6jY+cCvPV4iPYPOT4g5
uV3SLwS/rXFjvSopTJBU8ySQW3PK1Deo6lg7Qe8JXRl9x8ULGHV61YC3lYHhgpCp
S0iRv7CSy6rLi70Jlm7y/daLZBaKOXUuUT5ZccUTWqofnCIT5BwrtV1fVJQ7Yj4S
DKf1252IcbPt7UjhWuu0HOY0sgqOkdgePZNqm424RmltD1UxEpE8+Ax5cWJs9HAj
6FW4VBs26G3v1vVAp4eJW/TJGE63cEqIqDf2CT+oYziS9rTqzJtPphKT7WRWg5i1
o/VvhKiOollDtQ9sJ0xDm0AgcpMUnbBL/ThFTTZ5VPuIHEYZgxxbQuTiogpwinvU
lvB/do9UMLArZhb62zIA1UKmeUYHv+sz5ShpBkTtKfiO+ih2KbKYjHKoYGrdg2EC
ocraDAcjc00USGDukszYxWyy8ARpRTujcvW5hcj6ota1D1puuMTZ2qMvZzGXoUrj
zzFbfV9G63OyUV8hF8St3GRm/CI5tQfkzCG1hZb2KjQBC5A0M6T0bOxMVzUJg6yM
gVKSZ9W8z2TSB7052PQaQ/HBNTpBeAzdplKd9cDSkmJtR90fxUceRIx9mcOL0Uqy
4UCRVsGzsZjX+/xEnjuTBNWfa4hCQBddWevSs9MKsWdc/7RjlYor7kXNVhIZNsx4
iqA1ZMIi2Kg+Fmo/D3wpYgqZ81TYQ5mwd9vDjBuN09LdkbAdbgqEpfNJvfxsuss2
gqrlhD54dq3GfGwsDgQo7HzeUpKbna6C7/an7ngKHVnhJd8U7d33CL7Nz6CZhDct
fCnG1MijcBWJ49KhCoNUkatrhF5PTlbx4EZoaFj1IaXQ6IHGkJGAWXbynHVs19yV
caUVy0/ItYJ/B9NseWLFZ+B6XsZSsZEOedDkZcO3Qm04byW03HqGDXzkzjvM8ML4
fuTiQ4AteRDZ0BFie425+lw0MBplVY3p5+VSgY2xjwBijkEnb1L6I3+flBQDU9+2
lVmuSSIjQvzl7E2AQzDj/pKtxJC8yPqfbk1bxnMXGwyuwJ+0lSp7/IV+4K+inclp
NMT/TgolWz2/OLQ9TshPbj4l5IpS+t3pLtg4saWZFhN5TeA881ZcAjJH4VH5sISf
co9J/Ac2VKolQ6BxuWece8ZRUzczKn96ntpEVFjw9YF6jcF78zCkHPqJ83Y9ZNGf
x3LzMHkXJSaMFD+o5MBocP2tIrMHsKdb3DeQwBS5sLGo3xPy3xFCKPIPL5XytBMs
Nl1cZaNqtRZJ3mdaxn0oJxuLmeVkdWSSUikkEEb1E6pSaFnrg+cVyimS7vQMhsES
u5BiFp7b7G+K577PAZdrsKDLqcgiU6dTClU0PnM+P1jTT0HpaPYRne2UipUIarUB
HukV5DeV82H+PoNtauSv92OdFhHYdMR5KH5kxu8O8XKIhus/K8KDexerSYX/dZom
GDQP7vIaRQzDbx6q4UKK0EN5nmMGNRVD2maPVg3oi0CVsiJ30CGveouQCERs3nh2
w3uRbF8MD1d6HMUbxVOfPPgF3X0iwygMhNGLlWaUMULjvlZrqv+gjhoOcKwdj+4G
KGA7se6tzICLMvgN7znuPqPQdCyrz9adZpTBk8mvfJF96RHoinLtgwB7Vdh8Gh5S
SYoBnThZT7HC1NYjGbq8XJRCx2CBGlZ/72dssa60LCX476rb4J9kKZc0Xq4oF5lu
1DhpH7egGwe9tP6Kyhl7rQsO4JT3WhoFJZwtCe2OScFyOlsRo5LdoNAhgqpdLOWS
Zowt6zBm0I6KFP4a95R5a9oP36UMUoR3l2dvAB+xGhoBS/SMfQJFqakIxQwqtaju
mofDaQZ2T05Fv0Ixs336oR5blccD11IDO/M5S0EJ/3FUY6kfAjHWdwlPlO4P8nmR
a/aoTduHPLTflCfnreTUAzV1HbwwIqHK1rKyVIUzKL9RHgEEuAAkZlWmuqb0F8gh
3fUXPy8zgFk+Zxc1qY0iYrbiFYEWiCarAX8Z+C373y6BPatzyS01UBX+xsb/dFMx
wSdFZPJh3zcIn+fohOP8VCWJ2k5hjdKXLmHrH3VIeHcpyxQsMtAjGall68joZeDs
aimx+zf50Pu8Mz8mYPjO03WRGXH4Yv6CmsExd6zQBfDlOuksedRG+RejjAOMcErR
Xxb/5+pGpvmi+tmubFL2uBqJpX4rJtJg/Ra17QfXwQkNM/QVVt/zvVTGTR3bRwuh
I95KA6QgZXbLcduXVg7Td3GYwQuCEeyMhRWFZ5dHEUIcpJQHv2paWoXbpJw3tTxN
IEZoNoLP1gLqhcm6yx6DN3AHa5wPhl2ymR7+2kShCzrK1a1SFjZyrNzFs/smAYgg
OLM6Lqb4QO8vjn6iRGzvXHJ1DHU9MSswdJDJf0H8Bxjvilz+ED+W+yXEed5Ax2ZP
KB1lCJHYlPM2qyDEUz9VCgxjPmztZAB8eNRvLtmbNHc1+oBC0P7rLOf4sc86LDQj
zqt1p9JHDVgV08+QvQk0ZkC4H8kDp8Z2EsKbBC6cLm3ADHNSxhQuHICYeXljBRyj
TubgI7PPgyVzShqdTpxSJFO9Vq/jvZ6MgZx6OIZB1ne+gKhOt4FGfAStyw+09ovY
iRQ0VG+BPHMVRHKYJYn8VKJmlpGklvxWd7Dvp0AYPj0RuSdIIc/nH4IQhTuXL4Kp
T/czIutZHvweqOQpS/mwQqkDwlbJ7gAW1ld4Isexcjo+FpTnNDoP6Ps3rY/sP8AW
a2A6RJ6Iq0UskK1iyH90EyrcnWbukEUdpDqtooxPmoQ9gwQ5e0FEvQFlHYkPQb6C
J0aRnRzYmI8vBqKogVYyreFn2smYxymHMiTrdergFiSdJjOAvkkTP03RV/woZWfo
MvCJquSKuNW/C/TqKILU055teM9rNyEBOvVZCR+evp2e2ZdJR/aDWpnoJOxNPdVW
l6V5Ig7qdAr8/HyfxTbYCx4sC+fG88zUuKUbmFc75/CgQIhlYoRCcFL2AQuGcTBJ
wVayTBJYyM11NpkfaBR6HTW3WA0T8i71XrklYo+sTGIaX0SbVwspw6nwB5Tglpnm
IDQNk/zNsCCBCTWNQVZ/hNOxIMVqYA66XbJkac7XKDFOJEMsJ5Pf+YgKuUP+7KBg
E397Z0yYDJ6P5NYWOW09UYWCrV6bLpVNuOTGOqQKC01qiImnze0ZjnsLcWoPNzel
EuFASgudypzyDuvvkobKzPMWDaWQmjyA9rZnTu7VHvfPAhP1HutJTH1aHKZETMcP
GAD3+jUSrfCG6cnH38MBf2I/DZdMjcPrcdfl15Vdu3HeE7Zvkf75z+wFvjWmMvnM
w9EBZt5jS0+Ji+EvDrOj0ih4ptV4MeJOCYeuxH1LXIyk2cwgaDpHzOD3JpTfw9U2
yOhLbxdEke3EpxwSOXl+2r0b6Rwo44TuIwW7XFBLXeJaNuQZIQT5QQGoYNsVvaYs
0tC9nh4Q9LnqEZFc/3/wPQgnOLHzE/3mgu+rVKGJ3KmTLmouPnHsT5tMJ+TyDSMu
/MR7gi1PmlgfxQNeOWAb2EjGq1q812wmRuRFZLNrH9eCqfivZrE8mfCB8xoKFPaE
fuO1ZvpDtzZ2k7HSRojAZ0Zds+N5TrbLvyTLiiyFrLg5NescSOwTBpNKD0HP9pfj
8XWpbSSl/8gwSPDIgYcAphZ3u3H+1pDgACvTPi5qSZRQq3IsKR5hYSiQQ46Sk+5q
BuF+C+Vs8yA72vwpaUV9I1XFpf69anC4K3PvU0JC6yq2EP4drTNIjChoTzb2Ujoy
FmLg9UUo8vOVdsHTyG9bagp/X9Gn8xLIPJtgqqTbkd7yHip6/L6l464qpuQhxmc0
Uz3ivfHtyCJ7DTmKzcg/ShQOQcUGDSXuk23oFPYlBEFn3Dmrsiw7XJjXxpnVRQSk
`protect END_PROTECTED
