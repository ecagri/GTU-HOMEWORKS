`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3fERBuhi2YbwUAqc/mkJrmarfUkKZunEVPJprqgEdospF3Yr/c0xCDop5/Fh4UOZ
KeI32GLCYxKTCFZT2Nn2thvyS3Oy3FRkdS8di4Zbnez+ezJY3LBunBQTeg6M8439
mV20kvIW9myRaQR9DUo04wJ87ScVMy4DL86+kyhZtirG4xcutRLvFFyeAhSGyRfs
dHo99DnqFeOcZX0NDRcoM5c8ukxzVkitvandHBvZoSTQE5ZcrGdvb0VJkPKQLlu2
M7MWKauamxSUZKiIX7kdrVWlALS7YP18dJUE9bAyRWqikdHVe4iocroXDCHag4DT
HeWTR3ohyf43fRJK+kutG4jWduk9cCIyWLJJXCP6VNgR4MP6Nqf2Q9+9yE1LJIXt
7tcdS0E/JiaJ4xcO/3/AupWp15E5HhipH6m5zql3M/qvIcsdyfahjIOYQxnWzvcV
A7yf+Vqy26JgOHhJ1JiCBOhOGU9qndUKw4nAmrxoE18fq7Unlfouh+DnSnLg1bZu
47pjFA0VJSpXsjTnzWDNp4p18yDCN0B2D4l8zOD6veBLWk9KPyfsaOaVhVMAB3vR
6KQ0BimhXhXuFwqvwhC9AJ+z/ReLRuMBzoxRMz4i8R4iBqLY/DC4g/rlBqUIqjNA
hKMCkZ/a4iwGXnz65XqSllVfcRN3WVbOjI4vu5FaJk0VuXh9WvLCRdPuXW6BzXnJ
cjyYbr+CQuCCJiWC8fBJlgC3OMTJok+3/dyzeOLBFpPkZmHiwqWclC8Giep31Xaj
v8w9HhbX8A8eilXqHsUAhJ+hdCOAMh1MPogO5XfMJIt3lZFWviXUuBipr9HbAkuT
B5xT1BS/mdo9jBIqItARZcrVFvhMkE8ytNjD8svuRuanvyaEgOoImdXNYSXY7+V8
i42TxNoSB+wpvdpBO+xlE4khYkdjpHotvi9KX45R80csowB53ZRpSvqWoIdK3yHv
7+qvm57XjKzVLPaxxhyPvBd2UtFYARH8KmdUIqiAjbH7VB4ytASO4sGjsmII5yWa
MUu/MWU4icfH0UcIMqBbZT55f29/bWbz31vwDs5f7/2xYNpOUqajIIxnCcRL+pXk
ReOB3d9JaeYkiyzFaVPfD9vYGp3ihSafJUmULu6b3yjMBL1AQhEohvuwFvZldo4Y
IdnY5Vrkfq3NpQ8KPva9rMLpyyM3V6K+jfifY5I5PnEfOXR93l9Mez7IZ3USnKat
PPvS90z1ZRFg4pOL0aJSSLyfJu1mX2Wa7FN5g7rMH8HXBv5LQEtlXeLb1nnbC9AX
PmyUedU/aZ7yvqqMtFuwtk+DSlOK4YsFHu39hj/AiQBeHiRE9A5c/noc+TVJBmxc
XmA6CvuV0A4gxHoFdV+eHgQGarp5+89RLwGXkx9T/4c=
`protect END_PROTECTED
