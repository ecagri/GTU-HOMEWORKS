`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z/FwEli9AKv2pO2ghajajuv9av3GqswHQGcfiXXya7NDFcTiMCIFOJSDKlAzz5dx
yZwJMhE2S7tcuSVnZVlETzjDcADcyBWyx62faROeVsPsLxqrIITj4w4i8e0kZytF
9ztkO9jsU63Anrwq78kNo2/cph+7S6gWYQ3QrgBK0nZhq4jlVU45NwDDTMxtJGwb
ng4qpoU/gmvRp18G0glPq4ars0YSvD9GLlwAUh63wfQfh1nlW+Xpe9+tRlT3qQyQ
7RexHsPbDu63/Ly1SNKzC0/9elHjs1Z8tBe93IqUouu33YvgmZORAEQn2Ec1iOgd
W9mfXOYhMY0Nn6EiRjcLL+EUzubbQssk3oMIz6yj7/yptYUwXzkV4YiDKzpiZ/H2
tscVfmbXYIQH/60vbXHKeEy5tt/isQRzpDhtKEn94OZudAvpkloj8OJg55WX8JiG
D0S4l0RzUwWK6K31hlkPpm99AVNhVkYQa1GkOv5LIi7gYK70M5X3jaHaruw6D86A
gQUiie2cCJzHWmIjdxNNbQQmyq3Rr1+xGsA+NLepm3X5wZ83U1h7V5aezK6EMLcQ
gYqLDFUDndKMXCsnSXoRN0aMQdw17oPcxZPPPxzsc6fGLEsDHC1yuXD8/lDjWNHW
DnAnycSge1vYYoshhpP+u9uNdfC1S3hrTOOUOaY+NvvkLFQfoy52MoB0UIP9qrvA
6KFZGq9ozhsszYeRuidezMrMfT4Wsisvp8qnlph738riYfyPTyz+kucz2UUiRXHT
eqNT9XEX5yruCkBrHgFCz0NK7Yqsk9xkeuNU3VT5/eUO8XHVHSawWEp+uFHPfIV9
16rifAC4k2LRWVBiwUmO+AkGIyVjzUFyIoINA3BUuzS+k1POuZLB1YKiv24LX9a/
7Y8xaDJSCKCafbrRI+UBsrt917aOWWhC7BiaeUkhWdywULBTee5hbeaprphy1wWV
O74xBRRj8pmVVSbAzwnqyA5U6ytCa/ZpXun5mPBvnaLGMJrYZwE2h/HlXE5T6wK1
EWkAtxd9aCOAQmQ6rqQazg6rhkcA3ynJ9xqIkoNRh69GlCGl1DOjZCwQERlaE64B
C/laeCHOTdCJ6ZRy9bLiXe7UNfxA84qpNFjaBj5jf9XbL0G7xrHfcmuPSob4mw2F
ZxKX5DUdg5NRfmPpTGXtWWQWSsCVsQIfGQ/c39l0cSDQ37CmY0owQ9L5TrPmhUL9
bgaTRq+DPap4IuKgbRyQjdsRLup3RJ4U1eLzYVL3Ey39YV+TvK7YF4OZ+WaRpNfP
43dG54TEyz9u+a8LSsXm4jKqHryDJjaxlPPj+RJfQJBA+WsSqUctf43Q3L/6QErC
E3ZcWWx4XtFoSgOye/JzucqWwNSslVOy6u8pOhz+isQyBXqGidDjy4W9DnmrzABV
rmyl2RWBs+zU5bvPCMlmehef44DzVSGZOOz7RBm+FBKCMsOrmCVYrv96/qA48I0x
zNg3dH91i2CJKcytSB8nF6i1lH5d3DWdTFdq/oKA8n+V9Z22syvH5mwhIcbV3jYD
xqTl19c380c7F160c1nTYaXjs+pWbeGjsAgQ3lk1sy5kHxILANzHjOK9n8KjeRMH
fl3nG/+CFgPTOG+iMoQnMEYhnB5e0hwYUCkjuCaBGl/MjNwiwvseBDwmk6erj0aJ
BcPua7UIvL+DqAaRvdje/hDpfR1vKY/cg+xDCim1jFCfPtqSoVEF89RLunTSbXdR
E6D0N9pH1iN/NtQ6TPSRassFiJN5wNYhSS8f0IUCXQ584lo/aAd8IVo6xLaRdsT/
jeFeB6g0/eMHNUKDPWY3XXKUnrdePGHfJBZCVOzkneSwS13CG3LjsHDyJf0GwFTs
JeLPJ6l67x5oi3YraQpXWqkLLvfo31NPRjUJZ4OR6ZubTFxyqtZauzZuT51HZNwp
zXc//yZg9hrYtu3o1Kf0cKfo4vP9ND7qxkHM7sYEsdAdhBK6yLgkD4ob/Jx3qjaG
UXfY28MUsgO5d8cZD9RNQAGsQX3xbUmw/FRgDFRwdZOgRWat5A+vpohrqozFPyd7
2qdCiCJcGwjlNrK0/N7XK7lmJMqiheAu0TkHvbQZsnOt4RvmYqaOMlEQQJ8OheuS
ixECmf6jJWddZSjDnEVz0NwNXksZGZn2RGNx6m6SPbICZw7J9U5zG5VYisU6gOvP
8kEfD0fXKKpLQpqztNWcxuh43bxB4SWBNFWJ0htA2vruYkKz30QvT66U9/1d+sHq
hmmN+dyZHoZHmlZXk3/j5z04L9ce92LP3qlTQjk6yJKLzgw4Kq0sgBodkbsGeNgi
bXkn6byW/B3cBjHWAdvAY/E4noK4HJBwsWIkRxIBXJ6UUbUX80ORYfpYh7mwmwF7
+tFPoJA8sZ8DwNYoiwZ59/Cy8Ee31Zw2mLGy1gIpNCAPJRy4RGftIwzPYFQ6YabP
M1F14+jtf5EiZZlFC/gexStlT2SUf5svfD3t2w5GKvJGg7wyNxSQmVbaVztTBdbf
QuEuLJDi26dlaaU7X/NP03kyBtVxlI6fMHVRBtlWcr2qW4D+vERHklKEEkWYU/GU
gw1EcKWcmh2wV3BkPmIa5a4AXvPywjIGIMRt7lKfX3mmdFQPEeB3pMbRkWxRwiyh
nKeIB/Bd0Pm8yLykn3c0ilsyux8IcC+/NxC0XlLNtmqL7XJnv4uKGdn+DbJALfjh
hoQ5phaVVyzPZDu4GTgPA17ipEgQcaJB7B5MT1HjfN2d86Y+FjECgjNqP96ugfob
+NM9tlw1OmGRTw7vYgPoSiHiXJyaf069/nU3IPJoWyxF1yBqtdIU4Fyu6gQ9oCYX
3jsNyGc+7duoBFVP8LW9/LaCq5VVf03V3tqNxQmFTufrMOEzoRswcb76Zqp/pusf
ifUonIWnoUceD09QGNqUTyYVUxbgl9SLuuirP9b7YlIxQC4No4NmV39WWwybPjiQ
cXh2LVXP4bgPo+87vym5Ars4m4BcTBWPN7CXbAV4DA9TPMt3k66HQTYeqJa0u5ii
5kl48/Ny7syBjqOf5ti1en+rjo7pk+QZZODAbOYwUf9Y4kcLOdpenYWZro6Y7LQ9
e/7aIHBjMGIebSyD1r5mRzyL2/+Aom7aPzBWIaJJCjvyAmEZsXRtMsY8KSE+t1Ec
7N8v+WMFVLoi3nu53mm7npqNNbwf5Ak2+dZcoqeAj12rkjt5vUlB+yCvlEslBlpX
Y8TxGohCzuzbzB0ZT/bnEiwH1BDefV35c5YPzRkc2bVslR9S3S48TZ9Nwwf/qiei
H6wZp4c/IuYvSUZyO4OJsEBRACf9I8tEOl4hBeaHySK4n5T2PHL+rP0goWYg8x9k
zsqgpLil56T9QKbTZWwk5Iro5KVKWz4ZP6o7lq4anBh2L0ksBT9qk9gAv45cNFfP
Ibp4ZLrkbFPkxNM72b3zWqgt74DoMNpqJFeWpTgBfY8eHqTsPQRbb8jo5C432BbH
txPyTiT3qcza9u6n34TFq49qrSfXX0eWq99vKH8APFTgVeqaTWDnp6SFWpbsEOk5
jrKYAWbfcCvNNw/fjmIsQMPwAraH9jHLzZCsJ5Jyf89NP2bdi/VkcLRXux/0KLoG
r4N/B4URdLJYT1avdqteF/KaZ4M00E01pbN6J7uWsLX30uARKSaprw1ivIdTIKiS
zpf8TeeTAdjAhx+fi+JQEZyQ2R1RsKHj1peX6ft/u2XmTadR3XG1VBzBE8gatqlE
XWwZ3AVG/HT5azoLMHSYSshAS6CxjS6fv6LOYG65ubM0NdilHFhLg6Lo9wFcYo45
iKv9ld/h2XwYsRsOf2w8rRpQZV2KehSWtae90rEyfSYJtMYMcE0d25ydOyllX1wJ
rCFoPxtE8jRBlehLZwx/xjEGPGpofRWm8o10v3lDvWXligWQRijZc7mWzJX8fyd7
1BH9MeWuDGx1Sa2gNceI3B1BpiJzszl6KHM9nGkqjhYy+9Ctbp3Z+DC3AsINUMBW
VGTXXxgIegmdCZ4e6epvl9rYuF4tXjXhp7bOnghEW5Nujpvf2UhgSae8qmXcG8ng
uzLLSLSafNAVXXavzvV5hWmcNY6NLiV2YYp02zIayXvcuX6ewDhcdTOpNHB6wIlp
DLGzKY9Pp0EXDxSXCFbBjhJ+hmkPLnCv4gQSIL3grIY2hJpMz5ybptavhyXfB8VW
QP5fYS7aHQms1T5MVgn8NTtfPRM4M/T6vc7NWr3TCxUWqsjDoXmL/2Q0KPoBQWqM
pKx7Nwbx6YeOYCD4qEsn7P6QtnXgMqQW1OIfYynijJ8wwhNKIjNU+gucRAfNlTMc
PMRHQPNPWL8wPJWjlUnJN1VdfY2L6X7DVD1fJkW+EbpYyIbf0u1pFw8gWJRthvIp
qCRjxnE+c2dmrr3yjRCQMowz6lCPoaLIEsckYZJBuUWv6ISln7QukUEC7viH4bgA
LipfY42icjlFxz2MGuAAH1iJ78bF7q2o6QhRnEs33lSJ9NK1Mp+0uruw29UAE3Ys
H3cxLDVEB7KhVtX6z/owrvbTEHSGUdZ7uwjKLzgaHBHrt5KArlmhpvDtjnYX4x2g
V05Sf5zQmvPtM48HlgFFyzzj+Y/md8E9D2p4EzEKY4VNOwpsCSKZMAgxyeH+oGJC
/wviO5OnH4WrlVAg6jsJbADHJCFf6mYDqg/ZwhvxLl/EGcvbhLkYE1o9Xb64BTtD
LeRe70X/+3lsak94KluVCNXPfQgGenlVc3JDJI+ZYuTK5wAHFrCaAT5A9Og5f3Lo
MVG1Lg4ss8DNPdDGNGhS7q1S0CilvhZF7aYYnpr+9o6nSy80ZAbVF0BZc9uhdcTW
X1ypud7/ufbVWGpJzfG5iSM8lFwYqNAV/yDg4QwDnblxCoyNSY/Tl/9Tg1EpwpP+
RMZXHWYnrvIUI0PPyzBZV3rgxqK9NopGVkSUEIL9WnnvXuAxVdpCTyLDQJtZV1Yu
OCEERliB635PE8PmT8cnZmC+H+cfE8yfuv2REp90SCS8MeANLeSqs006STImZEaS
7Opq1A0SMuxTc1mdhM3OAUqrposn4GvAYPBRmUGTOuSSIk8aPaszbTEDnNCf69W6
5LyZdQzgDkJbwAhVrKI7JRMfuje9L1nl1vkqZTOcjkDlGkMD2eODu0T/9qw8O/d1
E+hhLjhma+HxxGD7SioWqaTSwvYIb/z7GIQfsSQtAFrB5qkTApSW+8tRC60zZW86
eYeeHjq8CixVhPJ738Xq81a3klerMH5qKQeCYguAiKnxaEznrVHvoyBWFxdVN7wA
JpW0/lE5mhpIZjzfIxm2YVJ2bH4NGgaNwtpRdbX1z0uTYOdSOMJPXaXPIWd3pnZp
lscqATNTEhU5fx5x8QqsanFp6ELM1aG+d5gUCJE/sj6628NxBrnElr5r5W1qAu/v
khTLHMjHVA6TWThzZgWwRCioWeg/sbjGtYKiQbsAn9rQwQuXitVJAQFlJ7Awk8Cb
qVh4VcTGI4V2EXxfh9MmqvFvkmThhoX+ZvG3nJM/wHeVTKQqMhCDdX7DHqPO9FFb
J+i6cK1aBvmmXLlxvc9/DHWDzrLxpiFyBGqyl07UMGQ8k5usbUbdZnOQrrPa/epY
DxF9XBBIZcSZAickOJdeYv42VeUAFSBDyGgl2IdbAvCiSu89SfMFX30XL7KRNmaV
2ubs2LpUfDcglMHN0BIdC016UNv0CUPvcKmVasgOZDbf4mM44EGuCNxEvDmFHju0
SeFUNcSS6F9hklt8dqUQxznXMt/8tS34Go8GmiC17JpTCCMMuzWOIlrMXGLUsG0O
5niWF1a4ueeJ+5YUtOboXayx790p7bnyxM/uMCb+phzmee+q7IpF+nmqBni1mIqN
EfDg1M74HfEnunY/Gpcs07l9qMibi/l/hKvAzvI9/SYnDX4w09zr9IGJ1yoxVTKO
iyY/xPQeP7W3dEsoNb45UHSP+iCaxX5LGzsj5Dp/drxlGwj5YCrBO/7aONUlvVQi
KQQn8Bh++kg+WMWLWvlBWfginTm38tNlbLs3sIzM+d9MhIsNT8JbCgxd+LqxW2zI
MPpIR993ZBEUdPtUFTJSnPLq7aWRKpED6szzQIGoac/2UN2yzMloqxiNBXAjr/Rn
N8uiQGAXXvIOETHbtPxIhYOYaKwStTszgBfpsPjlqzmreqDyNzUHDuWCGhFq+y2P
YAGsgpCnX3D0hCT1rcOknffVfdaU+1pCh4GPCIeEjmelOSXfBdZj6DLpjr7LlTc7
tQf94RxPn0HiJ+Dv5X0QPj+XXqZjNm1EbzB8PxguJ8ekfaTfXfMSbUSmuca1GgnN
hBnh7q082FISRO6FQpFBmCZJMw95OqPyvdBSZqfoxXkLnvdGDBVb9bHFarkL/xAF
fnN8ssQ4l/YuD6Gs3znZR0Nb7hM0dqb9SzivDGcYIAgwr9GZ400iTQ0AsLpt/un2
GmDwy/kDkq3qK2nrGDJHq/5svU1yUBXUPCYBYO0JPGMiGMENpgbd9MgNtw24qpHH
m4PDVJ0jt6NCyCqwehxDgY7aFCu9T6CtMBkSIkGYGCFmlFhz8TcCVqO2wZEpRmlS
bJamdnYCiW90U7RJQGG3e5/fcYEAYl9xlApfUulc27OqDstOwb7NZYgnHZP92X2S
KmbmNqwlVq5mwvmpWTF2hEhdgoytHqYZsPm54WZt2Nd9SOUh3kyntehnNJmWxNNN
RWW+nmszNKeh9LWPjSzHq5+smwYsY+S+MeiEAwQ3Kr9XEYixhmRFHLNyiDNk6HbV
0paAscXp1Ef4aQI2OiKzLw==
`protect END_PROTECTED
