`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3T8X0scv4nq1FMUOsYsTkzYFe6d6XOJ9B2rmh3Wq/NBjvGnrNa2XPmvuTdJjizcc
Gi7P1dy+p25PnRPUfzgycanzbd2U2kRgm2OaSqur8Q65Z+bH55qlbcw/8aGu5FDn
HBg7Jn53cPIWQyUVWJ6XWy8ZXZInHOuLZSOYeKemT12xLHZaUoL7MIle5AcmH2QU
HOOk8zqJAqpg28hIJHXVd60lZTuQs8G6Nq3vFkUV1PwSiwoePOg1LMZMTKoPbH57
f9+40RNiGmX4q6Zx8jpHR4OlTfa4qalaqH2Kl3Fnnuy7FAMtWwvl5VQC+R9cM0j7
Vn++TGBRmdgRylL/237LK1Zti+IsglowS+cWcDnNeK2OoEYWhZ0bXCLXLR3X7Y6m
lZB/D0IehpoVXBRTv49AIS+mc0R4RcQ3PS73bwAVjvc=
`protect END_PROTECTED
