`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MkD2d9F8InozOJt6cimsUmuwvXHAu91byc1MJxET4a4qvd5/GubRi0bpxMFxZVqT
/4J+NnobjmBoT9So9EWSGlWlDxc/07IhSHTUcSdm0urLLOCW+12PcTYEmH+TR/x4
5ncz/bh2OIdWgoECEMPBOkMwoXhsQbHvCHg4nYkumKKsVorvK7om5XEO/gawGUIP
TejrkzwOaaP6sFhWnoxmhdzFILrStavW3jZyw/bcXxUyBttYUjdfOlb7k1INuZgR
+PnTU1m2VFpX0WId5YzQBQSkwszd3AfPxiZzz5XJ1RGETmX8JtTwJAltRrIS9v0W
Y6CBAPkAo3AskF89tHfVDMXgeQtIMFLLYyPuNmiLH5Sng2N0lG2i0XVzcIlXYn3y
J0BQ4XoeUzGMhKol65Mf9MVUzRSjuDwzo7pnlTIQJu4YGerjKUpnBKlfG6JWiHxo
b1Wmc7BGsLz5x5QCjgeqym7/lFISf8UWsXfQGLxRRAG2MXwAcK4QRAPkdMcvYGXO
V5xrGpqgzEHUDGnmRtYahzriWZV8goHuD5u2QS9s9SteDQi74f9hSCS4TRfSErMo
hDKIcg1WIMfVIWEznSxAxZmzEZpSwK6FfRB0mq9+ziQ6z7RL98/EwioNGct4poyu
ghPAws2bDMI7jR6CQUSaPaepPVLfOXq8vrDkQNaSq648O3skwKzDcarViBnCNew1
4AYJ12vWQ1COx+oYjt96keZnZ6VEb8b6DJVfBmdMVB521RdT1bldR958LdA/Tjyg
Q7vcjz0XEjfE9+3G6spew8tEw9nztZXworcTUaWbdHTr0CaIq+PlnbmfMwoo3QxP
CkkpqVqFBRjXBiNUv7vq+89V23IFJfHHHroUy3uVoz0dbRZTIVKYbO2ajjzHtDVS
UMH6A6A5ife8EGgHEKAQdXY8/PVVA74SJ2kemarlZSgIIX+nbLOMv1RHB3iNk8sh
WKlpVRDcgEwZNOBL0QJyMo5Z5lA0251U+RJ8lo/dRKHCbL27+5um9HtHuSEEfaoM
/pilGoHsWQ/oAsyiV5n8GbNm5Aj6Dd8BEPxVEeI2b6r8QERoPTmBomJV6Cf82ZRH
ovcQ3wBBkLQht/h0o14iPHU0M0Scpgg3DXKRSmHPIsLPuJPm4QQa0mRv62mmYjky
2iNIrsUeBTkd7bH2bJz7d8FZerDpq3Ar7eRkGg+tJQ4AKcn2ec6NJ8r9SSQqKyr/
McHH1pf4iuI9agCJl4P6XF2DpNBdOWTpyqV7G6GG05C+FuwNzpOaNH375B0PyTr+
OP3C5mslI6Kvc7ikJLFo/r7YQOpKdvq6WUm0DnY1Nw6UX+eUPgdb3TKT0XCutBig
3tNFLQrBBI4vQcKOmTe8I9FbXDSu7x2rn1LPL2Yu1GAr2wRH2B1/TgMKOU1SFLW1
TlJLhjCwVqiAHm2yWUWQVq1SeDUTCdSFiNj/mBphnPMeoTC3wuc2UgcC+78MQIJy
PcIoutZGHCFJHLT6mHfuR6qtzxdJHQ4G1Abcm2wEXpWwQGA3lP04WtrU8M1Cp3M5
WfhkHvKI9XemxKVznoWfe8H9jTAV+ZzVaOLthhn1VI/GKNMvyGSbpnOIiUQZzmCx
`protect END_PROTECTED
