`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2cHEpGgfovJBEAJAbUKx8QyOTm0kaE4BRgZDtgKwSoMGICyP1518U1TrO6SKea2O
jKkPFhlb3EQaWm6SxKS/z6A11UpCh/hqYhzBIV+x8erTqQ/GoCfQLvVWLN5l7UjK
t7xwL6ih3g8umcs5wHkbMB1KgA0O6eQ3QNAzJygWjsHBH7JMk4AJbVd31O9jFgAO
KPAoIWPAPyWCmmZXE76eDslrJwezhXShnQAh5r+ULOLd5252U6PzFkpuhwHBHDQR
Ll3YSs0B5RSszVNm6v7W7dmX4ZdYFsKIAoPEnqmIcSS5AacSEhr8TugBe7i42w3H
ZUP/QudK7ZhuO7ZcWVF3znoUOMPjUlBCJ70+ubYHNMn8n3RK37l9CZtSt+cdBZJ+
0WoVZgBT2aZ49AUyllqPsdNsMHVds2n33o6jafJAwkuVWCNuaZ/XTlrzJHXNUNNQ
CLdbXpAos7encsJxKZmPhJsyNppJ+gZ1xoEaZP7Jf1zXOHWO+1Qcir+U7v585+fH
p3OcxcLRvPQod1vu/NunGFCodWVCcAJZ1+WHbY+jt8mRcOhYwWzbuzWJUGXfxQfn
G8Ovhx5E/XwWnrmIZRC5N7nQ4VQjNILZm7RWFV8og9MN1pyI62jtcMTfx2whfuuk
buZJBaHI0NEKDQILrowqwayVEjeKdcg6RZNmWKDYs5zlDNJiWeEoax6rkJH+E1H0
i61eQb53s9TNGz8tWmjUJXTImD+hBhh5j8iD9WYWwVqVObuXhfmJYIUNkl9dn5Ml
pAQjKlwzveuQ4X16cRqNw0KvQpz5xvWgJnbIEH3gMoXBruoWLYgCBSN0vLlReYwO
w9jghiMPPJ89++UMl1qPJJhgdRttZRXF4VVsjthIKzAxqvPnKyJKZ7daLl6o42hT
4KqDAOYVTOajQNRHdXhCE9UQemAHa/Xt0Efp5u+MOJPnWQu0mWaORxBU7TJ7jOUP
LpDKBS3daEPiRkM6VEUJwtW0NHKs38NXnYc72EaQYovgkUcj8TMeu9r4CWFZ/XFd
Y1KNMw9nZxENZGj8gRlCozWBku0qZvrhKMgg3bRDcqEgYNGmYnoO4cB2rrI8FxJN
dMXWakyETC5j7l7acmSHbkF2yIdrwfvNy3JS0kWmffp++b1lDUGSP1fkDtNfXb5s
3F3JYj5ynjyZ6kV7nHEk+WbyP87cyBqHjWDLgDU3uQOJfzdMI5/wdBXY7wL0CVbU
oDRZLXFtfJORpQ6pgRWceInKvAsbH8tF2pS2RPmgK0hI1csynDVGRr2qmnEG2sCY
BPg1VmLgTDg4Z7mpV02L8xgbffx3nmFWHA2w1iy3pEp2pcHBkOdODNp4xvM3Wjjy
o4K559HaVvXLXtXe2ar3tiuYE/t4ZIDLzBgP/M8K3lYGv6tb18ptRold0mdxyLjd
7MqDK5PzbM7n6IfVcAONGlD0lVCOxkDgD0RZQxMwy1ozT0ztVwbJN3GXP2L7FDBc
ZykUjneYXPtDRXeYTkUmXwx7r4qEhgewELysgYddZs5npffYydPuZTKNWbLGif0L
1rO5vGT8KssB42XqQrW5BRtlecHdvSJgI9uaBTILsXFtNkWBLUFJBB+waKqB4QA3
J75PbxhYFpDdGBoaICTkM/yFBoiY2Wx6GANAh65AXeZWYrVH8VtFWMTj6Hk46tSC
kz1JfcgA8pkZG/zmfGDemuZRLZCBBSKHo63vqx+KBfx/zXamOBkbc8jXbO38BF9g
+DxhfLFGFFQhLoBefepb/7zcbOJ/9POCTV6K5AXS/iLNx6ruxFaHg2qHijQHDQVQ
l9JTnT2IXZDdRO7MAOygd0oJr9hcs7kQhNW9/xPzKGMT+ZvnqH6qzJS+JYlxU2so
FVVAENIKgrN+4Rc+mftSBwRblAgS9MnSanxjOSqh+BDPXfUn6SDsvX32DoixPeJu
uOMIpPD7DEFYBAiIsH59LilwLQol9GzHW2UsCOfnOanDLI4V/+xn7BQDivjnSaF1
hfTWI7CSN5N33v2TTziymI1M09e0Zp+bJ66iu/93uXu8GnBcRsA9VqfOI034Z5aA
eFUQ44BO5rglL570QpxBXGk3u1I8+KhThiZosLvdVQzK+K7aSB/wTncJHiXs/KFW
HcFbdDj+a39qPgsf+JP9vevhlHFp5wagnf0cAWO+o1KE7h/PXhYhdj496IDylMmq
bpBuLFp26UKJtX32jv2U/ak/uKN6lRak8j7pfNKe/V7bdCDd6ZQiHfX3LM3uEJ9s
9sj3+kfhmKaYlk+57MXe/MIEUz9zhXvao7LEB+aJNwHZs3UDxvjQKXufY+hzGaJQ
DyUOcFFwxFenWeOfFxxOdD7qMDXQvrf+xVOTQcEtH4PiZFaj+UVJvAiUsYHERiDr
W8JqM8/uGaaLSGm6m7BSOMJ89XLbVfmD9/u/ADAS/hWKGKbdbm87Uj4fndstHDHi
5wI+BgmytzB4n0PGCd4yzU3Z4cbwOhESK6Ij/OhESXUOHam1SJW+cvh9mOxXAbYB
5tt36SK++xX2BMS2aoUvswhiCFiebBb4GnLMolmsmnoGrhykp5m9XqdaWQ8MQ6I/
AwTcCOqkgkaefe/XpemNvDiqiV50b9htw2DJjzpGlx0mShSnTHYRBjMDaNuNGDsr
zl3l0Lz95y3qoPQEXCc56MevVScsWUrUrIWW4ZUvoO1DfqPC0IPFyjMXnOhhyc4a
jqWFb3kyzjsd06NNeqgGATrmHboUWWAt06726uyCHTDCv+Itx+1JuusUYULU6hDK
+4VNgtQXga+v5gNQNKwxYVLTcmUA96hqe5f3N/qkdZYq1r9mKbStFMMcKrjU6W1h
cz2h0iM4/sWnNiJ5o6t1CdpjMCfHge2bfxxRJJYXHEUkgsdDfutKjStAh2a/AZYD
Sh4fnOhQOw1NTerWywePFINOhUd4mhWU7T2aZIC1jjOa06BsjQnrIcJvsOJORej8
GE7k9D6zE/YCaWDtUFqs+n9+gAiU3PX3cVmsYyDOG5eJdPo2kOzXbuWwYwUwac4p
mSUPXdmg7trnFvMYp4E5fBOfShzXUefHc6hZg5AsXIccfvUoapmzGOA6HnPKpi3X
pL0BM5JY6ejZ4ZGpc/yRcYS2fQ2fl9kRzeel5bJDdy+u5vhJsLWOczOQ7yKAtJfZ
+fsQTOqG5wM2OoE6LcZdT8TK+W7cvT9bzm4mPFqtLExfcY54vlucK4B0DMewv3DB
JZImtQlubL1k/LL6jWeqMrLGpvYokdcugMZ03nO4p/l7/YEiXukQZ/cLu2uoZCII
1wgegmTMIZV8AJUd7POiHXxzu6cgkdU97aXm/HhTldUFFoouWH9gwt1n7iaThXNN
AxvF8nnkkMxWG62qVMk6sDST936UC99UpHQ2MnCfi+MCS75xPXj4qvjqw3D3iIy+
2vEpsrsyuerpYieF+FAOZBteu8F1C5UjtgJE7hxNRLWQrm9pUC4BErYE1q+Y1INi
nHs5Vc9ly/zHqMYpJcFN1SfxjuvX44ne4POcrVO/goNi1GarNpiWW9podlN1N0vd
hjytqObytdSL8iL5OX2LcsOJuVQ83J4fUdkoDqcgfw5xSHYjSEIZFjMBrLbCa8K4
PsaJfkKYxjBzV3j2C+Fif2bTtoGUP1WtwXRXKRqk5Hpq8tZcWKyizpaaPM3XRKVh
2zZnjm6WNcIgodP7voGyrvEOv5qc/Qaj1sidEVdjrud0kKq9fpRCiqy+6en4n7SZ
jd2C0zWYgrIKdKgHQU7PFAAyKyflt6yrB7n3Skd6qcUWM+DMaJkKIPx48dvWEfeZ
p0C5icjqWxzZi0asZs1a77A50gJLLEWXXwTRANEVx+TVuKsaz6rThS1bHXMjMbkE
+FrfNM4nyQXTRzJ79yRRUGrDenH/exgNPw0DWEkf5BVczZHLbp5vDbtZ+r/LuV7a
2tW6x/dvn3qXrjfTAQVV+2iTQ3CFevhXPtiRoqT+SCQ/alpYD0ZMPoz+qWPoa1Co
yPKrSsysX43j6TlcQc2f0Z6p4d/shnaYD0Rwe2QhIm5cjNzThIbgwNERvN1WClYC
SPo2r17PuLxsPWV3gD49cudTTKMQMoSz543fveHiMf64dawiYoJ8otEETZEcl50y
0KRkjjTaN1AGKq0lcT5iGgKlWgd3rTkqlSiM8Slb8vuWIW+4OK8Roa1DS8nf3dIy
MnAB/n+6g0YqGE/p3ePE84vxiuwl9oHj5Lsr1lb1M/wZxNA6KGDGnDsJGuC19hfb
N+BeMtIMmORJAQtglAEbkHHnJM7D7V+KMiket1V5JC0ZFKT3kSgnar+FbSRbgN2r
uOmOx+VGABWwQzkT+rtIVtzVN31hc/GX5enyc6wEU+IIXffii8sduvda9ibXNFaG
Eeh9vuAJZcavLIun1qEJIErGu2Kx3A3R0S0YXjBE87WWKOEvxza0Ej2JRY3/Aqb/
SJAH44631v43eCzTvfYip4ZOEEIh+5uOzYgyHUeJLdzI7qUknLxD92kdMH09X6zI
OE/9U6/AoHVFXlBvRhCNffZvbIll07jKLk7WMt+zV2iRo7uB42zeblYd1uKdYDEU
WyvDVDkbl0SJQs/hG2B4TiGRk6zPxliAX/d9ZgTrq1QKSWwCKAJ6pg26/XP4nXtm
Kx4SCgiIciU9j1MSUaZ5s6mhrbhNHoO20+zM0HNrhqILWVQ/vTiv8+xyK2UGpX2F
1QC1esT13xeXFj5HzVFkpQIsUsnfjQWyDwHWBRlf2sgvgwitMR2Cm+Lr8ZI6Ryi7
GFai03wNBTXzvsLY2ORjLXcWuN76oUtYbDED2fSgGZlIRHwdI5b3kk4JZal+QeI+
TcNXzE0LgOQiqrwPadTOfdWvICPFBOAFN2Nlv/5NAbykDXRklab1TgnG+wBQjvF6
AhiakR1kkls7eWMw9blbvdNLSWTUHttIufdIT4K9YOikzqi521B7mTgH7g395SxW
J5kSFsTYcVxCvsCx48r96aS/koiLT+0tG66IgjX/QkRzDWzeZ4In2SSeJFlRuhcC
lg66bWfP9EBewh4w5axFqTxcqgcQoQXTdD9UgUXp3uW02Bn/QTTji/FUz19Mf24B
iR9aKw7lIQ7KaE3XrZ5oJWxKv+MZ0Ce6y1Khto8pBhd48XcKtSZnZ1RcPiVZ8cay
x2Ny6Rgq7pbCCMJxQRYhs4M4hS5333VO7QVPdhpQk0VEeZ2RfCN/wQYRXIx26rLJ
P8HjvGRMsX3lGeuFQHpvyj6IuwKhUyAP/hWnVxbZVzMg2niNTUhA3WeSkiGUqMRp
kSFPtM4VP+y8orVHlpgmtzqA95UpK4ywQFK5oB1Lh3fNkVKRI8sExm9bcz8HJobA
B3tGctqLrRUwNRTNJcZ2LwpNrYJ0ehuCownRovHZllibcpF6hNcfpIL5B1XzZE21
n6m2crU3Z1Co1EOyQ5Yo3cspOCrNqad1jht1wpq3DanglhqRuN7Km9NbKL7n/S3Q
1txYYVP52zV6UpSG+vl94LtazoZefRqs1yqJS5s3ClTRTeU8ty4eWKHTBkYmUEeQ
e/w8H42awhTD/E47DuI4JjQfR//Uby+j08zLwYi1H9brWaybYi/zs5EYYmHzUN/t
NtZTwA3jWoONByphkW6OmY/jhAKcoGW5g8lFTSUiLEe+4ICschIf0m4Z1gDI3bZU
jrgGA9WqvQdu17KwjU0v78e+Qx322QJwtR74Oqlsek9aih2s6X9KorAe2ZlFhQ34
g1FyEUHD8nFdQGXDJt1NVqwpcPPmtejr9/nomNJ8qhkhSsPdUKmdNYZay+jGPR9W
0MbdiKFzT+QfSJH4Ewa79TqKPqfISETzgeDDqgtrPv93rrZWlZ9Dv3z73oYBfT2D
yjGkRGUynYjpmTg9CDeQqMgSV5blxLxrtnE7wM9NKWwrQOXo2o+aYrfNQsvRUcOv
uzVQWEti7de14L+6OgkDIuolurldpJ2RI4vwLjXm9y2LZe3w8qEMnUr3PrU4jCif
BwMy3/nW2/bqMi4vuaMXbMlRjFQqGa/76imVbZNI6T+Zc7vTT/ucUvJM7/5fb/34
yaSxHVb7YjI+DbFBEGiBDDztTu0VWiiKjg1LXILTxYXGYh72no4vl07PV+YWTAWl
LKZgiiyhZmgPgZfEfRWklxoU6CcSqjurcqRI+tQQ3je+JKGCT6ASm+Pi0o/tLeE3
GHfgvyTrqYANYovVzm3XKlqCXh9g04uDPbmNfcbXHI8J8FuzHRJqwK+g/btdq65h
z7I6qREjb3TQ/Tp4eAh6D1oCLkMSq+xvSVRwqUaRfLwC69X9V2I9ZH8hOz+Jgrzk
CgaNmyBmzWE9Ll7Hp/oVlwVO8R3XLyzmqMI49Ory32g6+VwHKkF7PMUlqoLirDDu
kUoDqsxu6Gj1i0/n4goZB8m/zMIM9C8k/9CnK74u/0si22OFTPCh8gGgcFMui8T8
U1ZKrV/0Kg9IzcZvTcFRQLYjA5U7I0J/Xav53EWvJ/QbFfmFtLRgsG8QiqLvjg6i
JVexzCfDx2sa2GNCOTjUtZ225Uri0GppFGUy7Rwf6oFiIIo/VPG7GNPS92QwfMrT
UnZGDPYcAHu7gFzXV7C4TG+F45NMmHSsk6h0sSbBRtsEYQXCKuw5Ed5HxNKJqH5+
3cGGMYXFWx+Nm7OLB1x4H5qr5S156TUoEst8h0WqEe6UhTAc38ce/zPZT80py57w
SNPwuiHyGEEDG7pmg+DV2dwcjabPomOsE42j0bOwANLKziyOtbtrj2CwJK54i0fl
Rc7xCzELb/v4v0MIsiq/eDKszSGG/gnlA8khwwuSfQR0nEur3LpgYRQ+jUh6vA89
BCqQjMau+G5I4LKprFwdM2QnktPHr0ZKVOIRFWyyUm3X6c+ynbBq1rEtgwdAvynW
`protect END_PROTECTED
