`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vwjnl+aW4+9/FC55ZcNoOFifpl+zZfd5/n+21aGu0F7POMqj518itdna27ZabViE
i5hvIygoGabQAYDw8bY7W8no12MsTW3YoqLE6mOY7w0XX7Hb+04k24tjDhp0cDxp
OE/j5rrP9FbyAFHue7C/D7PeikAzx5JOOQe09n2SWUkXfeJQ2vp95cymGrHpVRWk
GfqTz7nsXDMd3NYOj30zbu8HdVYrZk6SDsfvdTFHp6oLk5VFMsiHRvZOPDhbOTqk
dKH9hMGZA48tN6Kd8LW2k3zGzH1TtH27U1Nb5E0y29C5Ccvc6zU5hQP0kZwTYUIw
fdLp0Qsu0JorPGycBY+ca+oxEkQ7rskJrKyBLNgoEdepx4z5FQsZDUEiG0m4GOCr
VIT+DQdWbJJIqzDJ3ZtFYKpa0ehu75STj+7L0jqeBjVythuc0B793HjrW3Y08HSh
ca0BCk3LNzaPOTVA/K6/DQc1FMUq7O8z4eFgrEftBJB2/rhWVm/fUm2S63kASm99
UlB3xwk+fEfCKjEYdU4Yo7hkrSNo5qBBI4wMz2bn3gyMyXVLNVoHO0YNaiLdl2Rq
46isJUd4e/erp5MM780E+DUPLS8NNpMYO3kCuSUv5BgEIV3nZH65WrkJCGi0izMf
/5/6h7hV+Yq5mESCqmPApoNFzzb3MuqFe3msKMZxTvD69lBLK00C+v4a5PF8Ik8K
8llgueJqrQSmlkkss3hXAPLHH8cIfmv2PYFrXu8wHdn/G6HHI7rGUnqqRwydbutB
hWZYAhYykOwWhifnL7YwAsJOFh/i0pognws24KUu3OIeT7EiMzv4Clb8yVF9jNof
9t/cHlItx1b4AM0RTldPpUuyaJdjNJrl98M8Vjb8ICmKA8bgvLXWHDRIzJqwovfg
G3/QXAuEtkgAY+s2IBejR0MANL7z3kLfw/70tWxj5lSJGfIodbSxVv97jfTiAtrY
+OvI688LJbC/pW/xPTvmfrRz3mDTyLiYWe/dCzvOEK/qCCEZ5qEo9PRIpHsxo4pc
oQhZm+BsiAQ5vvvFlMGk2Ya838GWMIrh0MnUUloWGm+25ozK6QSx/9LeK5Gv9g6h
fq0tEc6zsui8cGrEif8WDqIujegh+D+F0NuNFj64N9n+RAQfqJ3K9EUsR8TqLTwI
c5W1UkkGsA8FKhrgB39j0NvXLpjyjaq070Cj9U/TlVMppNtSx4UD5FovjCrtcgZC
mgB/BHCk/gXjdCvpm1LM8ZQnUnyXK8fpwo12ryPyqxRUeef+tOO+2FtID2e2NRYs
lfp/YxG0QEWXRhvHgWgkwfh0yXlwhNCA11LRKGBpo/nHYoHcA/L/5a1Uo4BC/QSu
awTXwGlKPruR/FNEuh+4U/yxuyPOUDKTkvW7o9WT4ZUBGwxTVCcX57Q0B+icwqM5
GNNdy74qnwhRuSEyeZuJM8J+bRTzYLfdX25q0ws/XqFN5mj370oO4hx5qgrekwwg
+oz0VN3IrcnEqp8dS1HQzWdWVaKiVjOqtHp9oST8MvFff9RwWLbYno7eYXU1BiM+
0NE1C+sE+CWq3pxql9r/67I76eYFiPaXUvxLwZ1E5ib+JCMAWJLyJBAEAP6qWIJT
ZQrMI0ETPpl25bEJKvuD1P07umZytUtS0UGqKiB/vQP9diRW4HynrrQfo1iMiSgw
4oXrUN7TLi6nNjgD74r60dVZ1rZ6Z+Y9liuTu+WI9GLmM9Gs7Gu3SDyP+vWmvLr3
P/waFhZ0z9+6SHN6SKqZXq/l0irItPOSIwmCoZxqjAUmuLDW7e7O9/pvUtmo3QyP
kAseGKnm7JZSlM6XX+fuoc/nsZ5qh9XCaMYe+pQf15HIUl6CYtwixstyDh8V22Z2
QM3MjS4l58/xo8CeIur+bh9h/nU86W2/HjERuq2MvjrFn88Sr/1RKixxohrZOy+y
4IUBv2ZOEUrS5LfWcvK931/cFHKSZsShfnZP8Bc9sUp3yPY9Y1umxLUZEW4Aja7e
dfBhFS5j9elBtKgK+xERmXak2P66nXWANb2aTsIvpVc3FnEPrzVlSzoNM6EN/+BT
qjXE5s2P2Yu5uBYLTHhv3DGSPIe4R99ves4txp+crzypTLzy3OWp5tfYP2bU/T7Z
RRI3M56vTcYAlpMexNGniTI5ETaUoc6+ifUOcsI5l1oW9DqxANnh+jeodnY9offA
ADSwNLu6JUNsMMDi/sn2xhILfTTkvtyg3uwC7eNJD/xoRdP4w8rtQ69H3AIy9qa9
CGwSWW28yJKnrUjOI29yQgLu+GSjNIMdxlqqLYV58Umn7WfSo2hJkvQ2zy/AxGe+
z30uwgSOBrQFy5hmxAOU9LkDdw1JPHS1D3hAyH75/FjS0k8yJ82Zy/LWlrkhuD13
PCb50pcGnIpA8WD9b3dyezkLIdm51Tm69oOhbsn25Du6sGkxge45l5OvtzeFo6iT
XNfPUY2TRO7B1LiyzDa1KLvHDJIeS1qpGIQKlNO9iKOk9FyD99QNbnAqkA3pdrC/
ULhPWreppWKKi0jRtJdQBavtySLvamQshhxM7Vo67O5JGl0mP1H4isXnM9XUH+1E
+ZIgeXSE2hlgZQ8egpqiWQrbi0ob+UkqqpA/R20D22t6WvM965SMeQK9xH/vlNh2
et8zL6jGF/H1QzOYSsxUV9lIv9CF0ztqQ8WYcHZR9IDUfjk8dXef8QBAwJkOLJm0
eR+ZvR4AXBgj1YxfZNMsRDgw43J02NNzcBryD295SfVj9Y3VSRV3n9HtzOXOs5xV
LzQH7Z/fqFl6YrxwvuYiqZ+6lNVtTlFD1Cjtm8w/ti79Xdwr9KyHRtTYzsNkgQ3B
599e1iy8HD1SJkCUtQ0bQP3GqpJAv1w7o5dFvgKLArOq3RqzVvq6kf86NKCfZK20
4CmKYy4vO+q4+9lBV/eI+Y51QOosSs+XXwaVW42TbPXfDEyCWquoTHiGRIvwqHuk
eDmaucKVZ38gmb5i6ysZW9huXHfZ9ox6uNt09vAvb0jXAMxZlVd7b/BC2WhrPXv2
vHKBi+/gC/MMWSEpQdZnfQ8+jMia1Zetc5N1SJYronmK2pcSouvUNcuE7noU3Ltz
OvrBw/9X5rzuBTmtQp+px9B+afX22kggEk+iASWI4fbMNR1XpGRews6mYiITp0aF
nG6cM4nO4izKVUBSt7+Ir4hUUeeTsYw5GeQt5y/ZmTG4rNzGR4cxoFSOs9e+hNoi
u4RkOzEGH2xnhYj3CsYTI5Fwgbj3FD+EDuWH/3hpG08mJpBHW+lcC9KCHuNiQW5G
9qQBP4VVSkNd61BLPc8bBJOv/FAhEoRDgkw/AtksE5Cy9NY8S9oBqBiJXZRkkUl6
7E273nDlwXcb3PDdU9aikr9ZfkwceIio/+oedkJ/T8debZy3BM2YM9utxTdCBFCH
677W44Ysr9N+rtRB4tyMvJThCS2fPQzrjjeRD7/sNST+0dOkv5F2qIGYOc72Q1kx
4sI5Z6EKrxphHoe8MWc6uMyuASu3mq4FQ4N2F4OD1D2hUmWPijlpVICJHLmDeMnW
3G9bcvIwJhnX17OkpCfwaQRa0Mz8kqRMa5q7NArxqR1lUZSnic6BhQZ6lqhk2CGU
6uiWspXpBhunEJmsHEra5P3Bc03aNuFS5vQBt2tQLAhTawVDBcw2lTEJXJdI0W+h
6n15khc3QpYY/pO8smomtEpmC15iqIqG5k8MBrogUyZcgf/GoDII2fgvGJmjJIat
u7VWj/hayhjnF3zZprVURR0dQvK0fLWaZ5iAlPAwg2t/02hV4yUTbOe+sFhNJgoq
lLzqEBQu3j7HAzOnxVzDqQX2hXTjskhFR7NwsGrdrpEilnh7JjkUCXaSdhwA1fFL
Jo1NOe+S75cqoJ7M0w6mjdiAwvtSvwcFSbHvixbWBnMxw87UbU5hShtD+rJsJqIQ
fPzOanvElxcFze2IQp4HMwCZsj4KwUtRLmAz2cXvo1z2sl9ezZ+Egz1oMRiX88fw
pq8EM2MM8NjzX5yb4p4Z4mdCWhA6e5BlcB/9U2JzSY3OQV11YTy9mNoSirCkm6mR
m+6+L4eN8UgQziSa5LSMW2W+4f5Kr5pJWUtJE7/mka+Pta43ETKBDrs5n09sTpEX
PQF+2R4ReTKf5XljNROzw41ZRzDn8gCVSqi61PtZ7ycWxyi1EFlagUO78uU8N5Y/
VOCA2UI3nVdyAhfB/afwQ50UQgi49yRipQuQzn3NXb6+tZmzwDPOSRFZSvM/WwVZ
60cg3Btnd2krdO0KsrVkrLGlypIm/MJruFduWJ8FfWAbaox7Kn/T1miH93wHB6q0
TK6cmVAizTGWsy5ekLBXM9RkpeYfmIf5W8zLfi4R2vxXivZWdlBTCP1a9pOmKtVu
+Xbc9QCcoSZ+J7M4fTmSR8G/IxcGErO6SkUx48e4mMyGaq63VAtta/En0RuXOhYQ
KuM5g+AcusoTrlEmZ7YP7ddK3A7PTeCCqAQOhVX7o567nKvkxzZ3mlqsQcX4nlVe
vlumeJBGMnkLbwVzM+d/yW3Fr5Qgj1td81BEuTOOBt+WWzjdSSfxj2Lq4WrjVuef
+fKbUwSjJO/ByiVlT1RNGgfiTBOhwD/nIkvrSJ/yfGtQd/+0uk5iEwqNBcyAD8Kv
ePf7dp3HT/2ZLIQoUfozMEPCuLT00m2eYxVKDpJLrOewaca++uzBgoJbKX0SekcU
zGrSBtPr+eICorOVctlqW6FKl5D0X8BbqleLVkV4J3wjzoZKLaiZ6QpukJMX+XVJ
4ci6JXYAoWnmDyoSr1kpTiB0aKil1rkbhy6Ollz6W0AxU2eLDHbWL+spWYrpj/LM
aAmlDj8VZwn1ITMagM1VrmeCG6jVYZYMw4qcFZDif2DljKTQcaQc7c1q6W6H8Um/
t3NNwiNgqmbBSqz9rwz6mOroAuoTzgQRwxMzlBZ/JH2v8nVMTDDDDKIq27hrKRpS
Jgv0IAFAPC/ZdU+Wc7KFRDfbqgoyMj8f/MzL1xwVFGCbRfR7i22C/PgGwSTD4W1r
XuP3UpiwN4JJqQqQF/hkLJnya1crhLglAGrQLwSp/i5JlrOVuTroTc8TKoBjcCXi
3jJGcy/3GTWuUmhqAJdsQRYwct6M22w8TyzDTqwpznUoU0yA2bGsZ/W+mMY9B/Eq
gfjX1IKz/1StadBRx5jDc0kFKOOxa+tgF0Jgy+Sa/rLQRoThV7sTSciZpCkPZ/u1
2gwHT1lAtr8ZFd2CYTZ/Tgzt8zU605RH9KnkJ/uUXgSkfW7APXSGDR2PfKeDEs/6
nqy7mjTx/BhDP9ngEY6MrH87ijuCQ3dGWYFKBGZn51y7ODIxLvtngSmwCQZ6tWJT
uYEdarC2FTu30UMftHitR2eEz77s76Rj0yD0qAR3UfEibqA86KD2mTAxWGzDcF9+
n+kzrRycDRU32plI0Qcb0/vdhY+5dGhOuXi5utXKLCpDC0OEgzBIQMJS+2YBmPi3
jpc+HqApqs/JOUT/tG6SrIdNGhaIRIIU2+hdJcY9dIKRNums/U0m/hwNnx/tJkw2
AGu4gFjZ9Q6c82nfEVW+mIHO3daYV4QsncPoeIRKUKzaWjunGheFhZSf5KpRh17t
/JrAv59w2GTYaJoJ2nqH/JPq/eEfHVTqf19eEOGs5Wf0Y0hcQ0gJlodADWMOnTw9
PCzGZVfhkn6rGrOnHzOZ/ceGxpt444umSdCspj9jWbU21AIDLUmnHRrXoPpIxLKb
FG666DANXurEifOUD6EgkzX1eDHAqdjHA56EDg6HqcLExSjwwrGQ6LxhVsL6x1k8
X78vu9FZsDhTl5r21DkKXnkfcftu7NqpHKmIuSThBm4LqtfK/t9Tur0Lyvn1AQB3
izEN3hHgDPBXV1HQaR3xwPlBzqNxgJeBIGyUoNN/Mj92oeULIgP/ZVDrId6HizU/
0/PTdB3HA6pEW9lw1HpGJoCYhpKNIv5LF9mJ75HjXazf+5GnXRxneL+eiv5rGmhf
qvinlflGbWqpuMcK48s5dKw+PMJQLQWe1vEnNCulvuHb3G9QWAvjNQsxAjO7a/3c
z9E4fPEKRgyUDm6gTeX4qtDgjKLamEeZ9kCURlpjb/JKMhiFpjzM1930Qwl8N/FV
MWZ+/5jafRyeRhIBWbMCtaXmlA08HVr94kQ8mIlww3RfDEbkoGbosdJQV8w501Dw
KMVuhuLoHZtwRPqtweb3lyVhhcen7Tm6dn/yH/Kj3DVk6k41MeLusl6QrPMIt2HD
4Xri29diYWggpbfQ/Yn105/BCPW4z8NY7VKPIZLiSXSjP5J0QVjI2bPR0+DjAKhA
j6mJvJmaEXVyr1ECHlQnQK+3FUH2RyeD2iKGpRCxYN0GLFwwfId6rGCh24fePpes
NKMc6DsbRq8KyvRrXqhrdb4jVq6MxUPR+VwEQpNwrqkyyrSnlc9VToRoKWXDE1rk
INdNW3n2tonSXzgoDC4qidywfEVHL5hoJDCeuHH2GbnOMe5Dm9Jt0JEcwpDtpBC9
nJTD7vC2xHaE/H247DpzUrby5NFCju+9H/lsBW/nAqJ6WxSB3D0F1NoLwkIL+BNa
qVxf+48TuLIWfKLgglLRywQsvpWfaDDtt4DSHWMrQwdwqXGWad0lfoBZW68KU+XK
2C3sqmLCY1Egtqpf7Sco1AOjuL4XQOYqo2E35ldSapYnjPA+7Ek9VyD4KkRXofgo
OEDJjY3+ngFsX/gtuXmZMxjmIQorjXnX6BkLQGrRh2kvjrfKcwouaC0EYMhmcDHX
mqueWGQdQstbsT7uv6kUfcYFYipWp1TxcidK44aMWqvfMWjowgVLEbzA6ekLKdiU
jm4viN9XlKQ+zbq5lu6UEm9e634rug4slPX3y3cIxylqiDvN3uwqgdW7BCJyavQv
BqsSmYIR5QsPW/iQ5Kx9jJPN0tg2nIIv1SFLnnqscZcd0lZAvk20Kne5xuw/0kvn
HiUJAUDYupXyQkxg4fVgX0MWbWJQFofrOTgt6sHUDmAyYHHTflIr0kc403HDccYq
CfcqmdF0vPtepdLPRg+NI0rzEpfhkPlSTaxBe6UZ3oVmM8X89vgcICLuRRJGiMEj
ZPVZAuHzaJAkHzutTWsZznJw6sPz6mGuejspKbkiLgi/Bd/Ro8dzGr1o4NdetZpC
/Kip+ivGq25inM+NigLur/tSBIlGUairTR1ObPsI0OU/xlTEI2INifzJLjYmuDYe
Kvzhnrv51Vj61oJewXNKx+pxFBpp8Z/Fx2RugMrOq21sMg2Q01LXsoH0C9tYBTTq
Ourv7E/6ZJ8fRDoyYps2/6DN3DdzS3kBakc8YYTVCGriX2d7HFI/vGJmSLrtHtjl
MU39KLJCLJyLKOC4MCNA1UZez49HffR6lct8LIdvfdFVITWFUrcu+KuebcYYQgXK
7CCqQQmXlCuvce2yDXq+JVamgyULrE8D34ZCcHNjH3UMTZILPEdm0d1gP6hjzrDw
fa4PRElJ+WBufvsQQSzDU8mtkJSjcuJ1edbN4I040FTZLLueQ5HOTRGu+s2pK8cA
OZ4diG03RiISYpuzlCSzNC3hU6HNBwQQtpUbvEm0NjwRzaXyO6OCuBiYCWU86Qcd
GuKwZRU3esm8sFuo4POQWr8divQIpGZYllNT5UF1mLtZ00eGAZp60+ed6ElfgDop
MlcEXJyu2BQpwskCS3rD/qNNijT9ofUSmbz+Dus2dkqlKL9D542J1vS8QJtt9zpY
I0HKb6jMPLB1ug3x2vpyPewjGJoGvHezJ03n/jAgMbhxCLm4qrgtYrbdaAVwiNsE
RoHF727akc60hNN2A7JdomcVjdrQulJxYSR8uCtTJGdqMF4/zvwpnZRTZKZkuetU
ssTlwMHeQWMd4ZseaShl3/3jaUkFVRNozEIt5au0vBdK0nub0QWZAJix3UT/uaD1
R62YExfxNahZsm+ZaHPysTZ7m+v3q2Fextjyt0rNP/YfiGCg1Bigaf4CpVWLLhNF
gT8LTOC9riB7LtLYTdhAqItUfR5lyZS5zJAANkYY0V5ZScQBo/wwZbAsW592Oj/L
8ygg0Sk27/h6xsrss4Kv06IrTavb1u38lw4JRh+3kr3/We21Bv8boamJdXgXASyK
y60kkF4+rcpB/PGFgzNMqP/XzqdrZPuX1f3SA0Act+B+pGo9nAevifQWUKpu6Uhv
EN7KNRKwVLeCiAmh/BcVJ755ceacDpGPP81BGprThVcpFgidTCYAl1wxvBnDkyM6
VyDi7p9LrI2rJySmp4+D1qKx0zoMs0ZXc9EUcCLbVtD9TSsmUfZDaqkDgaC5m5ql
mJnbcE19n7KbZR3WHZkvl13sXPYBNDgdavFugwR6NK6YcRj7TWEHZTy7ywFt4kqe
QsiGp6FqNoRg11dP+4P9phR0Wks0uYPAmBAyOiqHhTALv39jx+gm1+utgYYFc7xl
tZ6pWeqvHi/ClXbxy4nyQy6zUts7t8bEvOktQM0bZO3ezfHA204IjL+nE9Q04+gA
OYRfNLfih3BYLrwoxBsEoKsqmZ8MWLC39h5NlMJv5wNVYfPfLYwET0HeqcHpSoBR
STQ9hpSIqa4bZ7xmYxyByNESBencsaMTVx9H//r/XHje2Q94Vejx+ADLt8uFoG47
xXtTVJr8np0Zds3uscTUvCsoQN7p2ujj+z7asey0v2vVMO8opQ5q5Kj6Tjw0APii
Wb3HS5eidxFpLUjV4FPYgeYIWQBU3z3129n7uQrtBE3iojMjmjPrUu/b+6IsuzhJ
tY09Zs7Exb31HjF2McOMSI9DGSE8ZyPsjD1HsdCsc9M6uBfRwNN2sf5B9AEmwqvH
IArcxOTdDeJGpEvI/NovKkZCwX4M5Fr96slXO+P45MV5PE0iNyxwXilhtOi8n+bm
UCumZfUoZ/ZKzXpFivW4BZP3gGtKTTipEbr5SMsv8idUv13l5H8IQ5R9jKkEPFIa
oqTk9/IrdDdia6eW3ec2MF4k9I1RB4KGbIv2JAXbnu3rgnV6uNNBe9zA5x8ulk1P
xnHZWgesK+Lc0UmAumo6aQ2huTZ+T/oZaqvjxTBTuLE1Sc7fgX/STroBF4YT6Eu0
mOXrO4jYhL/obHCye37K6DboQNJz7LuurkIzWeiaPXY/68HWNcMulpdLo9l1i6Yx
vm1nknpn4FlzYtg5DUsbzEKRRqXx2YER10zToHLTpZW5y0ogK+5ki4c69Uqceezz
W54zDRxNYfqraCdf9lQcW4TsMykLK6bUupiOYj9DFsSxp0Apqw/Sk4QZA/SySmkm
ODL+UOsx+GfG3rLOkhE+312/NDlmkuU1GvkP73UMTm1mwoFKUVokTS/te9FFPP3q
AwsAPky+c7MYY3YK5xiGulpYJ1jZY7LlS8qyLP4CiZnp4hXaVPBaSLWZBDaQ2+0U
UewKI8pCDviXt+VOoUsO8Mr/lqJgWvDRyExdjYnUoP1+5Nb1E/crdUyZZqQY69BC
TzhWP1Oaf6J0idZKVKeNdN9d6mUepcS8fbYryFhuoELQoScxJgj9V0T7jvApY+xR
ZlZ12INzZWKqQRbcwMOS4gDon5ui6HJwHuWxwS+6yvVtbShHwhijjS2taReoc2CH
jiQ66yXKrhABYSNFzKRvNY3WcXF4KCsYQj24qtMl6/GTrRa7TNCXGbo+/2pcqfFz
YQ0qD8/ejksI649ySBSlFnz/PY2hReQGHMmFX9VDAgqpR/0WQGYKZUA/7ZmB4RoE
9iyX82HYBPBKBK90Rdws/HFLHTVp/j5c3NXUCNJ+m77Hdvko3wIY/IlLNrPP1wn8
PSb71rBIrt5OZeUWfuhK5rdRl+vgZxLxzYtQbxPa9qamed9fNQThSxZodCA+wKM0
0y2r3z9nOKCpT+frbFOgV8K4PajN+SZu5Y8FxMBMsFWiFG0JYFYCONdwTUIz++sP
Z8/w/zD7PXs3B1I7TUb8ImxTl5MhOY73jAp7DZhk19UUS+lkkdpbdL9pEj8uZh1K
PEsbUqL7srt0o+M2lrqd9rkoekSHz4eYi/O7rBzyw53eHnHsreBkWxse50SJg7uq
+Q/r0LbdsHJazCc/SiDY+kttqTd0I3YUAI50sIwNSMwK0hHItdwxVJ6a/YqSvY25
UG7AoJ7SrH7Y0WmY9KAeU4/HlO+0Q5Gfju92n2I4z50tUDdq96/FYNfUJU+zm+KP
FUMk6gg4hAr686KbVyHx861Q0B+tKrBF3G/cuyBaG+DuPjs8C/bK2nmAqog9stL0
t98NQKpJkH1vR3/jYzZdl1TuetbCBCSuYk6oQ51SeAhs30obDl2PldXWdlShsYkP
/y2OY9dC3BqyMDAiwyW5FbFEQ15sR2ftNfgotHZgn2bnj2BuK59JByaq/9xwZcUm
gkorWwd6eC/MrSrkeAyuKYm26vAe9BbNXvyu40Rs8l0vr0GHVUhhou0IwTV6w+5b
CSwAF9bn47ppnmHWBNa2MHqlKWVA+T0XNDIWvZRzvP5TMec+HTqjX+9ZWJYb8E+k
mXmY/NmFmzv1sKBFl+ohNFYVz65wJ0B48rgpu1yEbfcRO1P4gPjdpQWQMAVVg2Sh
e2gabHpdw7QpRxklin60cVx2tcLP5dsPQqd2azzyZvVynmnnnOuMsUoWSlBMeTct
4BgGra/P6GuV38ezyFylDiGnCJPiJ/TlTtX9K9tUdfKGLZvZ7bkXbEYJ/fZrBG5r
aBf545GFsxwjJZWN7PjRpcEYK1asr6qji2KIRU6Sw3EGA+h1F9M/0f9b9wcmPp2x
a/cpVn3Q727Co0U1yEr+MrvUGcIra4pCetTz9JOLWeBHJye7X1lR6jQ8dq3Kvj6J
4RGT81IsPgdD/ZgJmOI7WHiFQDkpn2S15CBEJsZzI8VWsEGe8HuQdewi0UA+uaB/
ZgWoiwiYHrhdTWgIoP2KwEKWj0jVmsDdzBtgvSm0JcpXhOOlzBJnR5fGvg7mqcqY
`protect END_PROTECTED
