`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GSROqoc3Hpf7cLgmJ4jM4+1RYA0T6a7klnyONKfSMUo5mCo04lQ8zy83B41olFD9
x5cDoomWR/83CtfLlnMm+dy4e+KTUR6cxwS4EwTkPIzHP78CYJxsNpQHIOCt8Il/
/8OlUlhAeiVXqoq7jX3IftaQQBLQkphjKvIWO0kGRL1mP65ge10QQUIams8o+FnS
RyoFQS0DRVp3hFngHoygGCqAj7vF8IuFJ4QtyHNr0a/88c9pPx+xvhBIT/IF86Pn
7VSSDYKJaY/+gzCO2msdvivpCbJmXB1ztBIrsxb8EiEejk0PxexmLCqQJ2xCflZJ
3AHnw9YAHz1JNUTH6GnjEEHR1+WJD7KR3QElJfWQk+uBSSBv1gyjhxnxk3XCMytP
ALyEF6vJXEvNoprI0d/5Zo21wr50eflajIyT5qNsVZxJNeIegctBFnDuJYYkFink
Xx/K1TO9nZadcUogzEJ1auSwg4NkPmvwvtt7y7M093t7eucP+L8zUkAD2faPNJ5I
H24Z+6bv5W83HVM0ESHX6Jmelrl2YoFTzLIZ89BeyCS3cZdMbRHepJt0wNbkBHd+
W+dKNhvIXlBTbVENg5QxrGju6NRd1RYE7aV6pg8YL9VOZpK6/aK+q8RxiTWxNswM
v6XHs7lBdOpJZtU9txImUvjLMHsa59Fwy0Rs5DnMSNsT1yKSnMHme3GwggpDJHCU
BAssX+lYklnUdQeBi9+jOP8E6AKl9csMsma67hIWLkb65Biqc86QxYkU175ax2Xj
5fJPgc2K/ZbgwDaepG+lAXJqifBvuauNxnAp5nYg27R6ugl03dSK/Cot21S9jxsT
iWc8TeU2M08GwxrKLYxcsMwsgiJfT1sNPxOoXx+L1sj6YTzcv67XPtW7OzFgmtq9
UE1/fhSNQ3cP3TiNXmAVY0t0dfIU2HIUPO+UKWUGwmX29JxD64e6A9UqxI+C+IdP
yBHsUhuNc05mpVUadFZbMQ==
`protect END_PROTECTED
