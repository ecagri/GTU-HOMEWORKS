`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aFD3yz0ksPKxHYSR2xLeFMOfzFKDvEN2H61DpshQvX3lh9b15hpAa57R9lugvjdO
V3IVZYPPmNZdp783UQ2KFa7uajHNg8ZgfTqArKl9ucQ9CO4yrXPExLQqr6cQe2Z4
A3hyWHnRUfuEIV8skEBq7p4dlXO9SCf2ee6lZrZKdcKEwuITw6pT4Y8q8PSm9lim
xn8F1h09zT0x9gH3irWXCanDH06O+2iiyR0sdWdFjqJOwGzLO9uhKQo216IjyZFD
66jRYxGzUVVi777Tw2CMFCeysedWOZ2xX9XxrnVyXb7EHJ6en6d0j36aHSVFzuh4
UVVOqNv3voGg5GExh3JMudl2/HUE0ZEQm4PQRzlel2pqIxwvBtk3aMbikUhiVMMW
VAc/tTjcb8aJOm79+CSRx9LwPZf5bmhY+I4tgyITkTEsF7fb+zDSiDV4oiFK9EM3
vquZppletqKshVSscDtp9/5dWZ5elPpkIvNj6bs9wGZgEqbCHKaXE+9woJVdrDap
9N+NzkUYcTAZaYK64TjxVmxch/tnkMOsaLplKvKQ4q4/ZRxvXujBHlLOnPhDv8OZ
H5DmWy6kPAcyhR/OgRaEth0BwJa44fFvMIgBO6GTW6UpFE4cMjeq4qlgzkFADU1W
MFkOLXEJGVdc5g2i8Um85TAWMjc7aLI+TJnN46SW0FZdZ1VfVSdzmlMZJKSolZir
+BfjfU88R55JnSObeteRfmIKQA6kKRIfOVWO2eRTIEVHudNLcWUdwqPr0ytG90Ma
Ue7sLEOodTm+im/dQfdP9uhjLctXfCBiWcMyUKyOQQ7g923OyTpSXgH+IjDKK4rw
I6jQ5DhTZbGj6EFFaJLoemHqMrPPOEcK9whz48730VcrJYm/gU8anM3zs3Sx26Fv
`protect END_PROTECTED
