`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BpobMBnvym7bGdwKYurBZ4zxKSZgPD3X6zlfrYBvtay2OOLZb4pfg28V+obj5Knw
XkoIZ3XIqKVmJWqmqqlE+huGsKLjTucPaZDSBr5Lr5R4OIPB+Db2bFc9YBJM9dxu
LrPr5Fnqyy0G50lIbBzANOsAoJLBNy4Qouuovv6MOzyLhOJO6/3wA2w5GMxHcvcc
YUMOwEcDUSzWYLg+Ei8TUr6NG/FJN4QTpQrja3YZ1PP0PRpYL+/Qy35YLaMw0w2O
pF7wmaC+5jat/Z3M24UjHlnSSWGz3KRY9wd4wtKUZCJOIFjs42nZdR9z7/jMhqJu
nZ4ZmbAB50lTKgvnEwNgRzavKMjPDU2X3vCydQz7v+HJ/45TfcuDlpNqTmmTOLo4
fT/h8YqEmkGUVlcJGbFjrCUbt8c+gqEme4OVmdFrf/TorqYiJSarxCvyOjWYLM0l
6bvrBacrrdk9mX6yn+NCF1oG1OQAn2BotzMWXb5AvaaXrOo9KO5RgpckRe87fgFs
W/+t9S+yhbijoBFyPUf+CTGqqZbejckvCnGqSJL6DPd2s71y9BqvXGka033NHPqv
6xFJoYJ2EyQOld0RiBZvbkPE+Cqsbn4dkRaztSXgtEhVzEynn+5He0YWZeVepnpW
B5joo3lfP9uA7JU3vow1gAtj6YORNOcxMyUZCQTGQ/I5NwfMrVj/uLDPklTF5/pD
ssWCa/qmS6zO/nlQDV8Xee4clOd4BzAm1PPw+x4FvO7ySfRjZW78owH2FiP6xmQs
Y1iyqTvwPsprA3kdUraX7Z/drwJF5qQtxLxBhDYHXIXg4jd0YCgX+FRnPdjkjq+A
ofZ1RsmVC2UfmCl3fGPRt/vAUpetaaEjZsSfd/SSRFDWbsM7/YOQPmkKPkAJnxLR
/ElFwKpdfE9O6M6rabUJx3AGILSKoiitIsFMy+NrHUu8KKaIuoS5k0bjsrpduZrw
A4U6m7kkGRgh38EfIbFLGYqUsIn9grFjDeSvbIvspsF2lCAVHtIfb52GR5VRl2bR
w8IT87NtC7kM+0EMIqtHU4ps5qxlv02v5bzt2Sa5QHHrPr0qcYnHVdMZ65AdtHVL
AJNM8GVikJ80kotNarse+dH6UbgjFK5fGItCj8HHnqnO5B/hndYLtXQ17282BGpl
bYjTfn0N0MN06dEb7T3qaufA7vHeJ8fTvcD19zARMayY4I6MMmTGWFWdUFB/dcYW
+MbOQ2ksSsQxuX8TytCaY69Cd1DeCeGrXrMqwMT3ApfLbsqYB7PkXU8YubcOLrRR
yEAqoqPvUAFX2xtWDVrNstqqiqwyC+VlD7UKAEkjPgcYNsErhAQgnKVCLYY1f9+1
+tdwGdnw8Zvzf0+dOtYuyo+aUgcsRzhCwRm4i1kFCkOUmFDa27yXtTuWRwJiw0Sz
k82aDOEU16ne9SLP1FybnlxCQwOmbPsRU5OEcYNRjD660HwosW1/D0AYtfXO3VrP
I2TiZ+66VwhBQzDNx/jt4qLb1DZx7HPl/UR7SPv/NaqittUmLqzWvpQQHgV85rj0
GXIQXROhVEPpjTHk9NdUiPxTzsRL4PiIFrAjVOob95RJock121JnvF4MW1K9gNtI
EeG32b+0h/HhJOI6HnLo4If1JNPQDu9thtWQpKXntmIB6AKRmgOIi3kt0Rdepoi3
buIPAKGE6+eq1gVcHo3hZiwAQR/VAfI+2KayvdRd/aD1try2ckiPJ2fZTv+24Z5/
CpKSswCz/PdO8Tb/EK6b/Hl4Cxr7ba29to2c2oQE5jFD0k2T4L+ifLZ4OMxThZo4
iufdQGp9aG34jU8GWwM/Jo1WzDp3jvMOhbfP65KhlRtN53Ko41znzvU4rS40MWgJ
9odoN72wo/EjHJZNB1ZCBbm5sg0/Ptj0A/LSR7p0M7+6fc6oOsIo/5GJmN9G2eEX
c4HR3r6T6gzzVhU+IIUbOZaIMXsd+hmq10hF1mBT5cle0MHlD1UtqiXPLYzxfPNy
BKZADCuSx196ahQ398avwhyQTOTncPc9nwKVG3fufQ3mIdWcFJf7eilGatD7itVm
yBajkg+JeJZkxIfJ7uHT6YWNqmwNRFE/Kt3PEp6i60l2/CjLzDAZ1+nhafLUkqov
L72fkIjMxFQgDWC6lUpI0+pXfd4l4BJLcU5vYw/3nzdTxwGZLsZEfGeZtFq0HaBr
b4iVVAjXvQw5WGUWoU9UyH+jn/paD3g/7B4F0vyVyDf/LhbnYUFoXsz3nPzHWu1v
/RTuuH9DzDMQPAKtBw4xftLIK9PM1+0SZtEIf5w7XSpEHaVU2R2P10PflBlmdc8K
tN9NFJRL8eurrkeoYHPjIHYs6z4pm1JNyxfHqn4LzUH/9HWznDHvLGoyKh0RrPjs
jBeCQ9CnYFnpj/462BE7dEB+mZO6hiB/OvhE+eIzIck1sF0j8EwLIOuXGVp39FKl
ygah+HFGuv0OHJ7tCO7GYJWoDU00eWSYfbdZGr1tg6N0vtDfcnOIeIH1AH3kxJJV
QXbCJMrvCOAZ13U0Ru7dBvBzq1sDsONgyKb1AerBCDki9i9ngKWV6ENi2tXYT0uL
Y9Dy/eVl+KpOaB9hA7pmmN9cF39hsY8wV36IV03wZ8pXyXaY0cgq6aLMc2QmQa/e
YtZhUYqzxd2lEV12YrcjvNiynamMl982ClBSYkQtkFmIZrA5kP1tM8X7Ue8oSi4W
HCt4tanOtq2qs4lsVCpxCeU+4nddh1a9mq5qzKGbYM5fepY2nRadtdM0svIHIv8F
vIS2JHj05Xef3j11DWcv2X3Vqc/otjHVs+wNRIhicPywobjs3WNqJxKg7PjfIb3S
iqJH+EM9A37QdnKS2UUbbWfymb8/e/RGR0pYbWZQm+O5PtcNUPVXNj5Oa2VmG3jh
T0IcjfmC6GlIgKXMlrts08DtX01V16covewB/7Jw/sxPQM+M9s6duFWXSwUnxPhh
UHEql4Lkqbcz5HrdqBXhpworkSiv6lXOQ8PNX58vRLwRLgnx4eKg7bD3V0aP4Cve
Sfu5GglR989AsSLjO/ujV+ObGCsn+AXvzhiRNxooOwBf7YQsBSECDoDpTSGeIZc7
DXZqUOFmJttkg5XSKi3/1GVUjKMjpxFXtta1XDyzKfl3N1rm83vpJLj0KG+vw9At
HYlVdFJ1jXJ8cEdOQe4hade+68/rIom65j7VAcxOqXbtavZrGbyDppBz9XWDmlUo
o7TJNfF/AMc+uNsQCmXd//2AOb1NiRHpS20Y6iiR0F1dDakpIC6xSvYkcpdcCbc2
a0/XirgYX4Y45UsgMM3MeuzKGA64IUHgdx3MUtYMNwaHRxklTSw7GZiSF6e4DAxA
NTsWHA2BPIIK94id1rC9FkxwdaYjmYykTnPCnvHiT3IORtUbuwLvm29XsAitSmYN
8FjKZsmesKz7cGi4czucFYYJuPYUulGHe9udIFIFIVCJbjspSKWIQacr6w1Edjnl
4obJ12fbrE6Z3B9KQ+xThWlV0Kcf5iCn5we3XsGXVGW4kqNOhggmUw/hIKI1UZEY
gVDVdT6e17yrrOuZhFB3cNA6k3YBdkF50TcjwhUC+fQZXlRF99ptceyrMsZsNvSY
b/ka51ddJuVOvh6jeBuf7is3q5suLJ/ZsEdUIAA1se22kZm34x1ui+9d3aiJXfxl
u8UuF3F/nPjeOPBhXwB5p477nw0mlicjuaiDNWi4N8VFAIHaqz6fH8dNrhgK2el/
`protect END_PROTECTED
