`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g2DPMLOcJxuku8eFncvKl52TxGAA3DLaUvglQPEk7QHZmjOTGsnM7mZ4HkHne0xV
j9mfE+QuPIsMViuDyoasrzNqaaz2DV999hIVeNFUOl0m5hcZnCLq7/y30YXkTQo6
8vAO7pmn0FjPfZC1B5geirIJhB7soGJ2R3Agg+cfwHgzUKUL7QHM+x3Rc1XpnsUe
7BXnSrXVoF62GK1IFWW7kW941ITIfVfZRFaTE373bk12h0jDtlWqInr9y0PBX2Bb
xme824wEerRAoyB6N/15q8lSMb5e1f2PbmYRpwJBoCA5oUhrkAMa37b8QLvE9kQH
rAxAYZx22c/paNF84g/phzWEFViMJ3hith9MJJDbGo/l4FUDQ/NUBWbRaJ3cp/HY
fpJjTrsgT+eGfDIj546HJTZb+Q60PrfJtKhcOw8pWPnG0g4uYfvTHo6KwiE+2wNR
MLE4WpiuF2vRM0y7ImZV0DCYE6LsRBpkPcECHBANaEO0Q0uPdAbG08chenjGPxef
j1i/P5K93pdp4jdT/M9DXr9vtwPS1nOHIvtXfiAvMTg9SbekIw2d9Znqe8Y/2ZIM
KfLwM+5sG01lfMMjSwnmzOVNjYB4ienIHwNgLjCjlwGYFPLNsFP7J/DOwSBOnciV
CQntIuixI4F6dk8wSL7q8biI739WS3eQusrqtG+1FMMhTVpU8IwCj7YGln+n9wnq
lEpuRA37coO2obGVptWaquYW7u2WKNLWB6DBKTlbSUsJogiKq1dxkTHnuKh1BaT1
NpRbW+lt+8h35LzSJT23gvnrb4dy/7KzVms0g07/ibbqR6Gz782MgshixNX0KNvV
Q1llKe3k/tEUuOQlERfPfiwbE9f+SXYKU+0K+S4xA/su0Xkm2Q7a44dHJ/SxqX/E
b2vO7bAE6xZ2jgbreXx22tP15GcevvUNGh/FqZOkwPGkGSGr0uijJN0p6jr0jRez
jU5EcLf8DzXtiJjZuQgE6AfdYCG3uWo5MnNBtR6ORmaDWnB63CsmwF6+a8G/83uq
OiHRVdlFqJ5yUiejdNR1OpfrXxC7NBdGdPVhmdKIx54RNiHRjO9cxGKimaAzpHKk
1UMSrNZXoWG4BGjv2rkwyQ9CjL7QAappJAEbyVatdMb4Ezl3cYR29FK6PszVF81n
Vvr5NGwDLUhmiD87UmFojr0LiedYukAAxRxMvYHO3/1bph9ESpWc+IrPT2L92YSJ
8yFIzkzckrHGA7p2z/neaWkJk6HtQiQdpN2C3qiGNRxiEIyPQSwkii3pLJou4PZi
poIWvIDibOdA5eJrkSWCXuNNJsfF3VXGI44PZbAs06mJaTY+8VJ9gh0lM9U333+g
mID47mKKT5LiBQktzx1GP0unQjsTZPNQoYS1iZla2upCkIY623Tin3wIhGqIDNgY
Po57CS40K6wX90pMg1OzTyV5fIWHRUB4jGpTHQJe9KPtdRvP7DeDTzmAWTHUE8mC
jltjCSE3y5nwMml2v0Wpopp9Je56sK1XVRijBWKuvB09cyPCzc00L8Or0ODlj0b0
ZNWG/imRDIGmTk26Uwrf+yW5OzIqngJihxXXgtny6Up/0jiJ1flhZ8msetERsjCF
IZYv9CceyLUZVOJ3hMoWvvyo6eAcaeCpMp/bFbGrBzdkPzWMnX7C1564eCXsvF7R
iySi9AoVP3fGlEolM/ruiBzfI6MJZB2urHCqkYgUZpviX/iOwNCwmd4dQKwrL9Bh
DvBRPOcfSHRIRCabFWBxGgR8vdp31YBRiS04gwa5A67tJfV9ujVbe3XrwU+laJLQ
sAAOOhjbtqwew5zoVzEkpgekPtywMAfo3Bq4dpdZ9rxvaZb7K4UgryCanY6AGcY/
cysBe7Quvq/X7IMEZHg9qN4QB9TxjkJYle8GR9fa+wIKIM+K4gG2Ho06eXulOpSX
WKwIqOPqCjfjTk+AnL+H5ysD0B+kH1xVXAhxFk+O7Be9/qNRBA8RmpiUtuEPtD7U
p+M5uFS0Gic6bNVs7oT1nylEQRV0Q+M92prJq9VEDrbFcDNhIqzXJfF6zBagAxt9
Womlunjznc3/XF/7uJqKpnKh/z5BhwZDiuOzoHlFwiUM+Xtl20PRkldLfZqXcBl3
4O1+hp87QJx4S4BH+ljbhlbL++gM3z6jHjawyPmA31Z9MAOO/L2e+mVYP7INQlar
0hLkF8SQ/+vmeJlL/tvhO6WLnvqSLVG0uU0gECpilM+OrJus2x3D0s/aHKnMnEgy
d1F7/tPupjZHr725bPJSW7i0ihXo7TgDNoN4YMiNO2oGpXNeWKRkCGDFj5jiOEZm
FEw0TYz73AbyHMCZouL0JB7/YuzGk8lg68s0HGYcXe/6piuKLN5iMDE6jMBUAhr4
CIosnPL59IjInIFt9703Z8eZ2+05Teei7D8rcjmn5iHLfLZ54lnfSl/+SLQW1IWj
R0cJoNJ/gV6O0AspKRSKQDXE5qLF9wXz3FXdJEMlIuYeH7frwvkCkq+4R+3ONesm
fsyTCp3yKD9FLb+uqboZP2chuoI42aXoRNaLuxXtY03Tz4ZRGioayEAyMtp3Tmbj
9JDkQxu/sPZjP0Z113Ie2NiGhNUFhr5g5GWiwtIl8gEH20zP7xWDkROs5rMoKRSN
9M7EYwYXTK4L6kHegIlLf/vP4/Izo33RLq8rSN/bc4ShDRc+q7xSgaAfMhtl1whf
Tm5OuaYWR854wU/tvnIOXvOCk8RWTMd2xoKxhvFs6TLSCqhLPZdUtjhSYJseld5F
`protect END_PROTECTED
