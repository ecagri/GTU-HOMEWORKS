`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KjpXJ7LyJZHKSHO3T7IridCd9KsZwgnc3gFtn20+K2NSc4c7ow1wfu0QFBZRyOqt
0zz+fIkrNdoN3bvbt+Pd5DdK0HJLuBezATn23aejmw9cNxjnHuuO9yPEzDw2hu6d
DQt6BgvHBVOYZ8zdWRVq1BFfmrDVuM5qMeKhxhsYs5is33b5XwbYQNIItMkeWcT7
PtumIFWQZ9Z0SRXd2yow88ulBLt0lT1wuBcevGoFmQCC5AJiy4oLDIAjCvKd5nxN
eJw4LMbEGaTTZctN10cV4631Nmqeuq8aMqHkkOyf/q27lsODYR9GDyy40Ae2I/2j
0Id645ZSdJHDgdiSmmZbySg7uTO95zbnzXssq5WK7j1n+Fhu3A/lgmmZWCVUS3Gb
b4UmCkmaJz46WQWReRPRAfE4LwGJwE1o4y7O562o8KZSd2w/qzFaCI5XgF9q6reP
j2LVr9Z+4+LvShEr+0joNshxHKZRmDT7r40ARGZfQ0ZgDGOO+az4tXHj8K/Nh/WE
8GykSZdGDUPnIpC106LnNPCcDLijvdUnUZW+Lld2druZYPzrWRUTeOEOOA/utXun
vsfZZ7JmcvbCR5vXPjmzSg==
`protect END_PROTECTED
