`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7uL8GjvjKcNL53ewq+zePfo1fq+H+vjvjnmSSBOGfXKzBiaYGMVNYW62LEynWqe8
R+/5lzoesFmWdnSrWGaBKpAS7rn0a4mH/2DNMjJ1413yllrGDyBtPE6sTH0RiR9k
v5OB1fM/lqk9bm3kMwmonOwJUnYY1lw3xVIMxtKblg875lp16errJ9iqsaA+mFQy
xLf+9wMkb8+hTb6qkM2Aihaa+2qMuGrxRRdfdjhn5q4j9Gb4DQOYptgZsJH5qZ0R
4/QKV8MD6TYbscGNntKZU1acspQDJFRYoAtIjoRJaLV9RuowgBd6XH/TTsWGo1QU
vIPa1sV/rlA2gzp5nJsNZAZiOwxBkKV+3yvDrRGGkPBYsU3jZTPOUlD2QnAcoZh5
PTVAOBCuE2VLG2J6MZS16FGk35Sn9K12uuqmy+3Z+r97vnGIS9k99zWTfd0o97TS
kt5ip67+CdFbb19r28fXjXEOiJwfRpi0daPqoFYzLh3F/pQp8W94zpdXVlg8lZ65
WzKfRSzRODRIhpxRdtPgesRFJQhL4RVajCkbIYWAZ6ANHvdWgt96LzsjeimNZzlS
nAhe5JmbUvfXdllxTdtZqXCDiOHxoAA4VZQO+q8+iogkZuEZvud1MUtEvy4Tqpct
raerV0pRxJyS01fckRC3UvyAV+EVLmk7Q/XQU4P0/IPaYuSwkh/m+XhofXZERoRo
YF0fA79i5ioUcuYt9tcNVlfkKa/o06gdVhRdLu95qRPRx1gGEJKv32wUYn7y5FOB
b1Ay6ZnsEyWGKVvOUkdBJ0VOfAxIUrIAzGgprWuSmMN6CXMS/qVRgjVf9Aq51qY8
Iv79ORd66GkvC5s193bAfXVc1yuf1FeaC1klt0uwoVtHZumeJLBe+U6ntInP4l69
ZkB7nAlWf/vRa7UDlvm+LmsD9MS/8iMYYFGwrTIUVm2Smb4+aSv3EkGyOUQSNd90
KtREKD1JB0cAqSdJZdOIFvwZ7BtPoLVY3c9Sop2ZCgZDYUIm3NJP9IqdUNDJeFRs
e2gDnl3qx76emCqRX3JNKHERo2NOhD6USEzJRcJ8NC4NxnkeOKQ9DGi9JcEc2PHo
ZS5fIGh42oA3Y+uoG8dr3qC9iyQZyMUDoZ6rQ/0xGzc2i4aKpdrKi59YDdohBveq
EmZRSRytwx3vUJ1XvmqjKwxopHNMBMig9Y2SiC7ZrAjgVuXMRRxEr3OEY1WWr8Bw
gFIpfuo+ynKb4dqEi7DOHRv3umBOTRoUfTxAfKaEuQMRhYhYSvkVXw3MjqR+i/Pd
z/jHKaep7sGAXK5Bdci5DqtxZD7xvSQQFeibPd+LJKxdbSJKZenpDehW6NqQRVVO
TY1jEJa03hjXHWq0q8Z2q/ZMJvNYIsElYGABPaS3NJdlXb/UXOpeTIRUhxcsFz6G
NEqCV2EnBr8MXiN0HfQyDffol6Ugq1qU/9F7RTLCg/6EItQKGIKsAFsDfM62Yd4e
Be84xzW3JsGhOYtAaSPWoEcc6WJhTEUg+SWVkpR/ShganqXy1y4B6UW3o4GYTI/C
OyRdODLgjcP32zN7Cmlrgj/koiXSAh67yAY0vO8T9mPo/qdyLhD1Wq2qNqeKfaPA
O1Z/30W+RtBiPURDPJITlQrpr2alBu+q6S7GkMV3QFbhjOpnkgsdgD1VcROTfk2d
eFcf4zwQrUae7OLMSzkUqpnOcT7AVtvx0iUYcIJ3gYuEyPrtuzOlFjetmT5jaEgs
rZNuReiLTwNleC154S4z8qZg9eotVs+cZcoEifqkAy0DICklh4PIj/CJ3VabP50T
x466AhwjrtXaYJWdXs/+PfJg6Ub524cJ+JmF85QJSTGquywYNYQ57VmJU9dVypi2
WRhw4VSejAZBwOs0DaQohxWXSpgfenp5h9sww/x6PsA2kgt+bkIiTxxkzA/athBW
SPDcGFN0wXkLn0EgWUt0/4fMXFqwxgaxeclK3Y7mHnlrK+m+39aGjhaaZDGveSzE
cNwyh5rJ2TuC2SlT74l5PwWYIgFYTWLi0bYtiAjaBztDe+mOZDtKznXKAC4SWC2p
VZBmhMc9oXkLGL37LTQI/Pu7HZa7AytyxE58Am59aytihNRBZ0iod1F3qPN8Ei4U
gVCNv2vN+HC+eT4DR+6gozh4sBmMpUc3woQVgZ4vQ26Y3idI2aQUK1DB5AwM4rKq
s6B0A4My/XcjDwlCjrC2gAXTgnCM7XG/F+8b1Ogv28x1bKRDw01oHaLAcc3XEp00
FsZPkw6OXzf/Eak+9aBGQ15irItimudcbZ1zNjM4w5mMEhX7cWf3L+2RFBQMQSSG
jMT8W6P2/R5cPgGSdbDtz1m3hPMocNgA8Q2miAwrErY/sXlmPjEbmzugnftgssr/
MohsE/FYH/H8RFq777Tz+wTcKOHKOMjUZQZyd6g1dri9qri8L74UJMk7HM3sYCu5
C/XMXF6+5yLxwJ2Ayf8hb0sQ9xwk+JjzpouhKJdsaDMwOQbRR6QROa7I8IJOwGSv
5X3F565q/91XnzymV6FZrkDgUYSUErHp2nqPyqxsqWHInMX46WBiCJLOjcgZ0OCO
xCW1fDnLzz31MF0naQ+GWM/EKqgoL5So5CiO7fPhv/e4JOkCWQi87zfan8iG7WHS
oWq9WHjdvN20yPXAsCMq8JL15mFJolxHKoN/NVKvLOFrcBqPHV06aqkfSp01PLSd
xSEQqQp96VpT1E26RVkWs8U8Pfxv8JExqG0m6DXU+deSp/Cvl+zsUmIEieR7Tmuv
JvnNKqEcArCO8tyyRRWlGBw3gv1nRkWS96PWL/xM3yDdXmkdaCXUzCcaDrOxQvYR
plVjlt/tTUb9A77Sgd8jxGoWMMmvNr49MdlYJEZecKrpiu7/L2IYMgr87tAx0kYW
alt11zdEB+wRgkQHbGZGkGBRnlTztYrRnN+dY7KX5AjN9CXEYcl6O8t06EHnxaL0
jrcInzb4olwptapF1g8CYMCBuq6kZKTTmfsr66CcYQQ9dOT7jioxU0TgPplPWOyY
tH3Z28EpgcvSN8KmrsDPDxKtkrUiFcc/kbgFivm0zJo8O6P1CHTZ8im82X2DXHjK
ocgCDofz1dqJzDlyPXbZyjK7uT81OgUNqkQNHmTSfKbq9jN6VcHVHpGLGyEnenXt
aOj8wXzh4VsaO4wkGK1a7AOk0dwRYQ8IE8hubMbAGwWYDCji9T9ThIlcEuyCpejU
vuCRmjYF0SK0rBc9GVhvJbB87R2p5Jv7/FbSqCB+0ETYktzpWWp0F57WYHqfldXz
rcEMft3V6ZEzL2QkIZe5IV+PW3wl91Jb5Sa7vlGTQNe73s7WjB4DaoWVl2MgSeq2
B7MpmX5r3Fz3QrBiDncZERBZ6gNuLG07YGI4Ltn1QjIBPMG0AbJuq6KyUbFW+JGG
VlaSFfnPLg2JCTaKt017GsQTlfsBPMATOgj+rH3MewR5CDAibeB1kXyz50a5ff/D
7S7TaL0f+mFCT3WIyVgBPXfbUk8ncPyrWANTVynnAh04h7pWv2wehdqEY9FzOBXb
vCCxB4mxmS6yfZM6a6y48AIWagWKdrIehtw7o7ntkYZUFUyFlAr5dD+Iil7JyoWd
xN9FlYRV28alpaFg03G1U+6bTkcK2cK8bPbqk+iYJK5GXVk82309squyYb3JNBKe
e+ChgCCqdydL3wGWO74+TikI1e06mDMcHtw/kiNbonbX0N3n5YUbCQMhxIzUCOgG
PVgonZfKmHAPhVkfpsJMFTdwK7BMBrkSpGM/4xMypNFcf4AYWZHsnXfX6zgJ2Ktf
owQRNUcNJmSXczh4CA+sKvnrVdfQ6GckDSqamaj62ykFAzafWwbn6wNDrNi8RMzM
P4mvKTFl/9L4/giu82Z191OD88X9AVTgre4nikaJVfqe9g9Y/PTij//PhdBthYk9
OX17/DMx+f3hNLhpLJD/zBXeA9/LkHkxSashNR2XKbJfJlSSMrEAs/BYcoa3RtMT
qWiaIYrHs6MDrWoSbREOvviVwAhcVjp9QQ+Ik1v6L+NOJjEnMkVPEDvYbtM3OlNO
PiOa4FQwgOHFFFkdkstMUbRdrUnek/d7SslkOZ6a6SteRIiYBWV6nZrnDfBMX8VN
exbxz7crAm8lyPo7uM/5Cjj8iLPKr/NJB5zGcUn62OkfahMECg8xGQ92PtJBcrIC
EZnTVcf5M6LMTKfjx+1my+3leZMFsSUTBpySS7BQJ0Q2qex7jTl13SYYx/W2xI/x
TvTt8UHU6208A8rUBR08ZESJqqJJ4uf6EDFIGc5891No4cpr5t01xv5Pt0bjwz1J
E9yDD427TH/N4HQyqnAebwW4vZmaFP/I3is6aVw3F/GUM+UEj4SjtsSvg9Ay2kTR
2VN9aCyZqH3izjhLZUBhwulNk6KfeETIFAIGTkhJJXJmrt2gopaPfXduECAD3Wz/
rNjbkt9bBW57kTccOUhp+UsjMuc5L/CoPPWk+ROot35xDpzVZ1vVKTMD+tg77eIC
+0I9L6J3IK9cumV5yn+6caKWIIvLlroJekrCsVsIhymoQe/CxSyJ9IxBaw+otzu8
qdUnejkbqf34AyfuqNilitVdaxCUfT6SJ5fXQ5MIML5i9+0gxII9zBYFkOD42ymq
kw44sLcjkjllU2UE3eUoQeqEMuvfTe5BGG9e6snVHDhZyEBboff5uVJZD8SE4/Fj
f5tcOKSeR2AYB8wqK7fCUmZZ3JIAKvXy50YUsgMZH0Wo2GYDlzmBnB5jHoevyZAr
yDwQyxwi1TstkIpEYRDwou/oyHmU521Au1bw2PAgWLn8vGP5/FCyhnkMlFoWN4zW
IrkKjmVQA69YxUbYVgbcHAP5A2Mji3sI7gJgclNR/3LzxCyJgbTVREAGYPQDqsjp
iQFGvE417ux6FMAqU4woixXGevZg50MENN8Zt2G7LowelOw212GciorNv3DZ9+fN
ozz/lR/+g16P5UDvH6PkX4Io7d+hpUhaHtn0RMVpdaGNMRaRNDVdmex55fPDtlAS
AYUl04I0QmdAEbtTHqbuV+nM7IDLuui2hGIwOpru0dO1RNql/GGSYPrZu+dp4XZr
fHeKKFbZ87PyyBWh9IKsMrEiIj+ZrCeUVk01vUV6wIIdAjttyIGux3Q0HYnUe1Qi
iuyBPfIXxRpzn8Uu8fv/HMTN5IPlEt285M7zsPCKWAg0y+hAoUQ0eELL9Cinozum
/fm9EgL1ltflbprx/CUAZNqI80IOPvJdevu/GAwn+7AvS32MdkqJ3Roq84xq4tYv
iKr7B0hBQTckUjcVkgD+Ct2WZF2ASjSW7u9CGLF4orPPQp3WNX5j3Q7LrtzRrxpk
wA+LUXOp9DQoEd0Jfj+s/BBUCjVSW0GG1NmhOtQa5RQSw18CMLxR81Ccprw+W/KT
lrjwqjCMuMMOD7DcC1Eh1CmQK5okcKhgl5eyubR4Uqk6rcA259wc7mIaX75y73Oy
7WT9tv1f9Pg2/ma7aZW0iB9MdFHB3t06XH0dIA5qiGdOKPWH5503IdO9AIIFg2pb
E0OX3TiknnzvNii97QQkOBAQLek1HKH4g0eEoCziNizBXXrZKFIRKX+wTP5DetYn
4C/7N7BdNMz4akZen0JQv938K2GVuven9R/WOBIKptx8p7mcsXGTU36ZHVfrJL0Y
LQ2qIgvxcxXnXhUeBg5QcDMuPotZ4msSZr/9KPsiYbxl9KHovvi0i97M1VagDua7
jo8uV4lmvpj/imvwIS4buFxCUfiGXLf9pgBRusj31R3zatPTfqnjH5zO6Bd2QtJC
BU0NPWAtXUpobYQxygbdiaM81RtSXSrEujtJDauQLIVl6mhHliAIPhnQPm3ylT3Y
qMzmBiXbNq8+9f5azZ2iLqGKsIRe34yV9eRGrVH541vhY/mhhn+7R00c9WuK7s9I
md+9s7LdluoPmsKlaOwd6CAgNXsKmoZAd5jBw+EfCc158kaaDZHre9KTb2ZUhBt8
9A0E7116kFZzePhrOPP9meMa8Y0JrNPEk93fL2zjHkoU+ty42ZZHPS3eY/32HMuM
IhJsDVp9Fdvjdo9HnizUr6lVFB2sXw0rN/EW40WF0ljpmdxx19GeSlDAaOqTTq/S
LIAlLdeH0FBPvd28yaisjiwqG8U6JSAZvNu49Q5ZJuCLdpBcMgYuKzwMkUkgHea+
++6aj0y8OagfpShLD9w3fV1K5zl+QqXdWjIhxdpwzvdNilyo37ogkmPEcVwK7BcT
uWNNl0mADbz/G0Geb0zNDuN49v7VNK/kqmDnkmC7wDWixUvEIzh2kze6qtckBZqe
bvCy+OeN4X7sYQkTbiBUsVDvb/R1ksVnGt0tWSVEQB+9W7Y2Ja3Hc/+vS/2FrCv7
LZ0mBtK15vdCoOXRXhU/Mf2ogqSHS3Csf3cB9NfKHjNZd4ZMAY2m5/e14VisuRoG
UfA66ZQBIWVWY3Ex3sNQepzvsd9TrK811LvNtCZO6FTG0FBY6/pzEtKa9IVhWPf6
dHQqM42XNqUeXdD0c/3jyRvBGT2ulNQhB3MHEpBlAZJZn6YKq5GM+UBCMk+2E1XO
+kM0lzplLi60Qqmas9+JiHxKYZlZyYvECCFT9ctvjxhA6/AXRhpk+J4d8mWeIt+4
KDTD870PWpQ6cdJsmhQ3m3EJmPohj7W1eopXaaelHDlFDXWS1N8Q7wJqVyb9fwSN
Fkf7ymeIxnL/h/C0cCeozRFqXRStUQM1kVP8F4kUXTyvBxK3w1FPay23LCxD42oP
T3nNjSxrP2K3JvboWwyNxUhhCfdiEQvAudmtFT4dp+mIXgkQ9hvcznL3GfNDwPNf
EU5fn7DrRoqCS1YLbiros8auZgJWjInjLMY7uViKtITKx3eDtS/ejnQsT1itTH2Q
TyHbCXTQcViV+fgYJwY9LIvvb5eD7VvVDOAOCf/h7qmNBBw3fXAwkDl5sWvAZTmV
v+s/F2j15tcmQS20lOCKkFwIcp3urwtNcMxq7qnRScTThqfZ9gtqNVQ4MS8VHZTp
gOvI1lUrvgvTEtz6/qt+fcjU4Zsojqk7a/vJF3DAjdJTHpaWTlBr7YpjXr8IA+wV
IekJO6hhhW5Z3s/FC2caEUKjfI0rYU8TtOTMQqWavGXwZP2iwZXKCpxXz7BkC8lS
KCiUxR6Q5rkfrapiMdlrGN9HSYIHqwcBfACwpMVQfowrcaDYHFB5NVJTN0koGd1b
fOAl6yYPuRTPyeNqeLywkZ9DlDK+kkjWKGCuUN3B1Gs0/+l7WfY8GFhIwfVhF6hc
kV7WicMkeYITerx77cMwsJ0EEjxw88MCnxhmcjdUlveP9Jn0aktCg7aPCD88dbT+
s2pSMYtjkwb+6894+nlI6RvoEW+vtxZ7Ewnxk3dHjEZrb1Nt3Dj8qUPL2Xds9erR
66lSh/rcpq16p4yJjiC0CutEYgCd2AevDVHzTPm5y1SurKVpgqMGe0QK/NjHJXBI
ZLuSbR+f1HaI8fawHXnpJZUJDZ8JQkYVm383D0lIP0ggGr1I5jncG0qvurgBwHRk
JveTMQNKpH/awUh39udcbmzpA6vP7JkqB3stDYkwVdRN3zqICO0kyHN/47Bn/51H
9k/54iMllgplwhbCFHFX4NQUtzXbpWINqSWCJ1na5TIaYPs8LCJ6tfBfBSbpjSJN
eo5pWnnJAUuj5atKxqvORdOId/eQgl1lkr6HtBFtrOIMiVNepZQ0aOB3GyLSRabi
q+Jg47hF2UNGJmpAALkdhHKSEhfQNIe8yvr6K0+Xo1QnooeOi5Gcvzimfq419kjl
j7uXeS2QEsAqQYfnscqd4/LWMmEfGJKAWz0T5I4XW+B7xjyTxW60EfGE+Xcr3Cn+
0uQQ+xLX+WkZWsm7sgz/YBXFOkiAEwaWvTPf1wh3+ShvNLdvhI/8YqdHqZ4tdWR1
aOIEN3GKU1Vy5FixTU7x88VCl2PTivYRN+b0Jo3aXpXDzl3h8rXKaZMq9an1Gvv7
ZzbOnVerPFljn9T4q0pbl7DqEmKkt/NIlV6F3jR3SjPnkMiqZfJY3a98VQvExtnX
ZQwh1VMtBn/qaKhkaoRjbvFxyyzrgceijbCmd+/QDcmSUXHBVnTzJZNPPmI3rRls
8+hAo6qG0XNQ08qq4y5pFkeb5zGK5sVBh/aX0VY3AEAQCFUeBFbw3L9tNgWpLLUo
+lzHIiq5/Bp3uzPDNfCrLi34tkxcM9ah7o0324cSvra5DGNgUWDnbPJbDJs+RqLQ
V57ewT4KbTvk/YXb9cdEAANY9zDJy4gSQgr1dPzZKT/RlKXGevOpPNipycuVqqSF
+h2TB4HSd1Z3hdHXOSC83b7ZZ5BEWReC6XAnzhcROpYaR0KvVNbGyIjveQ6lvJTI
3dYOM/87osU3ZkvYS7GYtl7z3/pZ7I2g5WcXeOBqeDgJV0QkgLqAyl2MaZtskQH4
ER7J+GdczSc0XcLdK3wQ0IN+UnXT2J6AoOv8+JskBXb3q0bFuKq7/kY+N72LTJsB
Ye+VJ2Sz1lTxI4wa09LE3HsWlQRJX+Qyh99vPesypub3hyBmmyDjmU3Z4hyszBzv
7xOuzDNkXemFJbfD7CmK15GfqyUzO6LmGqhhexam6u/rcJ4bt/CwuImvyZ2Z/iMn
qRyiKEtV/cUErkHYzhw6iQV3ZvTvtmYCQ1f9NsbgXeHh3tWsS7cwELxBCCoC+RRc
InCplEqGeJIpbQqw6HmoHgc7aU3nwaRtGuX1Mla6nyaHeokKiElWriz/AocGyc/2
pyrLVa56BW98KN87LGdPKg2nwFDjlSvtQg575YQJVBBfmZ7RiTazV2mUaKCdXyhA
ju2awG29w071ZZYxr+iHJoXQvgqYqoQQPFmXJZ6+nDMmTADfSObssjTBAopZBRQI
/frabLN2+aXDPBRLmZQtNlRthOs5ZjG1TmKs0ZvrcK+qO1ilcXbO17sEiqWAsrS8
Qze0+LDyVYLLrSoDb3NPkXFTfm3Cf065qtVR9vVyuWUKMpAMCZ9qxrO6Fcjzr5BD
B1zBoFVJHqSzOQ2RCijohq3IVbtqcruCe43iIap/Het978yNVTaAnKLdzZPB/Rez
93BarfYNlDkFrBgdQgP1dg9o8CawKjMnc1dLYfk6QHDg2pnEu8UbIg+ESiq5Pjlj
Wt10O6tsndoO67ZObW+OSA4Lrz5nRjtdZLb5yN3mXJoBweqFqBgzSWiiaPnyMqEx
bMSob0cgfCZZPggb5+Xk6Uu6/n+PiAt24c9miuENZPqErFFNYCh0iw34k6Meb9Z5
PbHXcNytdvwyN1St9Bkecd/ZmLudwZFkaswv5y6WVuAjDgNZZ7H05oZTU0I+3HJC
p0VQpl2pleAy/vGCGpWmTdhiebgJS0SR8Uz6x43ryvqBiHgwqcvEG2aMyL3Xil19
M7U4vdPMXlW2c1/Z8f3IWr+4lwO1z6N8uf9DtfCUgcvoUguACkxdxke6vDqNc8uL
yHoWGv1w0anGKMI00aAgTBREHPXjL8SqnQohbPt/6YHk7CZdH7OakB//W+zjP4+0
FizjVk0B0USMVwz0wgZJrL4dNERVPq+hc4XVa/pUc5+vIPpDQKI+C78j8DK6DPYl
eLNCAapsMh+cmp7uOmcfewPBrrb7j/esMMMorAdZVXMYDiaX1iwMeS6U/R+Y7uZC
r+cCrIssZSBkceUeEwJ7PFKTVJazNuYJCDpQfxOYz5O1DEA28FQmLrH9lq/5qNs0
gjFWKkNSyGc9ed+4Xdj9+9318R9mezGe/tuNxGN6T0BXn3J+q4BWtTlEh8AxE1Xy
RuQ3GTSXigqqr0nkTxj6LB7fET+xF97n7LCOtHBFoZa2zCN2/HtvDAm6VMF6WMXR
vb5FEQ/dSwIZTos/PeSWTQ7sMTB3IFFA1xL4yacqwIluokjDrdCB/okJ4CqzTmnH
VqgPCshonyjiQw56LMV/khubF4b0l7r0LZg8DUF5VuHCFSiz3jND9erIwnuA/Xbx
tIQOHfL6veBGC/oGxb++vs+kd5HvmaERAW/NA5eA+nJRacMajfT6aAfCiPDjwndY
7jJNwNdQC6SkXkzuuZ/DRg29JDcM9UENIL0Wl9/HTotS3+NJGRH8FdH2tHtosnhU
a2B0FTNVQIZhctA+OnJ/HT3fDEjQc6e+CUjmvdp5L84Hbx8acHzzIjMi1BK/6Y67
l/+lye+JVfS9ddt9mjEOxUJx1yZu8XczXZV3WnPfLeacZGyn8sT9rxCVCRtpOWdR
0QxKmmEzw6CVts9EkhRxTApt7Y3Ro5EPWHBmd8gzu9IxEOASquMz6hQXFKGxzizD
0JQ8vs8VQ48Ziwtz6zmbxvQG2AbayFNldeHhJgx1WSvSJT4Z+TBWSLqbG9fDdhqr
G4WPRNvG7HMktZy5xhKFyjSKsuhLMHS09VyMW1SB5Ib134ma88lqkS31RB1HVj6a
twvLQNYxunR8hUFEnlY1EnX8hDlvQBop+GzI+N/EKAO0r7Q+xZQFNeOAHl4m8XyZ
4CRmxy8KaF5z/s/SYsGfwGcGVOOrz4LxNrjd8+VQT035yTuOsawUNMsRsJydxkgR
mwA3t/ExfWmWxpxCp3Yhg5LA3WO0m469oLEBQptuhmHB9xlCX3TTh7MDJH5fwC+6
WKv8z8xUcDlKyYBMq1jvbJ6FflxHHKeigUG7NllgPafB4Fk9q4K/P+KnDggjXwo3
dWQQOdrLoPkS3aEDp8unopMN5dx7t6UiorLwusHg66PDhCnJ/VLF1KEUb0pW+Tse
FHSoLwGa4dnlkGJJZoQP2iUoQ6YO6Fll7Z4bk9XDHsyNltwwAAEaKhq235k1wnnh
e8yFsWNP5C3mXOGBjI7zNZCBJI92+cAuWY1OsjfdpStLjpdNlAFrLz4MGLO0OrxH
hMsypeu+vwIaMBAgCkCnvJ0o5r+K0bYy8WYCI7Kr+utdJ2PgnTJUViyquZny8gBH
S71DuNtSQV8TuwhvdCuSrN2R/jIyjKt4lIBGorJgFT0O9ZMyg95cDihNl4fnMwku
qUylf0JUAoUJZ2vHJqeSFJtipCWCxFXoJDE/sZTLeBMzYg+QelxAbiB08oeL3uZ+
PD/Wy7aKZAalpEa6OBbQz9aaGFovsqJ6k0i3Kte+4WxY+psRuqLDhaLZ4IGa94LT
894TDHPnEkQYYpnd0U94yEuONKrmKwDumgpxJEY5NJuS6wJmkPJ1avomgqq7s0WB
5adtKSH5AVrUUQ/Pqr2AWvKRkiZ56Dsg255Ta4Gtha2dNDNwkpl6phg4cBRtp5Os
Vvv9r2eFYLyYhgMMKU52YRhfH1TZO1Zvc6ZSHF64zZXr62CpII0l/itv8RjS/ndV
WI7LODO5I6tF2uhTbX1ttlVIW7brNr7aZjbyLBgtimmNexH5xQDiejpRq9XWfIPu
rPi3x7kN/ZL4/Cjw+myupxCBgEVzPsZNfIvT44VlZJOoQOHuawugznZBMTVTea7a
AELO4wRJZUC59s0F9CnCOXGs8bNrfvjqtS9DtrgEnkjNXo1ua6BZhW45/QzNx6bN
q1sh2ys0ETuLSuBP7yzf9/kb01V35o0hro34dBFGWEnbC1VtPxJB/U2ZqpSBhPJ/
p/Psq7DeYm69Tk3yZ3/WPRZ5H0/kueXepLXOIB2c/M00vntU+mJjXQ+KbuIM2qJD
6LRMZLtsKAREfHZ9XEuQdkXmrkZ5ZGWZo0acLjUYFjx1StyYsqrRtzhdWOnG/+1Q
mA/tusYjJAJZENSZFRQ01rC73odL0A7vXHCDX0M41mT/Q7KvtqF1pygNLvz63vK5
0BFuiRqLuOdilv2TyXuqh5/iD5SA539vnQNkyAbRiLNXayNiOrfQEXbHN9kvOfi+
oPzww1V94dzD7T9cUGl2buJwOQLiTep1e2qjvEXUcQP7YrEZ+3OyYHZWaDkAwJ0e
uXaIDX9BEc4YddVhVJYLkmbwGgp2HU07Wry4pYryjuqilO1+W23LkZYy8d+MEqOm
KVgVYtPDuSwLcZ6M0kyzPTso7QVgwrluN7Umdu8lA9xbJAHSnaJnobjJfc4G20Qt
Dp4GiGVrJ5P1ffOJhaNijJJQUOjXkdlRV32Vzqsp/D5ua1O7voVSWaiK8sl+sLHM
GmkOMvSqXUO6XRo9hTMsoqVLg0DgXH7k+Ea3tmhImSZztnGzLGsPBsU1gUwyB52c
4BPZTliMWgyvLNQqsB0XH62448R1U43KWH3ib3UEu9rkvNg8ebcOssTg1HiO9DLq
hQik6ARYhSb4B4FR4w1Wcipsl8prJcWiHHZ21JEgBPm8JQKv68ZiEjuodlIN/WJ9
R4F0jza/6wBNX43VEkLwDgkj0o7IEuhcA8GMwJVA/SBzFmrLtVbYfNy9/pwvuZqs
VL85RqxX+fpPABPTFPhlSTTkOYf0Wbv72UB6p3c+qQxlxN0nrjJJx7eN/VS3hwJa
pCGTwgW+9lILoDaK9ctyL7yJVOl9e3pJLT7ePqC21MA9WPueIDPj6AK6FbUQeWQ4
RaCObpvwcEAEtgtC1snvhZ0sHh7Zi7hZTf88huW1Sh85U6C+ok/m7bjHt6H0tdw8
UQG9qaT24aYSop+9kP0u+ThqXyfzGYK1+lz1QnAnFLPGktlQyXfnoOGPPP5EoC3U
qjLGZRUo3a7M5p0Ckj8yvav9yEaH4vQr6i1uapmM3eiz+Dv/C8Cpw2Ka/QzIvcg7
qcWyE3v6xZkJpHQIBOlZf48Z+1FmnrOJcisfWPqay0c840w4GOIt/BK+UErg8fme
MJMngGV/3W0z0+uv2iw4mCP7JZAocPWq1B/5Elx015k/4rMAGZX1J1Nu3S+N5g9X
PNgAaCvHQshO3AUlMEK7KBj2xuPZ8i4pbQcizA1Ca0lrHDU8XqSKHg6Kd0UtWhvh
SnUTrbuY2/8Z0DiF/c3EIDBe8EwU/E5DPqkiGXK+8jnIcGJ77bTjJHGcfSi9bhoR
JNPADQLY+z66QXafwYoh288szxwMZbJFvB3lfEp+nK/cv/ZIh0Z0U9eQ2IUD+n0F
ZWaua5gW/niLfC0jEZBt4lNJvvViZ0xXyuvWcNKRYLC0NkgJ8tKuFYGzFl3w+1X3
C6BPtyKH0HpWIf8peJzh2/jrxkPel68d7W4h1JrB7QSiq0tO0NbDPQbWgBnfTAcU
XESirofIWoBzuWNOcbmDBjCGYNmwDUlf1eiTdhSmrtWZbNkwP7ZgC9bZZiBhM2X2
6W4DtzGhGAUyZgDJaQz0y0SJq1xpo/2j0Ct6Kn9y/NVmWxnfG+KbmwPjQp/YT1lK
`protect END_PROTECTED
