`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
12905OGikXOlkTRYNZ0z279PcDMpapjEqrAcTcruUuBdyiOj2vW8yclT4UmTIAYa
2ZQE7esPmShO/XeSLpPfRWBEYvFl13E4AyDNFco+IvxGQtkbUdovDErT87amZsYv
/gYjgbHL50XV75MpY6c8l71UVJ3mi2FsWQ8xJjpB85gLcY26ei9Xh4tBDII3Dkx8
j6cK7ipHTT4nN6cQJdflnrx+8sYgXU3yw5YProldu7cO2vhvuw8QQacWvt6FO1HX
SyGq5OeiGJu6cVWBRjJxGnu+7OeJpfLhMZjDjYRsqzE+GDwaKDT7HDSLpi6+pI6m
RZkObdO+iax47U3axdxisCpspzvxfodVo92Y72gPqktdFRnpVQPs8m69ZOji+Cvi
NOYfABS+iqT74htIHSdrnvYaDc/yMQvizpIVhtrJFM2fxN6Bt2ACMNQRMby+RW4a
bxX30DYyRYE1papDPJ9aY9htblHyFpyfUt4YZxKZw0YmyGA3WGTI5Gsv9yScpXJg
cn90aEeaXL9hJOGUvb7qo+1bli9CCvPbXUodNwUSE5O3X+cl4Ir73dbvmfxGiRdZ
ye0KDYQSOfB7ijbQBKXv6n20jr8JslI1O88AtYOe08LqCbYkurD2QfXERDziPqpR
L+i9M6Kq1BPKvJ8TxrEc4RRmGyoX1rRPJ/ztxUOiWPxJW67sRHMNvNJIKmGL7qYI
OF5mcNh2m5fifKI+3WUtj8uX7+ryAJ4fcA8PLHZuAlx2ZiI7tRi+V1Xz+N16aVQe
Rfh3CMz9K0okq0i6h1PVEboB+AnZgr15z/IgR53XAZz31KW9dkahtu7KPoQFufOO
plWcHnymYR8zHU1e6iC+Z+v4QFkR5g9/3bMN6X5eVs5h/NQLC4DYXkXvhPEzgsTT
PDiD+ymuPc7MbPtxehLHHAMFS1wdck1pl+5SaaTgZoiXD9HUEjI9xWmg+BsaoQaN
bVoMWrYAmPtSmZURERJYUlu0i6ZyOS2RLihalOqJxxVn+sdDhYkM9NUkALTXoXie
PexOe5rCFYdRHl7cA8odi/mN0wjy3C4ekxKhcKuvU4RF/NRZH8oSayTUv5pCQewd
7jsLut2He+3RVFuL7pS2DGbmzGHG++H6EKSKl7aMR17vIAG9WapvoWVrs2lEOSpm
IOJmwhukGcxDdaliUlXD0qfo6IHRNiGvXdroMPORANiPuIuNFh9T+PD9/VBMd6Sm
lwkzNSNmvXIpUnVlOgSSY3SehW+5PrjVUKXVpi4GUJ1tPgXkqWOwVIV124lLT4s+
x4Tk6uXxm3LR/VZTocPidfdoldEJFqqlMJPeH/oGG07WzTWTJEIAWmPLVoTBOD8+
okCrlkx5cNU58uKh1Ppyd1+TqursipzVpL8eA5EfLlZPkh4EkiI2nx7VbIdNSpG+
VdOte/53OzKrmi95KhcRjE6gOC/742YCF3v82s3/xIYjHAFjO1crbG9HGrnynVUc
vsHkpVKEsY6FFFN7fi25lUh4JYMaXTdBvRnyFAEa64f9Gi1zpIlhjyhqfnqhbe1D
BhzNZ6QEp0k6kA0IMjTLZYCaEoCwOjHp0YxqflgxXETmhh2M/iHSRcWY8I7wbWA3
KhZxL72KYafJ8ijz2IavAl9meaKlH2Ik2BaP71XDHs8D26lR7AhI+MrperUP2Xu/
Wj+vDnYTSn/O5J/BqwONGew1yGYqZKlpnqkGrKRejMVg27a4gjwq//Su5bpUv/nj
x6+Q0zwlkT+wkURg4DVm1VksO4SfPWMI656PgK9sZLOhL5rPC/XKfcBU+oawCYFI
mFNhbXzv+Npe7xWW3WdA3nodB3WTwXfMMPFaCcVhA1spIC3thwUjk7O89SpGIMiW
rypm5vgaJgln/KeHZsKS9L6OzA0C5z8Ff87eTKvI4+hPpPMtJ/jeN/Nb+kmviuYV
DzZqWKnWB2aHtyZbAzRjxAdqgoDraiqiW9pgnuUirZRIqjhtDr3Px4qWaX/6Jl4/
VTEKMlzM1bfxXH0qegUZEj07VbjBoa7WgQqpTiJDlQSlpjiKa9yUCNSamVBq4btY
SeeUeJ2aiW1SRl3SCPJEHdVCe7sN5dAD7WAw0KFebtpgFkA34ZdAc4Q/sRdAwrVo
sRdp2vrc9ZEbErFGKitXYMIy4W/lmsiw4SPjiUSuM8mYtEKYPHzVECC5MfJe1XU+
1NgM2dHdR3XiFiuDva3hRr9RlGzaCNzXBkaNKM2I11+7krzvrN3vFE97Wl1K2Nov
Ke0nkx45ufJiB5YV7vk8x9n4+NXS1QwmlAorZKLm3pJBhROZasHtdotuBXmld2ec
SozibN9zyUbdq38PHuQZ3mJXEspRfODpfd8hRzK3UFBYpt/nL1p1COMiLd+8MreZ
FgvwW0iv+u4hIn66ky8n4I+wDCkYRfDjUiLoLtzd+9k/axFjFaT2QFuRU1GQxKHW
Z2eEMbToLdHWtETmKzfs6YAy1OqBDh0Ro6RSHenrmHLAhrPoAU0iaVTBLNzk1J+S
Adb5ROTU4czXxn8nmrwaJuGZFiTMUwDr0Gra8tdD9SNCjev01ZyEodZIh8m+MnF5
QuxATeTs8v8CLb2Mte4x3g==
`protect END_PROTECTED
