`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GtbM38804Lf8RuTZrBNDHDDtvd3ApEP2b/7Y2WJTAipHa7cTq2khvxVvy4hgOK1g
WZnIOYSHRFfLHu0gPGMy0/5373OiSHtJQwUduhK3LacYP+IxXIQJ96eEQHmU2tz+
qzQ1COcyYJ6mtqNzO4LM8JfDi4lj7MAP+g4EqdoiDW/qZ23NfXhgJnMq1C6c9EcQ
8vMO0ZMylH7BrAGoylo4pyl9ggJ3IWlM1R/A8Ul/Dh1qUaeThelNtKZ4ofroQDx7
rpnhnd9OQx0vIGlsGWstXFAqU/fasEAvL1EytGlm71kzOGLQrnU5KqWchWhO6v1y
ObNgRbh3C0SC0vYq9rDCtUK1NOQEOpXVAFOYLFxCbbTqPOTHqlcijpuphFps0cl3
OfVeD8QJ0LyVtT0virbrrWtEwfzUiE4GDuFb1Z8tMuIz8Sff2GQ/HvUBemE1fW2r
U3ghCUMvC6OxMJyAIZ3kVjzPM6WXh4r4MZ/cUBLIP8axT1Af8R75QyYWBbR8q/X8
WArCkla2Dd5IXEA8OsG+m9GMSQCnfaS0tFTugeX1vyRoGku2sH/kyfY0JXCOV1BQ
cCPcENVN1zoQgdMocZ9BPunjWy09kYXGqmPmS6kkQscLhA5cxVI3QJig+xxtF0Pk
2o+FTqXhk2p4KuAFGX73JofYZKoih/9jsNh0wmihcvGclOzd7cc4y8889DJ/W5qS
+eOe2qhTq1M9Ch6C6klTaauyXGG6NTEuFLLN79ewS5t/uxHcnrjoUdU+zd9yvKA4
pobi3U+6olB+h4zesg2QjNF78X4H8LqDUlmMfpsp4eovHVqIY6N1fLjHHH9r4lgY
DQbiOVNspMNsCjn68sJfCORT1F+huRA9/p8Wowk+i0q4NFAgTpnWh/rOsoAujnSp
2zbjCoaeewDlFbpyLsdkJkTEPDUsBLlOCuMezvK2JexWRPc9ETgQWSlurJT+Hus1
1vGtTiTBLJT72JGEWDiJ8jU074gcbIVo96T5rOn/gZRFLIcKJK+qMAwzfhfOT6N+
bShzEyH+D5v7ICr2ENrh7O10sXsPg2BwL0s4Adxh4/ixEr9MxZALv9ZcglbMz9v8
b1UHZJRp2GMS+7Ryv+vRrCXEGmawt7f6t0waIpAxcNjcvBJKKx1fSsLm+RdH/a0t
9qQAQwgcfnS1q4O40ZOwyofNpIcZmp6LEKRhDG5zXbK880ixOoHGa5t5Pa+0klXJ
+9npdBYla8fc2KbvgYfZff2CAFFQ7GNaURriPsirpsV+Fm4SnX1l1Xf0/tY0cYnx
V1iWZWA8yXhpII2KGGr4xyuUsPSHh7GHeJNQwOjzyzJCPm3oQrfx5sr0HWRuc1lM
Im8Wu8VPZoGGU583PsikPBtkTwkwdClcxCv+T1fTRxUOP+OJN2bZRKFdTk7cWYkV
hly3eZky1iTHT9oDDLrOskK1eeKCOY0VDs2+okjwpCcqnHq4hfR3Iq4j06vI75mU
dnuwscQsUOxoi7ygOSQn+PCRm0TlHQHIvqW344FwggFljeF/tCa8TgspHtk5COdx
QrGJSY1ewLPPAvDiF4hahckAgpX6o46Oms+peLg8TqCK8aeT39UdV+LgDR6X2U/I
yNsTA3XGGPKnC4LC99kk26kfJFUDJnlkRIUhSTozs78txR4FGZxLA2bo1iwJ6EbZ
de6td6DXJQzsUyWlO8xkfyEu8U100jnlvUhpzaVg3Yd5vL/WThA4/7TVmTUavFzW
+F91pvAEKOg0wnpqK9Bx9Dt4Ta4+aRyLB+vE4uxQsQIEWVsokuO5rieaW2V5eHZ/
HI8FRDQv9eSOiA3pr6s7pi0Z46QNj1pFNy3eoZSzEsbNMK/GN1y4jZnj210LTKe8
4YL2RsWQcCEytElnMpfmmS63BSSQA/xU/6xrz7u6MVUEapTGDIsQPA4x3EE21lKP
+uXdRV8siECveotjJn/8c4nx8wJK228dkIrGiYhxTAL7NUwqOR4gsG9JhsbD/PE5
AknYNOumPbV0Iqszwun18cTRSCGmNIyNX2DdFlHgMy+ljP6LN1q3dZavEavi8br3
JlHluJ03SY0RGmvaniHAZ6kI7UM74dcioUmqiSv6sJGtb+52jpE3E02gTjlI7FXF
3S8IInzcj03+E4+Ans3SAyf7+axxelPcMj1caOE/8igDIa4RHRrz4YwulPC2wN2o
8g49YHc40v7/xJUCP5dWFfQxg1kw47eE0PaIWYmSC6lhn+/xxgKWM4SCuLEUKwPk
xBI75eSlK8uBhHjdWH8dOYsw6fA8RMB0DGFYF4PXPHdhVu641AsjxWedUY4fmp4g
dmg9PRn+wDS32vk+j/e0RQ91PhMJ71KqyF7Hgh6TqdE9F3CAz31NILgYexp+Jk52
wzzock/qIHoQFk9tZwJOYHRz1ERqiDdsQPcQcpFSmttNdT3Wnwn6kHJm2OcGqFb0
rAfJzJV7ldjN9H9gIp7mm3X1yUc4yK/p72jLoygIJOH2R83zWvvhiWL5CfkPiKkA
D+BWt8ivpDI1OnmWWZdTdJdQyRQqIwjdbuiHxfCHATsyGRxJ+Sp1qTu0DOwfDxl+
BG4MFXgXnIFCxQP4YNi2ToXIDj/ujnf4wdcHTel8gfRwl7JuhR5Hszvi8nouFtO0
c6eXaZvFPQXGAq5UwBpmQfmX7i9vx3N0J1rmQmLbWWLbCEGHZYD+rtWUWZ7RSjaX
iEOEMy433YInXkE698GPdj6BxlVvlWVzW1hfAHDNCtYlmqVUpa88jQlZnYs1Qu7c
0K0nWkvSL92QwUCXfhfTFhDMI37cfaq1AUGvSuOYBMcxywf8of1vl8LlUfl5T0rs
m+E9LyIQDq88kMW3GKXeVJyYfAipPqEa2Ujex7gTh+RXMGi+DRnASf6jJdW1Thim
sRl8ZZQ3fL5dbCshoH/Yh5riSXsvtdgN+LJn6Ae0+FbqX64ZJoNboVfrGkhK9Fyc
Mdxl8YX2kSzTrL3rVP28UHfU2QG2IqPA9xZFBb1I6kGqwgztFrE5M+/7c3OFtBx/
IdlxApiSOVHtJ50gbM4bBRINm4DxHcyQVSbqQAKKtFE2QLOzKgMWRcEdKPd/6Ftq
vNwmCtYsEJT3qqu3GzOekGFlm/Z5tkNrRlNxSA7HGk08GiAS1h8YMF6QqWUl80eD
G4asy7k3LNB6z3DltDjzS1fBOKZbCTZ6hsH/HvXWqci6/qTz62BYLy+N7Ea37BNx
XEOEblTP7CzA5QxoLNtX3JezEoOUQDl2kq9a617g+/buD2CD7CtTfcwk2iuEPfYH
BhXyvD6ypvzv3cIBCuraqL5ooIX47Nod+eXWfxmuIS38wM28QmoEUzOktXg/ndpv
aC1iE9c5lHk2lEhXydAfboTF+x6vIAQYZ69nQC3L1FtJhdyXiLKTmAtIhZBIyiZ8
ybxyc1Yx24AKdF4FwzXpdVZPU4AHTwLe6u1xeTrAinbqeC2VsVj62igho2r7APPj
t+1TGb3ixadJ0cFvxovoA1rlO6WSqeGUX5Bt2KHBCKnhUgIYmleVt5SJDmHfWgj+
8j+SH7+BoDQhzBHUwLNIoiTEBZop1lwqNRzyaSXytfr8OkOhfzSFhE01PlbW6/92
qwEr0E39QVHbr0JJG58IuS5vrjD/38qV/jw1iSxjlgRPPa7hepEJ0XGGD2BjMsZX
21iLFOKP62XPOJ2t7csg3LRq1PKhB9m8lfjJVVTWGrCdyMAyVYlRj0XYgK7WbFyz
IHjpzC+MUbLOQGNEDqboElkqKaSqv702zVNDD6cnXevCqsOSP6iLZDTuMiHLTW7d
zNnSquwlwQ2v0JOpTL/wMzk0LqcJ/Cx464XMKTcAMU8j+oMYgz0/6Ie2sDHV0HQ8
pTG1adXi7i2cuFwSGqY2jwa99tkA4W2+oOq3cz7EKZ1MoZnxM2AJEWScKGXcgPfG
qC2l1aC9u0F/XISJvRizmmNlAonxQa6BM4ecvwLJVgsjEZmBcc+LnBClIM7IzPkz
teFq3okWGspM/forfw9anMeu+GdsoAMgQ387RjQL+sQ4oAzRRIqbe35zcI4Bqbew
ErjxSU7z9WfEhKanttw9gdUO+FwexlG4gj7ovIJVq2cy6B5kI2R0OOEmbhu4qI/N
jZe2PC8sRzd5Maz5wFKd7kilQnerpGDETXmOH3JlU/loOnsdnAfaodEUd5DSy+rd
4UegMqz0Pjvb0bTpCwhvnYJnVNlsf+QIb5Y6bwzjiW50C/Dp/i9w8LjSkPKQ7Ltx
3D1Cw1fv2ictCWSMQ2AnR2rktVbghlpR/2acJZKVM0Vw7mLNwJzL8JNJvJtkl27Z
GPBDNsU5R7UgtS2LNZN0mA1GCcEkCYJGsxWC6Lw1ywmsX0I4ndIsTdqG/G/rbxWp
AHaR50Qe+2+v26cfOlK0YZLim90IFeUE9+e3B2BMeeEUGS1+CjHhBwjvabTg0MhC
KNXC/Cr/1WPWbZ0QPqrvRSQx1Pl4OHPbdT8CGRCLoj6sdvJ2wq+IGOgehO03LYb8
`protect END_PROTECTED
