`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9faoFQ6MuurXTGNzhFKfc58dv5N2IEJzd2mM3Fj4sBzgzhYhXZ2xfNjAt39IzxrW
0H8OsAQ1qAfGXVJWnPs2NAPA0X9rh30uMAPHCciXgoJpa+xYDWfVkrJZtKq9qkQY
EWt79OX/7REz8B0WyejrMgq75CkMcr5aX47dokTC8jBs40fB8tyy5WGQ6R1CFYYC
lhyUgOTPipfSwG4NNqjZV7qtqB4GIBAAdazlCp+wg1Bpe2053q6HYb6UdC9262O0
BKnoJpCSHCUNiSOR3qjfg81aDAZbIOIUeXlIX++ExN6t45RCPh0QzC74PzKYlDuX
ljuSClt7ZnCHDyLKTNq+UmN5sRhTPtCXPu3/pRPBF3UCCwAjrGyDCmUdcTCrkW6e
Hs/kXbv0M+0U1OiT4Pze9weMd5ZTNAhH4jVpCULz8popLoiCJGv2PNEeW9PyRlQB
xpOFBmZQCGrhKc9ntZjiiAOIDLSz5cbX+BhCnKMiS7ewhnEB/UJcee8BiSDiEN8l
l1DjAkO3JZTKFFSMv/3PQPssJke0/F4YS7to/iAiuX4VRWT21pcE7gS+xT4nv5oy
EdA2TK+MipHOxd/lpMNUkDL/6b81TgQFdQf07sQ7EyjMGKdW2r/JL0mXVpl2JNAN
FdaKaEP1poRHi1sAIBYwhm2K+je1YO5ZEBPkKHirtrPZ2biHJ0hQjcioYrRz7SLY
zeKYQolWhGrZJg7MuI1ErLs/sDGXOaB3KGiJ8Oj0PkxNcQzGnSpbYihPrPw7puQ9
HcbtXZoLp0viQP2h4saK3+sWPxjZMXAUcP33npsFhGvVe6D1D2oTV46oPyYkXgp6
t+0N0E8LUvXsTfUzEAPF7R5V8kEJhuH6oHDYVfxmQ8vW/FM7b1cXxXybCDK0C7w4
`protect END_PROTECTED
