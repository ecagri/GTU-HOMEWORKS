`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XNixaD5IpWPLe6Ntyem2eSdsZ4dv4SG5yzoaenl2ktqk9jcFDK2DqvgafLy2SsGw
EuHUAKVKJ2N3kN3Ln9FA6Qj74aa9J5dv7GnOnsEpfn/E2LV7P6T6yfI8tXgSAi+0
IxdibtS+PLjGcvejHJ9UOK0wInklKSnBNzOVZyAgkonf+qi0lX/lSM9riTA1wU3F
+b5Yzg0snMAGGwVrWa8RrSOZGfboyzatr3I6JP6qOfixW9amscxA0Ut8olQZ7a+D
wvrKfT6q34p8Hm1NVoOATcJB53QXkGMhjfciRitkw6h8ta2cxfxXTKPmzYTJrQ3O
vfiPu5XBGmqJ+3YRxBiY+uW4KfGWz/xLhFlGIgfpdwfVhAqi8Veka1SwQdlsI1v8
mGn5OOfxIeS5RKeELQpNvWghweyIDBdMslRU5ud26bLmh1kEwa9KcrODl8T39DKy
dJu2dAE/79VusoXpLIFKfw+zMxQ/7me58Lki/AdAhOjXzYTB1dqqxKY0BF+AbC4n
uhh+7PIOqmewd8U6UAPWO0WDPitI1O0RxGW29jIqpZTouWPRPVL6BqC6orTwS0W+
ZSzCpKH9Clbu195Wrto1hsHmYwlaL/uEnvlnezu5r2AVkJuRDLC1I+iLo2WQKh/r
pj8kplXaJjPEeiyy9Pf+HiJ9iYF4p4RnFQlyeHAs3wd/2G7CGRLeJTwe2kqazZVd
7DSWTDpZYo0yoCAIgLI1rPD+wta/XYSse3nTmDnMQSbo4hKNThTbhlDhckn9+5hQ
vNmmCIrHqyPCUQCCNBu0pcSE788CJl2sZaqNzvkoQ074UGyzRU49QvfxTcn2HmQ7
OGa0YbEeF9m+5yJoj9qGT5Kg3152D484nX7AHfDAFzbw9zAMcXrZZgPlAt/kpaf+
1gaIV67GJHY/fBNfC2wnsgtStTrICj00nvQ1Y1oMKQIbLVqqIhhz8DYZAQgv+rcQ
HP9+gmML0pLeBZyMaOscPrsdPdn8hBn1Plz9erndcmL/Nc4KDkMxbuqYtbppYFSu
c20SugJxBH2r1+DlAVes2KsFI4P77mNTR449xADJlPtbTwzaGOYUKIauIVAIjBxD
2Tx9FUnJy0ct9Ii7uFJMQqDGQfwwTxc93m1KAjKzQxtxf7E8GhIL4Quj7HkDgic7
UWnLlzjat50Qm0vDmLr2TUNxD581c6UEbnvz5ReKBV34Id74PQqhFToAdAMjDPXY
OoSPN0oOKSJ8JuUdYvPG3aumRhFMrKZjoARkKfkGomLiB1N51YNMUhjj5lEiwOkE
PrEEyuWx1afRzRYnvPblAp+rHLTw8WEGlCc+GtNiEAOtjFz+HKSecqKhDDz6f9ZK
uFw0szhWrOfqrTPiGFPNWEEl0GCwEjiu1+37/2aNEbX2Y2tsOQ0BuiMIWqnEnx2L
wsWNSRD3twv2EYzSnT1l4mmiX0qzsuvuDwaVk+Gpxm1aQMyPGAJWgTt43NBk0/gW
gZl2AB295HQAbFru+fXXTy2/1swWWzObPiefwJnjMmXOT0IzGhSKuVaVH7VOYuS8
Few4nFc8c93F7tNk98qva7dmshgt6GnElDmVzlRd7Lc6mNCLCiUadgcxRxhWMCNo
lPdgFiqPEbuecHLpcCkto53WvpNB9XJHLdizABMUinqZOcEtsV6MAB7cXOkjWhUx
EyMqkRS5ZUni1ZsQ0xnJ/qEtbgyp8ovpGm3qjAIz7ypDW0MmTojDBOYIk0xvQoP/
iCEbEfCzmnkYRqRcZuQcLvHDQ23FANb+qNw5WFL3JyXVltuNuu9ch957/VN4P4B4
H6I2MyY717i076yy4l1pkuR//3NUlwurUj6eIFFTUk/l9iZC0pMp+qTTJBAAx7P3
libf/KwrVqXC2YsRJ7IQFfDRw4Ed+K/a3jrVMmoNMlhImADBeVB4+8JoT1mPh+OG
fKDEFz2cYewZAdYD3JQKrwmTff+de+T4T/3dNvD4GF3Qx608GcoB5dVzsQbbhK+Z
SqATBFw9eXoTBPUng+DwG+4s9ZUY8MTOdv9uGoAD6ASnxJ94JNSP5K3K7N+4Ghj7
OnoWWfJ5IODfGDbpjHNvMM3pZWwn+Aink5kX9DJQnybn76zgM/LNJBWJ6W9HD+uF
g16rCDadkYLUN26Z0SkyBtzpSIhEoeG9rG4JEqB77FDAPX4PCdQcDzxBzEz6Ok8u
N8kpxVLxtmo24Om+HVzREvgRD/+M81uN1s8EJWecOXDEA5duTMtySSu2Z4NeDwS7
ShtI9KoFAcP3TI6hWUbjVkSENx4GktwAFyMnUHLT9IJWmbfzzPkt0TfmCuZQv9k0
WykklUKYMKItdZySh2X3VioTkuNl++gU8ENvfAT6zVScW8X2r9netxOZonkFiiAM
hxTioPCi5646z364mRbwZQMo/3O/7Wr6TGDHOM+TNWh5SO6gdCg4T+21laDXc/O0
aRLNNl76e7a2xqYWCxN5HUPvqTPqzYRx5ikOu/JHgUImRZ0VFk7CSzrNHJM7u8/N
XgUzNTwm+JKo6XrAEHk69+UA34SQq1clbDA6pxpO+mV8YvEtLvAjMpqLMANJlTJa
q7gzIouOG+PsPL9iVYRt3dwNsypEyxrwuW4WCVqp9TcYayoF/Vqt/QBq7nIY4TkG
h5sBtW5zog52ICUkDAHE6N7aAjgzHUO10k1z2AnjJkpxy3ZQ5+Ncte/psMTq26GH
IJMY100s2xVmIl0RxRdUCaQ4+w8/T2Pg+Vh3klRsbXebdqDM7aPL25Prt2NRTasz
YSCLCFoaCnM6YJgoIH0rkC2kMUKlIbPG5j7LlmM4NqTcZY5rSJ77V18raJcDelhS
HSeag2Hui6gBgWJ+yOSWd5ZV+iyl78lwPbdt1jCAhZts76zrf0+/36OqrQaLnZux
kZDcAsg5u6GSOkG+RfG00eQm9Y3SbhNbXpsZ2hk+VH3VdeOM+myyBLoVNoiFTeEP
FrTlhNstAy6mYTpsL5Z3JUda2UO9uJxe47FErLXUSLs8VdOOgnFPWChCKdHlxjXG
H2bt30xwtyyon1IrBDF6FWPYLIVWMZLpPh1f6y3LLUl4e9voVGO7LP8HyqN3QADb
DsrzSuxbb1no3SXEekN0kdxNBAu+VQgDJ/DQgYZiEDJdN5b0vMSCj2P4rJGy7kku
7A73ddrBfc0dgcBT/Mb0xfQXoXpi+i0gLPAf+wnXr4d8o6I5nUW+LCjqwXHlnLg7
xHahyhRDr8gOKZi0Kc14I6Y73/PcIR9gftV6f1A+tMSinvguRK8AcYxOtP9rWKlG
iciSY+A+ooS50dMkbGryYBW3ZgtjFrKNKh4CZCptYJ4VRoSwF7ZvXT7/1+BjhExe
ty9LnU9/NZ+kjCj5SDlceqfhcVyhyKLJzmzfwJijTXgtLEc+uoCZdq9e0V5VpVpG
AES+j6YArhOqvKJeJHFZGOVjvm3AhjMRYLspcoHQE783YDG9pcJHOFES7/bDiZi9
GWG9Ghmq3LXu7mfRuiBHqJqdgdHz99jCAxxRNj5ASXd8n7HAKwJNurZCvM2loOVU
9e4ROsU8UFmEgw4pkNJPtkZ7XnDJQFflvJjAlby/y3S8+8G41VSYXJDAsuiT4h+E
GydEJx6zrwUbQJRfi6kCMdxC6KPr1Nvhrs9NrLlZuIkN6LA9mZohbUZPkkiGLucO
Wrf6Lz9VfUMwowLgAlHY4RXMVScNLfZDhAhhbL4hY9049fSi4zMxem1HHGCp1am3
lxfMdJfxSQ+4oW5V5ywDnsjEFnc0Cn2L3RE3FQvC/Bh1wQXSwBJNfkiHCo+2SXci
nJsv0HUYnF/o9qBZz5Oi9SfteD4AUkljYFKqvfts5m1HTiBe1dZXOPhR+ndX/0X/
TEbrjOps1WQwUDwPe3mF0G1ExzKpYW4olQar/qhBPBfI+c+n/xFRg9gjeYEKPPJM
AUWiAlMsySm814gFumUZr/VygHSCxs4d9Q8WQQY3ggnQ/IeiD2bNPDlgtM+8B5xd
Mrb26EbDgKMWBSboleQwxJp4iwqK1vt8biH9iFQLMBGqMXYqGeOCEdv79GVaH1I9
iy466zFC7EnTah/9StpXL/e3X99fLpyP++44sdGPAwwwok9Aie+Pw0i/d8gJ6Y/k
CFDp8fImzqgCtLNI0pdcWT5325vjV7rWfwa6J9CDpqVbfXMNIXztrcTG660hMDga
8AsIHkXQRtYSULZUmgeG+mtPfSYBqxglsAaLbtfzjFL18PNd7gwZ0IzsjpKztEmh
Gi2bPEu8dLL2XdOzMMnyxZL6k4//5y/3Z7FZNKLEK7i4o+0BIKypucpBMBuvD422
EThu4qtxhjfFNdcjeBTaA/BYNzW76TUdhriugGokGEmsvFQowLTI7P9uz5f6Ht5E
b3QAJO9Mewqj/+XJ0LBuHwljbnmjQ+0ZSCNgqyZ+Tng=
`protect END_PROTECTED
