`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CyOdo7Z13FtN3maiZWMNJlCkTsxwckKiht6+wWU8GjrYLjylTMedZ/qZ5FQ+j7XP
OvryU44fjb7SR0pp0n2vQOnAQ7AIo220zK4vKUEer0qmdS16UhFnwb/GhMhz+Mnt
lKZcpfqTAj1Qdu0DwGhz1zo+oRSkMfckSVci5q/GTzaGwDJLTOU40vK3dDpq2P8/
9Jk/gTzxGjhu4FxXeHDnRXKFg0mOCxsiQjXZ5df3Ni9Xtqs+lIlFeC+Wl8FKsjIX
3RxfCA3EbwmhHxfhWPlSYHd+BGfqdzeIoq2D0OoYW7BtAMizkgsgIwS0cq8mzDjU
C5LyTh9KHRvYKMTbDiflwf5Ar27ytjYf6jEnWqUzWqIlHeMkTg7ZTZt9CMn2kTDt
m5iYVRjNS31uQdsIi3YkFnnzKzuL8iv38xkV5Q7ieeLpEppSWd6wDVm8GSBQ15AD
R+G6O3B35+uoslyAkfmfal0jeYFWu6FwLaE3hHmpZrknWOcCn6K4bzn3DkwsDtYt
OqlsXFlHtfr/qQaM1Bao08FMoBT5aCu5ZPlbr226PAncGc/VRp3M7RUEsQrrG9kQ
8h9HgP0Ov89P6h0LmPOAbDei2q8J9RMFdP5itxSg5FwB5aQJIoJjMFVuaUiMHI5V
WRJGVPODplWK1eCO0kxwZCBlwIrDTouKeJxqkYNGyEMqTc3iRP1yI7013EHK0jaJ
tSbdVckAnAjDbTD68KxYZFJxlK68l0GVXM3GyEr+xuWv3sIoM46Prr6ae20+vEBe
wy2kv7UT+LLywMTElfVdea8lgZmqy8U9vR2tpz68m+/qv1kNj4o0EoFIqinmOEVV
uuFKZuL2/x7CwxwVN+IziLNHVZfsuCg7AXJnU6ZzTX33/u4ZlKqYlzAqzUxwVxwa
nFPdPeCGoayWlx2Fc64GYimWYzFs/triHfIb6w+iObNxQ7Q4O+EQxVPzYdCeaL+W
bawhYlQadb90J46bOI6ownnX40/Jrh3Q0mmRLhob3BusGxCpB9Zhyaepa2WI8542
+sknHeVr7jDu/5etoaDkIRJFn+iM/Zx+NkfobImfGUsM+odqgMKXGcfEFhabDryb
3zNsR6eo4z/gb9+WuRBzczlNidC5Np03b9GGtxaHz9JTsrORm72e9ywu2gtOlQ7t
iwaDQSUIZ7bp5jzfgMU0LnZsehUJMhGk/PJkXMC81Max/C4RBeIbTeuHrOkZJBXq
R5qtkF4mR8HGqBISYvXmv3L3vD3a5AoRMURjD0y48d08uHy2XPddJz/uzQLZEPlY
FuLWvXqDkrZNeoQv8glyHMNhgeIErj141SJekXQNHf0iZwVRO61FMaO/ayfqBq8o
i1QoOxfi5p2B0alE2EWGnWs9HzUvbJZfvUQtiy+2wvgf9qP6nQH4BgwdF7ttY5Fo
cbjcEfCzSc84t+rtpCcSOC21d1QnkfJLhL6H+8AOp6GdIXpI7rh7AR9so2NvcUoA
c1NaW4AFtIZDiwNtp/ozD4xfdNEjC+B2uTBSU5q9F25unXiuB9Cu69Nbba+vhFB/
so1wLW3DQWFfnQ/ssfQsunatarZq6cQZB/amZ3nP/6hhxxMuuc9QpAcKpwXf/sxt
7UZHy1UIv7hHoFkpK4f6PKrcp4Kd+sASce2AWpzOys8GLqvr2j0MCeAVYlkLq6vg
uZx51CRNTdRBjCVsN6BOXKMF0QT45VFHAS822IJnEavbGC2h0n9UV/AZD33IlfJM
qUfHW/E8AsrfW3V9aWnvYotOOgQ2ajkqRNPwYwwuvSe2ax2EfNQanEirZE/1/YyZ
DizWJu831n+g00RSiyYdEEo2d2+AQfDILzHtfIeehovZkMgNMrdFfXVp33qbosdr
CyTLqb8+E+awvfQTEjK7JpnWKPFTtZZPYP7Zmf/7gNXpKnWF7Oa3ExpibirckSmH
wdQckn6Ec9OdHGAdceJJNKmW0Xi0ABPBBJLn3oZMt/hlwM2zSluW7DpZeS6fA9gM
QJkmOHsrk6fX4zcT+HrdlNtLwm/1Clxnpefz5dPYcwhB53GeIBkpy+xc/l2mN8Pt
PaiSiLpCbaqaYX9oGJARR+qAAGjyvl1C3baUU/jUuUxb5Godx6KlImdCywON6y5T
rEpbrnOlnB1s2tXE3QdsGBbpvNvOREbTWpmF7pjyJZjOASSRxK5JH9gUID6iJSDi
+8gZMC3F/dPoXEucD+aKIyA5twaBESMWqaqilm6y2IBu9q0Znxz+G67Qc8Tgt4Fi
LVsPjAqX8YnvbVWMUQ/72b6A6jdW94SvTSGN0GWqi34arhIAsii8wKHWPOH3Mouo
yw3lOV4fAbp0a7tqs3fPK6UG1V0Tkn5GoS2gC4xSdfvpwDGn4AeJJ88OMYZcTRPM
XZMMYdwwma33YYoGRh9FJjunl/NOv/cIwdn15EVGUq5rUWGbEnQNIRp7bpbs2HBG
tPF87xhEMBX9ZOvgAntAGsVkI2/OeneS+WgcXHIlsgu+dJqYYiXFVFztwKWHEp5I
zSQtDvOEVTswJ2TV22scab8II59T2jzOdIypaboD8LSLapM7Ew63ZbXzIvqQKtH9
uYxbLO8f2jMcMXp9vnMPc4tPe/BbqcmmLHN2gRhwUiUz3yGVE8rs1wNZOstjIlV4
Ee+y3GVZpmuTB4C2T8V40KWGNiGtjpMiV3U1yXzW9WCtBpNlwPbRXG2mIcHu6OWo
BC3tDIYujBd7ySeU2Jti7xab6tPmCNsM6M1TICnXoUwTbhfXyUBo9e+5JYYzwnv6
9+fxRjxx5WY68a/45eTa2nMAujTDDWjhs+xpT/JSCVK977rKUgBvQs0lmTHn4QAg
PCGJ8B1E6XyalFOAE2AuFEHBLrEtIDfuP9C+W8GPph486g5n9wbAmGNS1ia1ehea
xpR4fyfKMCf5har9K7hHagYguqX3lfu0fzBQ9Yg3HdpowSC1Xgp6UddkcBe+5vI9
v9mQ73mRvCen95EYuuygW00cJ+gI6kvV+xFbGbdVokM7ZUvZ2J+tCCFmemTqcbJ5
rc7wzwnfCeAOzO/KYkHztep+jYhuGLJTLirAmtk5xhrrUh+02XeWBJsqLPMvIAhE
z723/I1e4I1SEmG038G/J1Bn3kZjroCtsHu8LWAEiKI+GCee3t8/fwPVjSDIVFTU
FhKC6SpW/MWgqH/sh6JBfF+dQ9bYJT5zpTGXZq+dG01cejC77Mo7uY8e2OWhPDTk
RPYWkCYJLTMaBRIm6QolUKJet7+gwf1oT7fw/mGGu1ctm+lo+Caj+P5etm812yqd
KRq6+94bhtr3MlNNz9fJ/k19gu+CG/LWHf75wZWASkgBoKS8xFSM0cg3s8Thhdqp
mer02DlAXFnJtc8d4PhTQ5e9RNzh1SAT3WiHBON7wzsbwoxqCM7w2vGy80lHqXj8
D8NGXGlPfTOgK4AZuedKEXiEFEcQRdGJ43HshRbb9IO1/r22uQXudRX+h12gCvzm
UsI0lktZDXyjj2x0DfqSB6CVVVUWIWsUTNhPgtPMzKJ2Cv08m53LxsJwXOK13hMe
EsfYBHMixd6E1YOGnKxd0DL4rlRHki82AuW0rHmuFIntjopZbwCZ48vzdLh+9O/2
bKMexDMXBQ6AmBZjN5wTCAb78LazTSJ9Uogbz1tyk1oxY1UVF0TjH/oNLgiU7buy
iu9mFaI5t39oEGXNHeRbK3lMzLworBbH3KXwK4cexGev0KEc9zdDv8wt9XAOMqBV
q61Bnu7tcplRt4DlBEVHwFYO4hIK776UrEboQNkFii/nOeAsMzY5TLjsQvP5zJ7M
jr+0brPGDoX4mDX3/RdNKB5Alfp+l42HN31CSJq0KjYHQk1hDdmmxVX0wQjezzFZ
42crK8dPSRbP4/gwYWNCT+AgiFfnwYMdcR02CYbsnc+2Q/I5Ot/sk2BygVHlz374
KCXr3vkm1+K1GClaDg114JVDSDsJUaL16ljgWjR6Op+bdu4qUxpME+UAOpyD2aTL
Zj0xSd/vHn8GZOQ/to7SACDXEl+HcfNFh5N/m5f48Wq2SJnKUciyXNNDyAOOuRle
5Bf82I88Xcm9QGRszRKCZDfZ5UTqK+gDrAtWE2fykqOP+T3zT4OLXf4Y8/TCG8Ti
q95aiYXb3Q3AEwr0pKAaaDNJPjK9i/67ZjFTKeHxEl2wWLH/Z6c9xSl0P7nUPP0Y
E5xlIaF3Zp6oNC8sMyE6fu2/Ad5T5V+Lau0kdv+ym2i3yfsftN4x/UD2RhPOQzm/
9v5EfcuPVQqlY+dBxcfViwnpK2lox6nKOdwP6kF3wFpvWGqg6kk7nU7G53L+WUx7
oZAmaMeTFaAgtzYx7ouccyg4zH5cyqkM3Tj9fm0LM0+SNRVZSzXr2Q0nO96thElK
+JRfqsEVThIoK0e7LXiSPca7Fd1y1zucCw8FYh37EHlerRnKwOxuPb+CcvSynrZu
xf0BaZlhbVdc86S9kYaT5BrK+ffd7U76rLJDAdg+dmw+j93VfDd6lE+fgSHDf1e/
llrcS86qz+j7ElZSvMcHvWfAWMA1ZvxBhyEySEzd8l4s6JUUxKmV/ltJhOzIiMyn
hDRGI4J6/PlCb+6jC85wQlo8gleKPqB5akLh6VK2DaRLuQA/zK/JkCysZa+nAZkc
0HFN3blzxlOqai9E43srXXKkY8+/KDs0YuIkH07oqFv/SD5GbPWTLxkn/sX9VZY4
SBtoSsX0c8ny753FKasRLoGBFczdryr+WzOPVFRgJ4NjlUw3m7/W1LEBOywpkI4g
djkv51DwvaSGaTleX0PUO9K4Jn6OYvCNRyQertbpLIvtKmsjtgSZ++G0r/KZWwqw
1JvmxOZnkkjGgGWukEtLob00tWPatCYFhM2NIZ4stfjXKztq4vmhuh4m/OnS5g+o
zjdaaIVFb3DwfkSbMU5WHzB75GMulBLiZvoKmuI5qLRhaEsiX4YCKsNChRX+cpd5
7E9V8z6DlwJucJAY84twJDgVCnuYszFLHThfTQsqmASyUd2OI1ThKLs8lVgRT6G+
R74fGj0mJvJVw3r2S/MrHSPIUgMDEmsu10d6xOWvOTmR5X9xYpCgBaS6Lu7NcUDx
mhZkYYdZ/HnN3oJSNzmMrkeUHI3CYk0CbqjKOCIK8NGW2Wa5WLuQmY1KYeMwYWh/
1w6QsnIAxrxFRzPQNznxc37kDQjzNCpIQjsFnyTgFswAfru9pNGy99yKnzDHWBon
is9eWnCUh0b5tSgt/wJg9d7VZ8/QTrgPm6CWnTHAXhJM96DKNifUzW/cL05b89aX
BiVkEh0g4pYSm9Lj7h6Q7ETLmEGqUv5+LEFiwKVGqlgV5Bd0pIXUzAidwQOf+ZQR
x1mtVkmUzDeKJc/wMQ6yRAAf/pCRlu3Wd/YyFOCaba5eakbxzlZ8b6prqRaAcUv0
qlH6AcOvW3q+2q6GpKrlJ9NGDY6I4p9QpL1ep0DksAePulKf9eGcSqCzicUfDLr1
KppT+R3z0+R6uUEBsvsRt8rSSntVBDfq9A1r7j11bj7yeb04xtl0oYoU421FiuOB
m9nUdc41A8FOy+Bin3Vcgh8vftpJGVcr42V4D+rl3L8Z/UkfWQy8kssBpQTtdlzv
7AJ9lnViXOa1vhVbXyEX2Xouk6qoolgT+FjiJ/mj2XXkk1t1MrMGDLcx4w1PsilU
URvvRRX6cLP3n0EzCj8roY8Ps6WuI/XGmECOJHBVDBdRGrXtpsAY6zvXb7pVZRBh
aU5xH0vLvmL6uoVOi69IppzHYGcICRudMh62qBM7n7yp864QdhmzZDHUBu+XpOSA
D4mCLq8vi/9k5jjgaSCAoiRrfT79+H1IRlKihrsfee+6vrX6vDKsxNeYfP4ymvtK
EUhuKZVW80sV83BooqHquZvi2Mn4nQAJ7rCY6OQ6GWfrWRdIJoGjZBR9lx7ZzXCJ
9Pf2HHSC+nCC9sqpiDO68/JFndl4FmNPEVoiOhIEiDre8ShwpuGbxR7KdpJrNzd+
Z4nOEAYByb8gqt7OKTSfl41dIoTlCPWupLZ05UZTva84ujbaIRGu7l0q1EO71Vj2
3Yx8+h7geCL8yQDIqxLppPozzTIUCWcu3nSUvH6n78dbZifs2CNfsra2WY9ESRt2
7MYCd3ur+DP71mLmz6j0WwwGXM1LZGf701PqWdfmOMQvOQHhVpsxoLu+S1H/tPwF
k5FRqnlNiuaQF0NfFiO858OEZ19wjC9FUZ62xPECeAJ2kJlfx5I2JGS0fLGRrMCp
V+3FviPqgsaVP4k3LxRwWDEjibjz1LYZQMJiUkVbyieGkxkPG0G5Dat2qq7Qty6+
1FbGY8cAloLqV0s+Am7QS7kQeYYDnZsv0wunpfy07OoXUG8yl+ZjalNtqKHHzLaf
Tm5oyTTNC+VcSuM6prL6lyXcAAapKm4IhDJpZSXSPrb+G4cFX1HvxIbH3rMDw4sS
CPJ7iua2tWsSBv0iLthFNi9Mbi+MKsBVK/Hti2j+KpIZCitDor2geBsI/mx6ugkp
6mCl88H3a/Q0q2zWvkqBtvXQNpIUX69ICFugdaR4p9MbIb3K0ueM5JMP4QcFi3Ej
BoQ4LqFIh7G6hpESbqwEVqmnHEMksWazc0r+hI3nUBVu73cDlrMrJ2JHUOlRa7OO
BiMqRIafEQmsuxNoIGPy8fg5oTMADFQw2Aljj5+FIs7ZkMRSrYBnCdhhGain7LpH
mWeiQkjvNejkVoii1OYol8/PR4h98hZj7U4GL/6LJqsg2u9jI6GBD0wrtVC53Ao0
Qv9x2kEQlHC+vZrBp4OlsB6EuKTlI3ZxbNHuEnOgsrAKl7Wax/ihGdqsFrlWmdd3
OUMyNrJXFTefD9VB+jWwunONbn9BEUdk1tCSfrV4LC4fP5q2SwnnZ0Ik+cJ+pSvs
WaDYZ3oghKXaq+v/txtALLLaPiKT2po9itGd1zYyEpQduiUk6EqZsAvISb2rb/ZV
LbeDLz2JCE3Q6jgr8bGXkV3s49DGnGf6E1SkdOS57qbMnEl3qnB7czf6y0ZSD0L8
jtL5DF+L3KyG89tblEuD1Lw1bOajK9CXVM+9tHIr51m4uGWdhyOInkELAESo6VqR
+/0S+yhaheeAbxGHG2hpVfpss7x25adaiihG3xMSheckWtFQlBUfYw+YB0npHztF
UrqSZt2DvtGkv9z3YbQMZuemTV4qrkjq1Dkg+JhUIdGIoo+t15fpJtxjGxegdb7U
O0EX+ZSWfr6gDEzFuDxhPB64HjnFIH4zAtxPfqGvDpqBGwj+berDhcprBBL9836b
4qlW+KZqMoTLymvwSiTSxRK31l+z1WTLCqkYqAu8i7oO7qiNQbFSUQRZNFZyah6g
ANWpzSfnbAAn7ATVoqkQx6Jlgy7g9mpDTNYf59J1c6Fjj/5OWosnlO96zxxLwVRQ
Piou6t/q7VhiA570TxgkvYalRZXz7CQHvvHtlqavUGBQOi5lGc8XcHB6Wkc+drqI
T3c7UfAg6OXAxtfKzKqr//6YcFIXBMP1GYW8etTFSsBFe73Ck7I2XwkvtzmebiBD
hk2wbvb3stPmmSFofvOJ6jvyUt494znlBYQaWW6Xi+JwWe6Ab94QWSJOhuj6JxMY
yI0m+kGSV4+80jmqo+9lliemJFMtbAqgvPCE/149N+Xf45VtEkWjxrLrluOxjtNX
D8Q5cBlw/vpXL9PqpgoBlis0DqeLr5XZRM6HPhz8x25AW3F9YA+/LHYkjv/sDy+4
pXEOYrELoAv4rlELPZqJKaqEtCCk++f3lcDn5UxkKi/lTwE0QXGlIti1PER+vmJz
L89GV+x8LKUI01zrkq44BjQo/htdG9ZSehg2ayeeIdAtE4lZlLBwy2RtMxbgRXH0
Bj2TiH8Rr/kKq3nzRLlN3YbRDLdKN43CSVeOhW8gwPibDQ5vCBN4Mm2MJ+yjKF9L
uSJ+LPdwuXy9Dlrk5jr6iVg8y8l18udYFJzmw4K70cPO/KdJ5eq+8PTn3OrcILsq
5ZsQKZgKaXLzo9Rl67qTa5pApdKjKZrATLlv0SLHqx79WDmi/lHM2XEbzy8j3WYe
9iDiP6+z8W3hgS/y7Hdk41xbcKGzDeLWloUq5zwX3/vIUxzYZ6X/fdpXzK31qGF6
0FzClJdkIa+VwvwMXQRSg7uOZ3Zu0/RBYB4mFRIRw2EetQBmcpDVRRutj74RbzxK
RTajBdGov8NUdtLR9qUdyukOlBR671setfwL1gcOLERYq8MIhfIcPJF47154wio9
JvxE1/1G6WgEO813Dzepoy33eg2RXIyNAPJNYlgLSwgbRRmpzzdqayQSbad0NVrq
11T6C2Kgmwbr5KRImCCq7bn1KLWLRv5P2cdP8AQn0zKIbKIEbFDFhMUFnM8TGT6D
Yzu6IEmPm51eOu/WRS6BjOHuUgERNGawLs4plpTqKl26Z6un4ut9EyeTX8TyDYT7
WTfGO3FD6kGv06sgpfbRKqsuA8rSBCfzYd3bcDiEYQayUPs3ruXuBt+3sXcT9NzJ
x5s8zevdXnao8qUUmLtD88rTqyUHEZh7EHTEf+pLlo8lcfo4Vhbnt7HuC+vNutBi
S7UfpJeibmgSbyaankLtGdbQPJVQzBLCNVWrWZLtqOiXrPnkejHbgg0IUAaO7fpL
vlGOfn1VEQePcZaaD1gS1qaUrmYI8wms3T/E1YvSPQKMLgpNq4S+4xF5RIQelP5l
4sACVwymhVIU6nlU7oVPIMx2P03T6TWOlAnYHEdFwKEHzQaF1O44U79lLdS83f+p
xUC8//EBPEsP4i357LxXV0l5IvGuHbQoD4GK/aAoC1uNSmINkNr2R37aVn0xbsEW
xvSUgPSLpVZtfACZQRXB0mZ4ldUPlF2BId0uWQ7mybqB9qN50un2XeABeyFmvNzb
hJ/9bJwSIJhLqAmxkLIih+AFFDiNrX34Ldovvj2MpaqPUoQXz3u1jKfeNRVf5a9h
6Oy3T7XoTYMOQ2mH/P+LcitIY2s+86ghd1jrtO0aH0ktv36uN4fykmzkI2/d+qfF
Ruow8wCzbar4KBNsczXkCWfKfc6O3MU5zIBjgamleqCuT1twuGtrx5NbV2WTJzA+
EdwCtXRIH2ia7GwKiNzQP8MuoEc2Hpnl0DFQDPmsyYywvILmEJwmCF2k/jYB6QRD
L2Cf8qGjTkJd54KI7xd9FSFywFfIsYPNoOV3KIlo+XD/sCnbgbH6YVPJ9SSX9qNk
7boskOspzi9OGOM0nDjFsZu5Ydh/LfjGXyIMwNFOa82dlN8llsjE2CgTzfz87OY9
cP68+yvO0FCEeBzumGwHBV6a/9doWha/1jprOlrx3V1UsiSo43XilfvLu8T+7Xuv
1aDxy11f+cM0GlcehuZ+zGvTHUDUAcF0Iss71atZ2TcfvDQCru8lhKhw/X4B8k6U
f2WcalHi+vJWQJhDfpIqO83ePAWV16UkjzQVvms8uPyr12P9ziWn7KkxAvUJ1V+5
8L4iYHLR32YUjrsG8/QhQAkeQ3EE4/X5dHUcbLHcoZM1ixmX+wdDkMA+sl/XcC+O
pvWJq3nVtEOb9MlqnNqg/xSOS6W7EL60zT3GSnjFaQg7q3QdhJPAauqp/1r/ogRD
T9HqzO8WVDt8S2l2CITZnQLpbEWT9/D95JojEEDGnolR4EFgAObbGpbM/5QT33S4
xO9YYL2Rf/O8RcBVFgxlVy7ZjS9vm514KIecLYvEpGhqEgOW2nRI8dQAj3CSF3dc
PHNoZcj4vZG5hChCXIwyLHsyHZxDXBAKM2vlmIMNiqek69KfIKGv1MymvU22IbfC
gVXSm4ClYLJCYmdof/uny8ejCZDVr1pqRKDTCoseSFUFhq6/sWKxrNW1S93AWPd4
zePPEKfyjkOFZiggsCyddR/aLNQxcd86w+EgLtTe9LVADj/xr1hmIbi8DjOhpDeb
zXAlOFUzrv+RkbQfCs/rhdZgtYQWV/24nxFD1jZF+ThIuujijAS1xmUvEQ1QbJj9
UUU0ZxRNaiibXwwCGbCusxPJZwqEP6O3zaJotGmq6lxlMXvyjYFT5leCY8gEvNpr
NZeHayGarIfEQkzYnalxzQPHP9NlkQ4Ws74tRXyMxdEkvK/Ld2OAgDcLYYdwRNov
tE+TPhiqxEhQcZT1TQSBnA63Zx4cjIVIt3lwdwjs3vxQRRqxmMnyM92nbMi7smAT
FST1Jxef0qkM8/sl3CH0Qq9whFXYdZWF2DPMKMS/zw+OFpypmZaKzcgqrneJhUPO
t6UKCjoo1Wx9jUeVVWY/PDVpT0+hR0PPdDs07z5wVvk4nWlWOpn6G982g4q+LDjS
6OtV42j3yeE/uf2ptLSz8omuSWEjvrImrAa8pPEiAkN5Kqbn91QDJD+qcJP6KLKl
pXozrY/8SJIfYt8AODnJqWkHpXHAhJ+8BEm1aeJF3OHXZSvpa3PwFwRMCDDGSAJ1
5NPyh2XIVjY5YcTSucnMLo8rpPQ8I/eEz4+OyYERLXwz0jS5SPVU7iYrIv40TD2+
vUkXMeTZYDiEpqUfpEKq6AYXxg/9tnJNrfR99iB9Zqek9whSHceT4k+71JWwBk9q
MXbukDuw5mHNGj8IsrdJOjvMNwfCJc4W99A7fQS6LKc/cIN/jJ1phzdyan4rfHAB
ZoObktfxIt7KnC3aXGNqyGyNq5QwutuKLhPVaMv/LNnzk0LdpaIxpVQ5MmbzCt0t
ScFfDMUerwdhwvAwbNf+YriN8RDnVh+/DdvBKysW+vi/GoDIiCOoDBTnSW4i1zfV
LN9vxohjedI/bDxyeTqA8RPHAhJMmXVlVKbsI9pkGcN0anbyiABSENqZ+BCPFNYq
nnU+MTGP5wtW8NZ6nJ1OfptnXKauMg7EtOGivxBLTV56OuHp/RAOeTyJn+8hZH7d
KvTKZ2fjQgKEhd7uMLUQnXrqRlshApOhNSaZfB1WVGCYNeRCbGiwSX6TCIt7SDM8
oYhE1DVIZOu8rMvTd8sxIZEExyTfsnf+FKFEs3rWAyrvDkN+lsCT+gXgrwOvzceF
JcCHeGcdgrKp8QUdqPDe3Sa5ZhVgjhV4f/ejbY6dm6prq/ojAK/RX9Vxe/qBabwD
BgDoICm2uSQ49kA0UjCIl+fbijuVwH3MVh5tnU+JOw+DkF5RC0T34y7ONmuDFycz
Pocc2C7hAbH8zI7bcPvJ/6UbyAKIVBkHY7HAUJPDXKKzYw5V/YpA4wDvKt9OqIu4
ors5Imp8HIKaWVRMARx4DD9yHSDJx177zUuz3YCqmodMHEK7KuA7kLuonfisrrs9
k6evYwgzdVOg0lEkZV9x4kCbI6ngXcY5ZpvePUyAxR9OkrIOGIxzHnO8wX/yTI43
iXc74y4K5QZMOzcgY2Egv9OJ/pyEAQRqaFqAAMd1eVOQT0IVlm2S4+pIBB0xzUP2
/tmYuaYtKoJwPx9PYSKhpdrbZcPMKRhI66UIhOTIuR2BUsTkz8SFi2oE6xODbA2e
iz09x+CX36+rGN2Fvzuo+4OVOarerLi6SJpgEySpo1m8AAgzreQ0J0G/Q4GHx53S
i1hNh3az4U3J/qfm15nLsl7ZgxbVIe4ol4GVJhqBR20zt8UfGah4nt3UdTRkv7CA
4tz/pm1ohNO5O6PgsZRWCMSuF7V8x5U8etTPo/xFg54BHU8mII2azfS+0ZMqkE6M
PvKD9fi9/2OADAjAmfbp6maFcsG5MG53PexI+Y2HqYgjXHQlJwQytEfnHkd1QeBY
s/ie01fKQnNBGByCD0x7aFQK/gQWCA8oR23GjgV+tkb17tPOt26ZaKafrxrAR6NW
LfxRM15siDIdHPJZ0zDkKSVp9QkZJppBxJOYg1KWBBg0DOqIdyKU6j1LwomFEtZC
akMShaLwKB1chdBCNOVcsdjXaOdC6GaAVK0BLCe6C//HzKbfXaC2Eu6a0dfHZM9Y
zH4xKF73jEBHOyeqUqEVEwrLgjibjTQofkB47tG12VG4XF9p98Adridxomi0nKbY
iIupsQfWxZZTwam1z/mA92PFSXJVS6lWlumjoozoft7trSPDrtkfStadnAxwPY/X
HPWOVC+AKu7OQYUYoSB+x0dHmr3SsNloG00qLWDznMgy57U70VuTb67xCooov8Ux
Efwe64U5mPX9ZF6mqIK4uXqoIpl5R895b/RH66prETHFm2439dKBIlp5P+cioPK6
ncrEWk1x6LhXbNG3ParmnTDwM4wAX1wNyE7pj7DIlkx5SRrb3I13WwH7Mho/nhu7
NvzJ7M5+/a/SnyKDrYjWv0qyX24icH4J8Z7tjEuCI516sLc8CIqj4YfqHacT3aNF
/tONvhcVn2puBdc3sY09ZZyVXRIlACUFd4fIT8R0ByeyabYWUOG4++UdwtACz1w0
QtIwhErnr+wI19HqjWJLZq56+0vYpto0v5HGaTXxksYsO+qmUw4jcNOLjhWqT1Jb
En4ir6A4gmxUH7UnKEMPn8kbdoME+MRtqWv0AMezCJxSWVIunqza2oIsqvdu5hCl
AEfLc77avVjBiLNL2tpUFIFSW5wKZew6V6bMx3KulVtZ7K7oF4XMtvSKQkaqlppL
aNIU/I6VIOwAGNywJoCjpZTBWiRthESNW1gSdKC/Cx7HoO1+w5sdpnJceKMx1V2l
qtiZBwtu3q3t27z44pV7KOu9PdB/0tNvE025+xUkphoiYfKb46TwjSIpFBZAeFWP
elg1fpXxRn+hnxGMZ5cZjQDfmFQAx6rKmanInyOKZjvCx+nOxwIUwTLLd4H9R23F
krSX8q/fNlmU/t2fXCzUccJUrOYW1S5x72Y8EalpSNQRFRnjTPj683v8KF84Fi5K
XnvQMscQDkgS95RNuJ0rdHtRXEpc2CNDmmIxbTrdcej/7u9C+o99LXNO2PBUjjVz
DQEOuznDC6unD22goW/tC3v/GYWxgfXF9wt1yBRqAhCtzoOCFVD81z1tcfQrdYVe
J7HddVyKa+czgC7E5QsprP19/RQmkLfMcUIN9mUlqrcqFhPlJdxZitnZma0TplCo
oyYkboOclp1bf/TK1RaZd20DyiqAo5QE9D+v+HDG53LfG5JAXzTK0qiZAxu2RdTi
WYmjvN/5bAmWQI5+Q/XBMYDA2DiX5BgcZl6Zb013boLf2ECUQz4ehpmFM1yfnO9V
TIkJgEIpQ5x+XGUWxg5NTgVPLVR9LzHP7Zin0qDMpY05a4mS9G7h2EBw5kgMkw0h
5PD158Ff4Ccl0JCm4rEd0mBw0veXTUXoCONFxeWYCndH016gNNmjSpOh284C2s6x
IPcjK2qAIbRmNoNgdmTFL1CjyT27p/ErCWwXUgOLeWVPN7DYsDUmT5dV9gBN/Ny3
bAEOxD0Xxlb1ev0Y4ZtJAhesgEeg0GLxVolAXX9fqE5lqQ10wBG6rjuiracZoNt0
ge4Rh9MtwdgaPSUs+uBmmRBhNtqzuEmwWB/umGQwPES9WRjkvJ2PFZvUfO5un0dH
SxdOTt6WeuwQbICsfxSPR2W1pzZJnugyC0KpxcMdOwMRzSzbGRQZ7Nkdo12hoK9B
9bU88jq8SXqxPPuFUnQYamSdFfKj5rAXnWlsPLXm6p01gGGbJC0ZIS1Gtgfd26QQ
SZG0i5nuvhzfW+6V2M+zmcHgaa46L6zjqN15cgDpLkkiG4n2IlDfwpcx99e+mKqZ
aLNc8h3p3l7USe+sVBdN9Go00S39JxFyxrZS/dDdGSkY7mapYCAxhnTIU2RbVV94
Rgn/v3l2rlMLBgCzUWO1GNWl571Cy2lQm18dm5wy3Y+xuDh13oVHMy7JdDGDVj1j
1/3kg6ODn4xqD2+Vdatc5Y7UCEDREZbV6OxwlHcO1Z2JdNN3MVVPtP3//LeXXdeE
+8uzY/0eUqtt7mgZk7eyDYyGvQGUXDf6Grff2lMBIYxo4yDUS6W9XY0v7x9x6qiG
T8wBeseGppNyJ6GozPEhrvoxI4CkX4ol+Codav0ywKTWGofjsxEt9QFFRz4FJ3Iv
3HOsBX/tvDPo92fbaFouM4IbM4uBEqPl2GqHRQFbBRg5NC7FEu1KRAMegRkTBNJK
SEAXNP2ehj1dJUM0C0sRa38UXK82YIXnsfwzms2uOxxytgm85RnfdE+HIMLbU8C7
SARWTSTJKwrp7WAtO3/HIBL+FeFupj5SWLW/f2Ix/xg4KE6apNZRn4GGtbB66l6C
HY2+95npKp/lmcp3P9zje4nQ5Ds9+yViZ/sycpMNW71qgsfFzmdOKAqqeSKEKMQw
j0EayyL/5GiSWucx+UD/mZ3ORXmPJb0t5Ggbg7/O1Nq7NbLLbSl5oEmYVR0fhiWr
tRae1XA5cXIxm0zR8AAfu6MYPEiDIYgvUv4CWGh2x134cXTJLE+bQFWMh5irKtLt
Wb3//VMQNLuG70mKisK6PEOD4ss0EdPBtXSzW2oyuIOujq4rR9FptZRV0XT0hLq3
V4Q9WQ5LcdeFz/86STQam9aVzjuIkoKqNo2WsSspTVIVbodul34IB3YJ1oC2fPpL
4NFEXQxbc1qOMktnEIySjPqRg0lFGmXK7KzU59FTu6dby6JU29GNECepNXYzyYox
ByFsq7O9bYShJCJH1fo4SaPs+D8MLywgZKkE3b5IdQqzMC+Wmj05YARndrkrKzfv
BOaVGzrMSQYCeexup897/Elzyv/oKn2fN2j9KnNCCTaQwJdFujuq3aU48fuHSveR
kbGTCYOLwOkdNCUSaAMekHUvfBkhjRVTaqXjf7yLcTSf70NvAi6Alfw9oBQeYgiG
Wwrqtq99ozwMbfvNmBu3bSV9ZtxBjKwBFiX8HUsfIz+ruKxZfClaT+LC5eUbwjG9
+CtBfj600ALryVf0a/0E6TNo7JFihHvrjt82XKf7HZYCQR9EXynttLfSNfwkRM/2
9JAIBxb6F1qitbl/Fha1zqDP751wDMLAJrhu+SVG3c5GzsJpz4FISSSTml26xKD8
EJeDx9GyDOuJr2LYMLjtekIkxi88e81I7Ew+1CfP443BcCTQwncJ3ZVzhLKvkTK3
IdrXSZa3erpjR1ipyDbhfIWW8U6TXntq4Gu6L4PiHAgfr0rjZNhWEJKnImeaieFM
r0YCKKZqO8kMo2fUcLq2TCTJa8KvAnkcxiu/Zoied3pedZTzO4MuTucOeCU93ANY
+0WKtiaSABrb7xF6XTRMuJfqHqpbSqaFG8KkTJ2+zRIX9dvH8LUV6T+7UqrOHOzN
8rR0mG/qieDbkzbQyjWMi75gRs56vDN4JlLbcrNR9YK6Z8oeqXkC0pPzOvZzMSBI
58LTW69g95EUS/aiFTrD6cY7oAYe0a1WY7TyfupvhZpDkDrsZQmJgCENcX0NixQl
na9z0Psa7RhBP7Oh7N99VjTiX0s+Ny/ZyJWSeYv51s6f4hCN3VDyWFQbgT/kG7Pp
o6WDna9/+HqwrQm8OH9Kbujls/w7vj8saWb5yZsBtv+ansftuuIdbWChXbzEsWwt
IN+tfsEKPGjRt3msMkIF9i5KITrPJbz40x5Xk4T7R4AaaJunyVkL/vrK0ZcranEK
1oKHlbNHD0UEjO56Fe4/e49hDVeDRYsvPI2FdXWp3A/DAKtGqOGrwRMpmfSPzZEp
Nfa8PKEBSzQRM/qvKLM/t8m5vClDJMfeLWWm4uUkNHmkNMZrd28pzTPSsdVJy3ps
bSDscmLZhmNHdgmxEO6R+TkOGvO+v4s9duPo0z9U6TjHKx+ZTJL9AasLhbsn2k2N
qbEOGuWjQEoOewLFC6bIkpWY93OiCBIcJNhbHeXYBFBA5gOSZ/QBSqgTNGebpBL2
5/AyQfu/HDK0cDFDp2C4BcpO+OsAwZ9bDLBRklSDpfwxiRgUg+xgec9Y11oKUMkw
SFxamSQQTH4HyZ3SIiTW/tfKTxzSe/WLFLgY89uBXHQQK2iI8cjY6Nmdq0uko8/x
dhPfml6PK/KybjeMlWKbE/LwYpzmfKY0zQ+fH4jsv8rM1+FSxB3akeoqQhLit3ll
rLWubeDqGAkwFfr7VwMa2IJdkzACtMGf/YLiWUT06TrH61e/XJnT/j7eyPu9dtWt
gVW6ZqyRu3Y9EFUEdWOWLGN7KBNHWPb9igfkNecO0DSbzQFKZGfCJYVbiZogNsoi
kWElM8iZpQQQGG+/ywj8zGslBmj1wnOhDbwe+uGBohCL5Qn0Rge5GdTuX235rVJ7
kHcJj7QYV8E02YOTy8MUXmZeQTzwFSTHs3ZqAUUd1S1qAl16z/AG001qtj5qYk4r
p5RsLr3qcIl6Y5VIdsDrT63w5DmG+6CLatvnd4p+xwDc1RoIhnPSmQFMWKSkQ6vc
7LFG+n1nGU2oOv0SCn7Qv8RR4K6k+N/wE668sbtKmY3ARSs7ROQugWtk3MEqqdjn
Ts8pppfWBx6iXnSCAqRoSl1kF1FjwEI5nw5OF8TocOYOkcZFvm0N+UJKHQKiLni8
jXTWuJGw1DA8oFMSOy54oMuVdlmG7We+1Wlq5CGKSpHonVnYCNw6eqxLL2eY9C7B
A6yzSAwLTNxEvxDOhpnQA9um/7lqDcLQWkzuRtmHaqgrt/zv2ffuzUuNz28J746r
yl7pdVpZy5L7wKShzE1r6KiTRWYL0QNCXKCoAXa4fmw1XWgqPuY54DMyMuHaHzl/
Mr9aWcCwhCtrXE+JMmjVTn2H1/lFYw7uHw7meYzV+ZTmoY4E15Z8LXFZPtnL9El7
1Q/wUh5fK3uDFK8QADCkgRe99UaPUhEgCsfMw0OYHRzv49MCDvw19hACUMoLjKVl
FmbRFooMVaAG4rMXbWmIrjaQDm3R4eaLRfe/3R3lX5kuc2IjrBj0orkGXLy7QO9Q
fiaaTDIFXmPvU3wwT4aEj/5OHc3Y5QVoJS3uezdizTnFGT9MMvpEOH4FHSBiGtjx
lUmJa/UUsUNgtAZyUXSDlaoUS3Kjcxw25TX7WjZp518ORtlx0SR9kxwxV16i9Uzc
ZqAGyc1JGN8lXpJhtRPcOLYsMQH5VqUr6XbQu5gUTIbhVC9vMB/K2JTU3gvclbZ8
ZQCvPVPHDH0N0P239mOOhJdRPRVjbGsgFQAtxQ7bFyT40R66HItFgIT8rnTuTL4R
k+uWWdJWQVOOzEr5bLjLyjO5TnTAdPUQ5jZ+J5Dl4JoU3CS6lXG8ne1HajAx0t4U
S95+BC+WsQgU0R6+NJSDRjnWl9oHuGvxq7GEkzxAokzKuf0R3etKV6951rmo1GjN
KFuNX346bYz9m6p3907C9mB+WNXEJ9x7L3/gjucQNf7Oq+BH5aMw/maVt6ooek8o
zM6qwGhZW2scvNFT+K2698X3x7+oRnZEvtilQgM+tG3ilADhg40BMKiVvIoB01VC
WMKAIYDg9xi34d4/ByQeQ49K/5OJjM9UMQAYDr+5988+DnxLZdBryKULn7CA/RqD
R4xe/PKjT5GJnjpqbxzvfRm6EGtL8C1of5qhdpVN2Zltwde6NLZh9iyVYzuFI2NQ
Ee0neh0awA//iockfsEXidAaQa/C0Lurh4aoWcMIudDINoqT++w7dMNEVLy+iH3r
Pktuco9rfhWtPYBNcQzZ9HDekZrsivkVgu8Z29rwp6PDUpzNFMyYUoVIVg+NoFZn
i6cOpzOeQitz/Y+iibT721Rr2k+CeZ9zAEGecPlwBKn4tah51YIQGquPoQq1Jvyf
dSQWqTnpxX23mWh3jIIY3QkZq+mJD1+XQsHdjUD+p+vz1MD5VycfiZAZLFrxXct+
AFjEm8vl+TPM6u2jq7s1YSN9+6KxlTWca84+rIzROQ2cfLbxWESGsCZPZOxnRU72
izSwTyDF9HXDaivWXFoJFa9+DWxb11Fd+wwWmKMxOpsd/+SzGNXOIbFaduffSyUw
7rclzaAyjEC2DeCfdkMEEeE0NAK8bg3HWMMpJZbHMNKvh77OuzQROdOJwkINeoB1
0D/sY7xPrUYG34aZs/y2K3Z22xRH9zhGzqNYDr1ZORrHlAOntH0uvwHvByXJDyzD
ZZbL2AJhaWUJj1GRMVAK1cSxRIrTkvCG73ee4LFLN6RXasACJjQhRzDPwJOhkPvm
q2RXuqeO5UNYaDUM+423JqgJu+34mQVM1yl6/xFAgqyMKCzC422p5m/3shXVYO5Y
d2db3fpeqU7UFiHU0MyG8rU+qk0ehH70gbm4bwXDz2/89KUsCFhpZO+VFo4ajEA3
8jb+7h+kRF9Xhl62122LlORjvNl4Q4iQwcujfnTAnDKaB5KfVS47d4E2nYUVGXzd
n/6z0iJGRdOkcZKgUY26fCKrEPNJ+O6CiXOvUgjVQbSy+J8DSr/6TBQz5YzymNYp
6iYFpr7IQrsWp+br26l/+bhjOIE/gx3zike6qQGjIcIU/9BMPpw6+EBJgfFBiRsi
5EMj9pPFMwMrWtkJhUM9QgpXZRJnNxAUJRKuQTRjXAZ+hkLgV9jr8sNfLNj8urJa
mZxHJ6kQanIRa8CS9+fPpuO9navahRyNeq6MFIfSVIv1KHJzmwIxHLhCMAqfJ+Az
f5qac5i3EBjpGOOGKuO/Sl7wRVakyATsvhWa2G0h9cI/8lLvGOm+fjhNjckkjkrJ
msIObdaB1Q6YyAD4XaloVy/z3+Ln7Y1EtfHuQn0lmdPgjNlECFrFPDmeWRt7BLe3
63oaUZagt6hfnzmDVABQl/GJb0cS8DbkA0YejJkYM+XgozQmFbZiEHiqeVClzt5d
ZpidbVIEfMw7pat6KUYuhsUIbiclcjj6Jc+3U8Cd0sKvFq5tqeDZdEXsf6gsZjIZ
Xcg9RLwS10OT4+5G2BzWgEP/fZkJX9+3w1P7116VrsY3pwJ8IpQNPTVskd5P3N42
rGsmcf2si5DjkQIwNtK7JYaHW8/y4BEbI4sak1/PiaM/55b0LrNXvsoe37lbm1u0
AP51ukWh1qYnv6tiE5ouUKk2b/bJ38Tyk4pGhy3qQJ22mswPlsWruie6trmqcNLE
1MNQXMVGAeC52GXMYDRkmVmBcBIG6llxdEyJNMCFRRJM4OG3dwrgT+9ZpZ6v/9f7
xw14l1BlBpaFdd2iJWWs0ARsVqc0bhMMPpA0fnUD0MaCpwuJl2Dj2ncYwH68uu/V
/Tt/dbkxAGhYR9DFwAXAyGKOJGyBfyf90RsBWupNeKtUeiBTgI++9YGfHwmUD2r8
YOXLtdzfEZOmAvRkVnx2fIneSScOlOH/b9LEnBcwgposQkUN3ZNjfwcg/apOvD4H
sx+8oT+UUucBhjVfLR+n3/JbaWI2+VCEJEhUIgnsT6DxvZivT0qmWZkTGp2XLHqh
mKaaKz/HYqJOT8AqqupyQeFGwlh0DfcY9/dTFPxB34kNuCFVt+hrIaticH7HTFs3
aoYHBoOrklN6M9qEcAzCiuiECEfnfAAPDt4NWK75KMYCDIXJnYCsh+WrBFKg10fu
KQzBpoZz2358qImMO92F7R6BlKQhzC5KWlPko/+/PJ/Kbd1wYdD9nBJi1tSpjOsp
zkr7qqFFovGRjn5eZ6LmzJ68fFP1qv9fsxrWxXjCEMIF9HHt9skIRvMuosnyVwX5
zxfrZkNAHwoK0inB5JIvbpoG1GZQ6bwWcoEAlUvDHiMJZPRDvfz3fzWX2pxnDDvN
txGO3BicG8e+tC0+G8qtzOwfLG8AVRgdw793609zd4XuOGFnONEvYgIxdjT2oCwU
3qY91dBBjTcQVQX+ISEKDXDDfxcUcTHgwjoFZ1iAPAqBbN/iEzT+SNgKJo/uwTjL
ThjZfAprPUJi9YG9QdtNamwr3II4HiXweIpjlEWkxZJ/2qx5IrrZhC9NvceCgR2f
YgcL45yZJ2lgNnZhba8GL8+85WcYXIDJUvxgi78yzUzZn3OPB225897WPkZixpJN
Z1qh7Pvgvmzf4fsJEBkzPOyguJ0BpwgSd5rJH6Cybgx4NrV0o6EmZ1LQ4CAeizMI
AHdWvpCQjOZgUAmtoVkSdTxdPNDEL/fffYnmbR+0aKGb3Pwo7KJeLQJPiXwLIoBX
emZcPsUzhhbCPf99qYKGI/6aeKqiFRxNJ4oXUqchn42NDX5dIldAkt/4wNP+ENrd
zme0jffPD9tqdYw/0h/2MEXRKxfrY8CiavQKgWE51EJSRjJ9goGtaWGaAPChlo8J
pClGExE90Iyp3DnkFD76q0qgU/7DvlfZkS6c5Xk3S3m54AbuzEbQEPSNIYJmsI9Y
zdAtKJrx+dWkL8+lELCa2BY+Xl8ELLMBmiufhzli0ENqsiJIEVLks+qic1qWxylT
ymhers93L28t5UkAz1l/LFVfIml+/PAXm2HD2vsVcJUsWQQSXyHTaVJWFOVTzeeo
kqt0JpG+4mcVWYFLCypQA/tjsX9Wsq9fahIY2HgtenOkEOyX37CgVVsDdezYxdYr
6vf3Z8TqG3k0h8A2y2xzVYzVoRQhgCMuG27HWmTKVA6fVUjBYoB/yEZuF99rLxZ2
bKZs9OaOwqHCl1QpzJu2BgMdUeU1yQ9srqKFfB5waKx6GRK7Aa0esjV4XL72QLyV
FFnUz5lvaoxJvAgAF2kaCywh+PPRqhDcVPjbkahhA3RrYnq7cfIwBdx5S1aBM/9S
RijotQQpi1wzKhjdymSmdZ9j38mR9z4wfF9bGWJORIsNSRAc9jDMuFzaEnPbE5lA
deIGq5vALOcrrQbnPTmSFYdMDVk3CXsITT3H5rTIa+GK3qeF6gJsqKUR+oJVybhx
d9kmEoRlkqUcjpH4L2hJRg7RmVa5kMbANr0BDT2qxRqCk+8KTU2NW+lrTe+AIerR
xkRMGPtCXVse+iEWsyqXORA3tbHbCAgGX7VBwSWwMH/IZYKVjfrE1MQtmtLXy9wM
+px9Z8uQ24v9ovX3L2EBF8lCLkLsG+3KweqzABX6Wy7XF9bO+eq4BLjh1scmhedG
Ps2U3OUGT3WBRg4rB7tBoHpVps/LAjK8YHIp/2k9KL7ABkoveNqixZXggYHouvIY
Jeo/HD1u2bvkY2rF1gVGM/E3IXvYFhFVZPGBjQmo7bP1lKFSuLquqLT6JXuIUvC8
5h355HhmbqUMuk0CbGhFNtTa24NWdB73X/pHPhRt6GogrFPWqaKFnh5fxGJbWekO
hpbNUktmr+Subz0/hvkyMUPSCh9ScxlAhQB0yFEF6U5dxEFYgyG8rEb7ezMLezlt
scmS7DeLYR6XEKWQB+pU3lc9mURDSqLuhqGmv18ZGedy4y98BLk2Cyju+AuYPYIB
J+ybSy9XoKIPOH6JOQXoKAY13vihS956BXyTxww8F9Ub+GALftCwEIegA/1uyT1b
8rMoSjULSR0xhmOOPXlAAzARJ//+f1s2Jv3XyOLwp6Nw1O+8tYbzQVDzAiNU25bg
PSWI57OoXNuBmrCsyiBR7sKr6gA2htP9uHOqtW7886/nUIre32FbG/J8/C189xoJ
U5D9K1ZGEc3fVeE0pgSQLDVKUmEBR8Tb+QwGryCV+lgsKDzg5ROZib62MOR9q0aF
W48+lWdWJKYPJwrCnqzVRgOygUF3AU7NihC49E/Y6TCN/CTUGpOP+fJc+GHxbkOo
nhGzW5qgQJcGU59hbivoFaGonCUn5RjyhYMWS2248gZyL/Qf5HW8y0ZyWR0QFqtT
nUWPHbuEyQSJa1quKRcJ0JjkUjlzc6JOdi0Kv9l0ueGd/aWIxRM6hA6MDfq5FvCh
97LNfGaFoQ3q98qPGvX/LP7eQMVpx2ShCQAgTiT63Ylyiz77EW8D4/uma4se0i9U
jqQWf2yHD4vF6AIYATAAIDsgXv2hEKUm02DhSapx5ohcBPHUPX3MZi08E6hhrNhu
DZk2M/CSWl+fuBRyhd8cv5qIfZouIPSBLoJ9O+kJEEeTI+SFGQDMw39gO0a6Ip/c
Esdlw570g3GPAzgTe7/7Nz7zJl3BAAfDjU27EMmAqMl0Cu15UP6MgcAlO9BQNxYp
PBZXXFYBah1Ab69r4c8L39gVyIvOswe7Oz+KQAueWjCTcspzrx2XuEz5kA4Ik22p
nbmKqa5LzddlUnQNRnEGH92aLupeFDxI0Guy2xgYJ72BJeemUOc7fBugBG5W7/Pl
vBdk2AjPMGc7sqGUIAqb51HdZrsZ1Pf+8vEmVQL0tREDyDbR2iUdJQXMUSPbYU7e
3EqWvjNiJiDnoZGfOdBkGQHEiG0DkTL2XkX0HcncHPuV9Q5aAdHhgmTXolJUhBq3
/6aPXHZwplZ8lcmxppHULBxexfFF85oep1HmPzTz9V4jfiHZym0tRtHpsIdW6yYu
oXvXUp/JKTiw72O8hbD0otz5Z5nyJz6BWSvEMOzBGZf13G0kZ3gnAQzR7rB/Z7Cr
1R+GtrxkSiw3FgiVhzliZhmpumaaXRvMFLcUklCfgU3NWv3Cyts8eTPdgU6R2fU0
QFJz2eZS3RJqUkPfXuy9vp5cgftETdhYl2fSJg8B8DP2JJI3KsqVQj2xlDKsRl3h
+1dhfy9ksuLRsMOXrvKrwc7a5vjp850RJNxln7CySpWV3TNYIFQ0glCxXYzz65Go
OwhBisA5fOTqu33GmAP1SYApSJT7p9IsR0q78VisrumADnwVOirXOxkC13pSoooN
IBusLx2puiwNBIFOUaAPz67g870QYceLd1PrZYu+YmpImXpG3GdkuueUnO5QDEUN
tsmbKxNswBxHqpyv1hayVFZDYMZODrfS6jgKWSCdHydAHZ/VD64mvKdEFBRwWwbF
pkPr3NG8jA1PtAYdYVMKtjzh69WgCo9czpZS107krye3e9XrttWGhY1pzrDmT1Q1
P5D2rHgvtUzKvAktJFVLdrlJP2CRus4hpROE+hAi+Nib4WOi6Nr+oaDDjuPGKFka
yDnR8K1K4mC0Ql5uUUjfY1YnoIZE7HOGswNw4Nbhj86tRwi8qh29IwoDAEfRG3+A
eo4X+YDSt9MOseiiOUqGEcB/fn+FUMldobsEEUcBio6zCrArmjul1Bh2bDwf1FoD
UP7tgCusB/SvmwdZ4jL8LbhV5mdurCkgbiZVfZXp0ognQLbvtcXsU+Fhw5m/lVv0
PUyjvSb3IUxQuCaO12D7tAYDBPvSOWiMzbBbGhmLbVxAzfdPtHVxAilbv/i9xZaG
3RVgBmPSaKvHiIP9kRWNifWed1gppdntPIMf6mHbzCz+4nKqKadVYZ5EpVGSh3hf
+EzphytkHMizTy++3a0+zDoFEvBxoernluWho10RNvO0m46rDBxVbQBIq0tONr14
shwsJq4lv9nnTLA0vmJa0UmFXJIDIKYGaxyQm/jRepXfk4G1IwOPhM2YkMAndwaJ
wqOc/0G1G5TolTSr3tlQxBtCElUrF+iMTvtpV6pqFufpQvFTmToZlj9g1EWnNjBX
iaeNAD8E65PMub3EJbD69j8MgZ1thsEbuuX6IGi2V2gEbdPFYScT3gqC+wn1tVL4
oTgZtzzmWVoPHc7GU9WAy6zy3xQBMh9YgrHbs1z5hNpXiqTFJME8nlUX2T/gYzkB
91ypRdIR+1vbNTw0bRYQIoEnoAr7/PV8MQp7gIZMbv7sgxVR3O/exH7yGDC6nCdZ
WzJbWrmha69cat1PKsB4Ek+h06pNNnFLYRQPCZc0cz8fRA02lTl4NjoTMEQlf7bZ
SoD3wlSms0erx4cSK9oYXpLaIHfygqBJon4VBKlIs6XdJOKL15G2LxUpae9w4Rvi
GIVIWMTPs5icJapGxSAya03Kk/Da+k1KAs5QQSy2bXDv+7Ir/knQMBAOK0MDyvu1
aHs0MM0jjNAUnjp3ixeVl61PiLrycr+ACwub4rgQjnQHxwT/8o64A/NWNSEsAHz5
WJkFQJrtcR20fVP3TPZACb2AisAphOxN2F6cg43GNQeT/5a+J5UmjCVE93WsLeR5
rASCTU5eTSadQ9/DMvBeLu2cXMyljgVdifcqqVorqSoThoLx+9T/1fWrMFRJPPfT
qNF4eSOogQTQWG6PJieO2oYF5NSZjKU4eHNaHf9cAY5z2QQUephOVlFcFgZ4qiiu
183vWYZUvEXHV1Id4pEJFF57t5pamI6h+fo8GRJA/rXlVCIVGg7yGi44eBKjMiVB
VF+66RYo53tofkdaUkxIXf980c6AmwJ70nyKjm66kccS0f187+1Mx09C9HHi1rbw
asMhYEMUW/MDVKcWWT0BAc+5p1EJfJlIoDalTchQbnkupjYw2NRyOUmfRSrmaEpp
wKXoBnrgfLj/LmC1m5QV2kc907XEk5acMJLOR/8LBBtSbDihRQ0Va2KjnH6maZWr
kPGhXyTVBZcLqYnZ/eeN4M0aFus6KmaRK1W09UUAQ9cmqWAkzXhvkT8x8OUfsDAU
fgk5zVaCeVKKpN7lxWbbVKL4N2ekmJyG/M707gH41UMy3eVVY18dZllZ6HQLoQVk
UmVLGtAfaaRXlnwFGtRmH8CewKQ5Sk3BSB3o2nfr+VpeIHNhWMmpmkUPdOMFzHF/
3KLuEYBd7iSOlhlgit+G4ymYGmWyWhxDMq6hiEw7qJ/+yLeTVNWqyc6R79LiGMKE
xwagoQh0uw6lYN/iYtIgrno6Q0SnC59EqLBqT+IOKmXG4de2U26fflnFZ+08TkTy
ZounOl/eAUeOfWN0sPPMX3zQvBzIDPBY6zi/+7X0HebwGxqqvGpe4Fkbg8dNFjav
sbvYJXLoEbS7A3+T4xpsX4nH+RBo0DvkAaa+fkqlK6ajTT6GLdprRMG/Iyx7Hju6
Pe/rL4B96lIrWC8q7t4C89UV5QpJ02G/L4hg5XjBwob3aCSjNvQTIkcfiYVvSk6D
+O6bh5kQ8k2oNwluFlE1do6jKVOt+SCXjj09BsWBbaCDYmyQqr0fiXEsuAWI+pds
jR6Uxv8oMbfywrgKqigNTsYM7GHrHORKhrd5NhaPNggoNDcY753hb9FcI6n3DlqS
Gw/NtaLzE7oFPseFsDwI3Hb7W479jtNRwI/iWkdgNBYhh6SkX/ZzSvw4Z7HJoecZ
6OblHygXVvvgFxw2a+nb+regszCR591dA6J/T5oZ0jQCSmZmVPNui9FLkn9QkvT/
FaxKRPwPowAwIwXbUfCaa/1rJKbgMH09NRdnUVNUROhgpqHmDdwv0oE+2wZOYUXJ
hMRAauLb8QB2kcgWQ5adJE4cRnqTFHYo4ffpfHv810pszObXw1VgiwmyhzVynzvD
W+i5rdPeOos4ZvhkMGRnVngo1chx7KRLErNp7kAH8mjuJgUWSmpG/M7L2bMeLszj
mEoQlehxP4soHZTRvUIoZ+0B9+V4WHZ1LaoRM4RWQotzQXpcEqVl9m3//9FVatJ3
hwnNPapzTw/migp6ImnRcBGtL1gJIvAXzwmX9Qe6BpG/3wZ9Y1UofIR4ccr4+dlU
cQVByc0ELAPsBoSh/CKBOjNmGY1P2DzN7Q8puHLxknlW0gJwLHT90SfG/9bBuXkh
3OumK+45fMQJnrjyAI8i455M3MlgMCKEz19fGRlgiPnyh04cuWdshSvQf3Y2ZP/j
DXsYEbPFdBQ7vZuGW516E1F3M5kLZD6/RkZmnUTN7FE0xMcc7S4CH0C6fG2oy8w1
GgNmKfZjSbq1B+GNC35MSOGTii7+SPBziiwuIphmDrcgBWPCPgKNkTvoGUvDdBy7
uZfIdF6NHV82Tju6sNSf57tsMWmaWXZly07HMV0rCKb6Lxu4o2CteXqhERFVsQ6y
wGiz+6dPNebQ81XleQyinGz9Qsbl5ysT8MKkCShedhrgBI4WbQ3iL2eh004B6r6i
hvAcg+PZCl/bBSvmEy67h8cOlrBTtdDe42Ful93D0CBshQWH/kDLEI6aX0oOhtK6
I1uv1vNBQc0/PeWcRZn/G+0LGBLtwLc/tXcijTcMlQZuoCoLxsBCJCXu1WU32n6g
lUSUMm75sSxjlUW7rHOeznKQZaJ9tlQdNWyZD4+fAsqfF6X5MdXfbk9BP9rJOeAb
bYSRqDjDXsPmerOosV80IVdfT2hG6QVEwfX7v1iwQIaKmPIWDk37LDxU7KazPLJ4
PwpWK0mAQe1K9fUR4Rw9fulmTU/2HUVyqbfLW9c1+nVRsBIxCmipsg9CPkWNTd8K
f8OGY7/Sfq6gc2chHEZVIr4X5vtpq465kP7GbmXjK/5g88vCHDCAhcLzMuqL45AN
SsEaaNh0Y5RDJfY43Rl5MISpZU26iSlN/OGW2xo4XY5FVhY7duJef0BUpTDneALR
f1Rt2BqSR1r+CWgNRKcRUJRKomtApEthZ449+vgjcoXktSI3EDsP+CxLV1edfrlO
FaSOwfsZY8kZYg30diDRlfT5BAHMvaEVkMJXVI0QmnU9imMNjtzFJB7SweEPBYDu
+1+ZSPmxsQXgH9wtJVM22n4eOKl0gjAH89HlwTIY2MXGOS1aMM2yBQWRV2c3Yjyx
J7TvH8d2oz+bmA9UKmBGsWVchacr4gSPXWQhui1psvnjZPQVPZXfPg6bV5UVIL4G
HWXrdjdo19rQCu8ADDBwCXjVouJrwdaYllf8n4ezpOvALRZQd7Dc4LlIQciKLqD7
XFY86YZN5f+m09IpSChJYqbuxtHUYV9C/iUZnxPgBGLYsVfomOpDX+yWnt6vbl6q
Nw3/kq8bB98Dfthy/wD4h4nVjvLhv52aGEJwYk9IC0ac/UFy6WDOF3ghLBX1uddl
QEShr2Wii26WoG30j/hNmzAOLnq0iWKRa0XiF/euwLGUsIPNBc/w3F20QYjHdVgb
2mMVlnVyhYd8mxoxZJN7jmkRdbLWXKYRj6a8rFbLHJWecNbLXRNXjCKd1fccNCdL
EjULtUM6Yz4vgKO6N8l5i6TkqYiWAD/QuG9OVgKkIZUZFpEUvHbCQiNJSwDEkEu5
QzuvyjD7G6qxPlEk+jxDqxe6XijytkG94it843WXHDTCsVsuxKnU5l0LExKz3zz2
Ug3V7GaocY0KVuWdf/Qs/Dr9mn0bF/bsLoN99yZRc9vDmqoj/ThLdC1e2vfG+buX
r4GRcYMP1uGHSWIttFzBc40YogSCierTM4cJcgwZKsnwigLXRkmGDT9v5uGx7O5o
DzLhvBPl5RBpgYzPBhOk7+azuLLI8A6i+yHwyw811tVJv8RiB4JtsZbcphhdqSDK
b33LLZb234HEzzHBsZBawIgPTy7j8y3Fj9zFCwb6RDnl4dtbcCIgTewp4U7Qwxd3
8Y5mtswQmXH68wW2Fa1XcNB6FnAcYzl2X9H2SyVQq0a9UyYGnJ/Dtv7aaRkl3Chf
QWJ/RPhLF179aRVbR6K9XxWL2Tpb7jT7AakIaKoRtgwZ59xZMEEF16x3QXXO/Y6y
V2Y3rWahsN1dJHDyCdTb6PotHvwfLgYh0tq5T3fGbMRLGUYtTOh61CgbM9Dmg3Q2
WFEE6tvrahTuyLkiROfijLFUlkmDBdUR7kqEDWNj6kUw7Cp8rfPoZxr6/HINkNWu
If+DGiPYqazUwH6cfiKKALvvb50zM3iALVS2+nIX+fKDj66hyM6+pMdGMZ4lf7YN
vW7z5b9QZv/nAAKZ/SNZ+3MHx75uUC8ajY9T6n9jAXYv1G8/AcXsXwu7KFVpSD6W
JMFERHAfAUojwNJaHv7pUB/pEVfZjlVf35lwve4qSBOKcVIGjOgilEDeXFGpK0qB
8U9N8HpRcJJsECii/SdSUYkSFp7OI2LWE+Od4QKxRfygERvagy1vYJrd+PAd00UG
8ydgpIweRgnSB20/kn9ram75JXhBrjGSq8d3n5+LbghzNRdnrq+9L0YfMyBDLhzn
YDx+6+R0zRQPuAbdy+eMqa5BZ7liMcODWStZF4HImWMIK1Rfe/IG+31i6znS/GUu
IhWI6FNwb1ud9ZN8iHKbcYRE8oPER0dkrVOa4DJBIVgSPy0dDEw0nsG/MoWjliqx
zmARO/nb/hqVtfcFBjjTfgjgiWtIOnQWHuWzPonaGIkwn7yCCw1oh5ZwUvLw2RNj
kp9CEJZHD3P8fCPnTMigTQFYegya3mXtB4/PSbGQx/Erb0Rk60pgRjGVrwNfHwRL
Nose7lOCcj1ySraWaZNHvHgifEki7Rusaj3Zk3kJNsrmQu/P2xocOeunK1jhTxkG
GXHxcgxc9T9kiHi/jYPd4weYWXUOYjJdI+at0gIDUNqrGXpumxfiGYL4/nr0d+fS
Tj1kBM0jIMz1HbDKbJQUr/lCWMU83iqeXbfQLI4/x2S3V1xkoRemmkjNDKxAaAX3
BQuSGSAYvHikMqZFFz4hczz64MTZ0lAbYb1+lkNa3OvZeNypR5GMEunRt5ng+Yxf
D9XrfUlW6ol9tQyHHrBmKPn6dOy+IWTfdAUBBXwqvoRwlOiXeCiG8T0ezK/ZA8lY
dYl17lTsfQBYZNaXNmII4fkrsQlrSKhovU9YTBhZ4/XCPEDqGBSbnsFN7glZvyXQ
9YE38W80HCH+NIVJRHstLAoXMrkhZfDBl63m816TPjh7dLg4WSaN1P+nxvCS7Mw3
PeqDIdBznMF23lHkoyTZRKQ1qwVWwXR45+clHtkn1dE8HDikLTT72NH28iwE4Y0u
pQg9ejzEDDsVB/BcneNj8Gqk2imfRr2fZhdhzVN762NQ5AEX5njrFnTCUDnWCrW4
sbIWu9TpkbBM+a6+xme3kDb5v94eQ7A3qk4SiHhRl7xo0t9WLOdwoPtT2hVqZTlm
9h6YcCGBp/QRvXSfHmcwwf61u/GHWfNUDz7dnbJUG5fdhncHsrYa8Vsw9MCbewI1
k6lhMDTc2p7/yMk6e5dZlJfCapKiDRZH0RBj15rrv0H9oLcZCOIdc1IfS9fH3Txv
QwQ6hc77LWbhA82lDLNk0J1sqQTrFoRaI6q4PSgLVJnqyu/My4x3FUbgm3Appwxy
cGHjbNseZLBQmemVB1vaNboJezKQktUdfd2hPX5jb0cZ0TmExkGPDBgatS5ze5Lt
nZR/YPvYwoPj5GKWmBh0NHGz1kcKoYcN9Wajwwy6jp1MVMOuhOazilW3Xu1+zuUa
Beh0g8GtHZXY2jZXTQy86fwcq1A87YY+ckO4prEK4wDsNcXXbgHLGTPIvyJN/Hmi
0EzX7YcZoXNbkFNVj6JA3zl1Md5PplNa7wZNjglT32hpFL8MCRvaCzamJzcXJqtE
xKpyNiYMBuwq2b3S6Cs/FkrLrPjIsKdmdf408BzthTYM8y0emjSw7hkum50QylYU
odPW4xGXwTDXwvt7UIlghCN/xouCk/tbNSHUW8d4BY686IaaTaXR5qFBcFQH7jwi
MjapFg19i7eU8K8GuSTi2TEvlHOCEMLDxWP5x5Vw59L+6wUsE/p6NXy2RpCnsLa/
WflWzrLzEc7su1fbQ9zYwqkbHPXFcFB41bvFJJJ5P873FmGj6SqHXB/EF3HIICjt
4Agl8CGgm/eln2DFd6uKUeramAJgJXq/ovsP+yWc5sR+d31Z0EvI7w/YfddxwZie
4eS2phUon4SZBhpHm1xFjVt0loYo0Ye7LhO/lSaislQW4MT8UU7kYg8IGkV/zAjA
E1D2y8cuquDXwSuMZJXXwE1Pw0MyOarPIO2mJgXgGGJe8B5jwnj2J6moqlYfC2QH
srYQVS+QlCtJ+x5+QcXQ10QJ7qCWwMw6EAoG9nsGyPYPbVENDxkE5Fx5lZaZiXB6
gdl43iP8+j0lLZGktii7zJG/3BBgBgdndt1f45k4faXBwZnlGlR+XERZaTuXxkp0
SvLVoeUXlXgCAqcnRsakCu2fr0e2Z74fUdF8zOAMSSg9cwGUyNOtV7gE7ls06peN
SxDeKAlWQN7Ucf0juHnqAIXEAtWF0o/jRAyDY3Xziiw46EYZzt4UiqiTiLFYmI+J
ukpx9KfL3o3yeTAxhT6Hz6JLt9iPDqMRlgmUAb4il3E/1BPSRGksfaqgAuwtbtIq
oxMpsXUyJfcTRJ3VexGVdMGq/clDoWQdZj77k+F+nQaDmgjkfbtiv463hsyjcokk
CYIUeaLeyXalA9p+DEu9RxikMjPoJvdHW4W2hdIhYAUxU1K/OCLE/pc+Q7GoGGa5
sKWomkHYYGgQtq5wQeYpoEcaB5RiOncvQLFFSciF8CkrccXOjN4e1rNIll6kXM+v
rrSmat70c5aSP2j1Qxb/wtY9VFRn8CnWtDHnwsLk5FbJBlKO7+7RJOiELAOdnwcQ
KMW/5Eyam6Drqw60aH1gXhJ0eTzCfWZX62A53bWvnGxW0yu1OxRYuEi7A7JB/evx
PNnFhF3PHcaEq4yYyEpzE7SHIk/8xDtsgKszuoPDjF+63xEB+mMWN1tjAW0ZD8Kr
RNVOZB2W+KHLoVoRIX/T3881yFI7BiZBWOCzmzKjk3yMV2Z+IbYsPM0uHQkuOnLf
q3g/st0jg3s5kpo2v8Dtw7kue7YcrMSQIhYLLMllX48eIM5u+FG6iTRj1F5EumgR
aPA8+wcbycMUzUM6oP9L8pNsBXRWBamRPXXDbQMBi0MAhi5Lj4gZSvBWzjO0PZQd
MTKeqivPoGVbu5Bh1lI1ZhVRbgtMnlHBUvl9Ff+2nvetonRrrDem/xpS4blmDwcS
cFz28feM69DFElEX6w8v4dDTV7BYjK1x0q9m6uyR3nQMLvg+fsv1J60xkXc+sN2z
EfFHRz3xV4tJoZSxVahv3Kqh+/JKYWfsQzZ5uSi8YayZ8fTUqBPxSzr53/ACkYZZ
AZymNik1G3K4B5ViIaE8HQRdPWXUlgdXlMSKZV3w0gwQuYzt1urU5vvzVLXvZYp/
GVNNorJH2KQpR8NFVymKMWuEmLHWb9G15O1wluKrxiIpcO+ZIc7WO0Mg1F4VxUDh
pZSUOnT4skEJSYskMMW4eSEQTQ3z6cvMh5YzPE3RYwIRSlOKiRbkVVvcWzzksVXX
EmHJKs5g5ivI0Bbjel1X9brKT0WMiZXGXnr0+YU9uSQeQ+BMnY6jpgeU2WSLV0Hd
jO9qov/hdeFuTr8mcff+YuWgKtVwEl9x92g16IQ/s6b6a8pqg5//rqmDbvEmhqvL
/8PzuVMs/MrxylnQ9C/8O5uizJsjmvRn+Dr7LhojTSvQMrY9htTauHa/Wcmx0rjo
2VctlLgwCxa776JJKrART82XLnegfVlKzW3vuZdrhtSjo8KjCFzzsmZIC7XrxoOQ
NanAU1HXZSGhlJtcSmzv3P5FYbPugg6p5tQAJv+/noKs2fFPTDSqvJSVNeusFI3O
/GmEY+YNrLq+5n2xru4KBctef38StRjgCryuMoA2ZwbVhNvSix2yO2IsTlS07d82
qr7ILsjcLwpC5Mazz3KZKg0CBG+vqzmE8Bl06Ewj3+gxMkgOWIXirH8LrV+Xfcjr
NzQmIOpaJ9HiTTX5GOqz3zPk5xmbNhIh6HBZbqcjcliXYsLo+e5viB97N259voNR
J3y78MDMRVFZ3RoZtlKXuyrDS6KIJTEEaQbi0sLIjP1OC4h3JS/AVRK3fwn+ibvp
SsqtHLo7TgIAnkk90htJKn+gyu9JxMKZYHTEVl/QdXxR73657d4nvuPGj2DWeO4S
MYVTRCpXPIhaqj5apx8GS+IsoJsj6NHRwvU3+KvHsCHITXkurZFiZgI0EAGPvpbw
Ud2xRkuFK4Vkk0WkAm14mhdCqGd4NbhbcD2oVGoPHmRamacvYvfU3h8v94gDmFJi
GjzfsfBF/gnHyK2ZfFbsvPGBCPMF2CNwtKCexusVbvGuM5OC75R/+MbKWuA2oYdI
ffKmXycn4o0A9DpgnGENEkjzuZ7SBlvMD3zXcOAeKH0vqU75tZZE6ACg7aLzY2//
WNwL2EikYZwkekKsyIiFi5JQSGLVmlRimfEkkvRPKQHgWyaghYF8iDyGDY5Gf2Uv
l2d3JpNsFxHgxE+WUNakdgbzB/UEU28OP470+WHbGYPuGdaVFo4sUpfKWViFZJNB
h2FupWFvsbbCJA/ffnzP/sz55r1L6OiYawY2qhflJvCXebjyzdYkCaMhp5rkNY1l
akTjB6XHIu3SX3HLT5T/Uzp/rivmbKVXnFxYqhzhMSqIXn07KDqVpy3d1T57FTAj
XLZRu7rUsrCbLnnZXLSrQxZReMUnjU5jc0O4m7OznKGRnQ3Jz+6dnG8JHSHY2EfN
jOFj9uxK3ORe41vNwCxKE31e2Z01kfzGzB5FzP22V3xWaGbZKgXWfFAMn+Jw3J40
XoiQxTJG2U/tWiKfdcNLUC3j9V1nRzrNgGPSod/kvnR9owbqlTTIcJk0+yGfD32H
GltVezf/+iqNs76vY3gdHN0ic1i4jK/Qd6KvOOX82vSKfqbxXeTvmrjKwkWbaPWd
lDtfkjwHxNjjy7XK+8S4Qw4CCZV/DijCKjNhiomdZwg4ZzXSxH5OMexsUPqloMPd
Y3+l3GmuNzMrfp5KZiUOB45rFFzY6RGuoKnJ1MjzFbfIPZu37UJoIdG++aM0ZExN
SXu8AmvtP/7pfkF9baQOBQJ3kF6U6DB7s1e4s3APkemQh8a50DeZCVreGh1CQNaG
n8V9tY/ktX/zarIqV3yEZhgDruV0A/Rw8PNNSP0sulscicTHxizj0U9s+EqjO6gq
S6iqR5S9CHV5mzxBdWENgCciGyzg1SkL8/ZBqp87A38siz/Z/YZUqGesmBCMR9Dg
ITxUEheQ8YYDsQ/UKH2OVE5exGMcUgE8dpGGfiLFbsDmOaEXllcjHxV8ID6zVtKj
xVMI8Jtj+5sWPI2jBvl20L1SPxdbkICIqjSrp9DYz3kGcArmGuOEJeEcPf7398jT
zA7M2HxIgcSBdoKxMGCUGf50UAJfObuApgJrJ+6TfR8s8oUD5OumCufWRY6zLjFB
in/mlzq5tQ5v+9++bB5GR07Ytr12Q8vikmMkoy3BmIeD2IJ3E4aM2HHKqb9KESlW
qrlnZXcRXaB4KXHMYgyHQSj3SUiY/QfLH98cfJeuMhgjYRdt9BwHbotG5kyLB3rL
BplN9IrjwWuplUYm2vNRWccWv5GvPDwABv/VA3qvDF5w/T6abRuxkgEnYCvThkD3
aAuQt0JJhxbk6B4Pu7oSh8rCIAV2nb9U14HMrjNSmB8hqguINZT6oKOIiIwZEkpg
sudCzB89ab1PuDElYcsvWHTbFI+zXk6yMl85OutS5ja4SaBARvlHDcVU0XE3xg6O
LZbjhAAoEgOafcAtSXtjCrjfyEdB7tHhJetlGspBCOtLl1fy8I14FUyeRyJcVTGH
Zl0+rh/wki/syDN0TBctzgIPYvsrGbRvV3kpTeD/0Bo6QVG8YcSOn4ZGEo/JLs6X
ymI9ogTsPTb/BTmduHgnmWV7QPNB4w4Pt7D0f0mYWf6msTSBBbQe1LYwafXmSgWf
t9I+7W9hxyqxVmY33r63Oem5IbVH9lovFZDAoznaj4tkByUVvyni+EC02lv5HIx7
O7mb3e0yN8eizCV4Qi2O1tgqZZRwi9YYCnLs3oa92rvgZCw5qGaeCp9dQkoQeSjy
AuykCfLl+ZRA51e89jFLko/bGSpwe4FXi8iS/MsJd17FhtdLpDadnZWh08aksmMn
yUlL6XBjDk7W4SHMjzV+TS6DgoSAOp676jJ6gNct08Oe0rIJFUVxU5317UMGIWq/
V2G1No/fQCoeizfys4jd6tMFwU6OMPcATqXr0C+0W/Rd6L6YCq2zGqtG1b0cN8Zu
5h+vvsV+b+xOnrhRcILve2FNf0iRN+sfCk+JGtYISnakfZcgu3aoTepwLXC7f7jX
VbhkefCY9ckB9Gbi3Lk68QXe3aYfDTsv8v1ILfD9xfDO2cjmCIIQLtqQsgSZO7gL
FzGdarItO5wR0CeVSbHaQhXwXkX3FVg3DVr3XO86+D9rLyIWrfgC0+6gxQyrk90u
0co3lsyxmApIgKSA0goAz1KQBibbhFINRX9wAotwVJD7TT4QGVnwRZ78YoUwB9bH
UcQwLktJMXQ1khopyLIOwLaNsqR0ng5NT9hMpZ1ivhUNsYCOXqwqL+Vuic6DKczl
YkxCu6jHJwgw0u+IF19G56tLccNU3UDQ/4Rk7i5kIqb9pNbQ5G3/7Dfsv1NrmyCR
IGMHPD5K49+w+1FF52m5RFNLjsl1TiHQYDo/50lPXqVQkKZ/A3jy3CrLiOTVY6hz
zv3CTGcCyUBjpq0r7SxmpNTxltmOyPJb5Yw8ZZhAQmzVLh1CJ5qJQ8mweEgkD2Vg
NkYu2IEVHKBmc1XTsJFswhrjGcjTH+5L034WXR/xRZE3vVSDY5yuYPQWT0wDpXfe
YkUmIHvKqgmtvEK3KGKq37OH+kC0piTolOeX6J77AhJj8dNznzG/1HjODTZ+57uV
Xkxh4ul1Ndtf3UTzUeFKX+GPtFZDkuXWWomrSvzsJiAwxbelBbSTrieynomS3wO0
v0hGeLG+6d0gb2Dv0HHv/MVoB3bUtJMM7m4AboHYwwuj9ef1/cWJg0ynUmXVNzgr
6NUBhAasigEf2R/cDEa4hXWkfNlOxahORoCZ3PFNkGJkCUs/y0TwG8WIylXQiDZy
ZHgxpBQNaSmGE7Fl8XMe6dejGIewG3ao/ifucdc6Olf1hODk/MoMIc+ME7b06Li4
TqUJ4av3+t0F8zEMgDEdO6bXuCI1mIGjBLzsjZKhk1Js/BcemIZpFTHejOcpZzU6
AslTf5ASmrH/dmZa/OSdwby1R7KHkG8T1VNkhjczmKA4L0uvByukr94C5/h2Y+ko
erluDIFNjWHoPyiQ/FYtXvo4rbckLsEptZ9BBYkteFDGbUFHbeIKBoo62VkOlfwA
FbNu1wNi50D0K/QOMbYwWXApS8+b8eMPea1bdFcgosOhTw/s1xA+j4BkKaT/wUjN
ec9C1SmAN52LppQ/WtMPyDs9TiJuCIVkGsjZuBiEG+22MbsOZNkBJnsDFWreOhgg
3550AbeiIOZchmHgUEb0DveErP8qR6ZM6LtdAyq+eLYpyIb41xabzPzOPhPjvjTB
HEEKu1qfxqd5qhMH7sUrij3K7JcYhFLp/hBBuZ+5GBA99xA8vgnr6ukPalTiPnhB
aIhTwBy2cKIaG2WgHlWQ8ou/fbRCfG00qxhr/8/hUfLLC93uJe86Wno9qapMrnP9
X24l3VWE+rPfxi6ON/cPV/cqsgLyTsqAbwicOz6EMBJ4sM7a5R0e6xcZvwbUAWga
O+PzIn79iYuGhL0RE390xWbYkv0QnPkaRgIMh4oOgKeg/fjrJG7LRHJJvRyH7PaB
OkdOYRP76BMih6e90PCVafZD6jlt87ybgYdkBLEzQaCeYOVzhZGg1uGajPS1NN9r
Dl8qs5W0A2JPX6VbEg4g84oHkq/bC8Lbf+LJOVFb14ptlJOgEzl1PFbkgLaCLQd+
ZQl3q61u/882CMbN8n/CR+v2hfKCd0lwiyx9jn3V+Lfl4SG4QFmqrnkZ1M4xFUmQ
Q9ftQtivvv+8U+tCxKUWG2/iEj3JmCQdBt7waGAR196lpaRS3F0WjLZtZkauu9lh
ZbKxjD2tTPIr4R8NUsVRxILqLQVbrdICfIGzVaBH4Ms/Ody7MFjPDvPE3zmMPycu
kQBASGvwQeg3+z806eaLJRWLPN9XH9BXhNx792ONZe7Njfx0dEuGM6KDLDEyvjVx
CUmhxs3uOTzty5sLpinUDVTGRCzIsa6PhoRoa89fkEKhaD86Txnh5BYOTP1cx7OE
MfTOziyMVYZPLcvDOEMPrOhqVWr/HfMaHN1Q0CsbznlNZprKHq1bgjGOpzGmYMkb
PoYXToPS1d4Q/QhNNdNeD3AZar1GBcVURYcgDaz1NzZ0Q+w9F30TyNGKr7gcc0tj
Bd1Od+HJ7Uj57xkKfoZsiQfPieW4v9BWlDzq97qz98k3+TDYyqhAApJpbH4C2+Nd
Nz7fWKqSd9bczD+n2q7qcSFG51+7vqx4TLDpHtzfbR8WcafQx1oCGGDmfyVj9Xwz
nXUmk/GrmIQIdbSAMlTE86xazQ/3C7PBYnzqg5eZiuGWu9OszGzxFHy+MbgjkV50
Sz6xKbXHZ4kkLqNtuasn5LKSGzEFy8qx1V/f8IjQbJ2sTPaJu3DaeyF5GfzOq+wG
aVxsu381hKepPd15Bjwc5S+adXKRbcNlzMJXyDIkLsCgI/pu/vPydJo7q3dg2IwG
0Sb053DaagfRvJBJfFVRygBWV3/WAa8u5UvoAL41gxdypfJNJyZsGBB2UzZjL5+t
l0Foke/gWthyOR0b7qvVOtIDh1WZUg7X7dzpNEwAad2kjpHT97qyfB7s44lnR9Tc
AKyej8E/diKMimY+6oW/+QRtE4miRXsBJgyEz84A6lM6OpNYAyPXbiHMxuT+fV8p
YH9R98zmgD/MibSRSBBBJmTb3AYZ4YWTWM/gs419mh7LotVIQYzslJlWDBgm9lCA
0v21Z8/L09CzeqQhei0OB9k5eJe7p5x+pfIPkX7ooE4fHwfCZBHrvclnHieg0uyT
GRbMwsRF+7T4bIXRRNhi8wm60Z9YGPUSVXpjW6oOEJCkWJpyzhDep7WirMzZPGVt
XGUJ7ekStQWufk/i/4HosdrfEhetCOd5UVRaLjkIRacPpARqQ7ZKj1Vw6ehKrVph
O5pcngwiRsLpGdA6TdYFlO0rIWMa591AZq3P45W/xE7N20scBdlmIdqqGZox+s5Z
wfwqLgUZ1poxH1ss6Gts9E5WyfzcwX3XRnuF5+BSqJodcmuKW5YqTgBgr89er12S
GqJcLM+2MInxG5+xtngVPuX7NxqSkGEczFccpsu9SloCUqsM5n7/Jglej1C0P2eB
cvHRO9QdYmYqr57WgrzZmyQ9vmrHoqXXnIJRmv4VRKgWlWIGg2DV4UarFfkN4yNk
3xms9x4EzYcg5OXzzv7z+kWhta0OGGVR6q6j3F6WF7ZyPs1OxcxDUs1+a4nToRgp
3oOiwldkEicu297y9XfdSFZTILU7YqOAgtJqI3Jp0SvWAmJXWREPV02JkdlpDxS8
+DJ/s67kf3elin1CK7c4BwEGCVkEGRxqaLDOBuJDRQ66Mv8k7+1NgzGKd9dRc3xx
3go2e0qx0AMumF1UvDqytTgvgjmrsMgBUnbz93vi3pjWAtcWl9K3IQU81aRa7iCG
BxVLJVLR6Tl1tbVYGH3wuu/UU1Cho20j/RLPPvKCc2d/fa3PHNQTVuJiw8V9+9Yc
FMblJOyC4trBY5P0OyzDBtow1e+KqGE3j8MNHwXfPzHuxiXh0KMrgOLE78JQDBAo
gt8TkA88UJuvZ9qNK5oJeFZ2fwLV+nr2469VebDtclxRqPW7+WS3aF0E1DIVSNpF
/CQX9JK4TO7tZ+Fr6nE7Xqg7ZJ9PmudNhgUnQ4IflQ8DtoxkRwUruChTPHvgkHRE
7baY2/0INTW5zT35LdR/CqJW/RAVeEGZEXMl2byQaPKDJvHoUbFt1E4blur2Q6gY
5RN5uaIAFObJxGTZksPceW/dmyYN+IEJRM7GhTR9bkItu5w6ZcXUoWUGHKHcWh+k
8RuBYP7X4l/15floU8kthzZD9vbzEOl5exXpo2MR80GPGOfI9sOz3cWVhoaIt/rP
vnlZG8RJvMyjPDqc5s4WEO48fgCmfFOdbMdQS3aCu9DT3gUq4gkRTKc1MhBZ1tKu
Kf9AruCob3H2x0qepjxI4f54il/agCk+YqRb1W5Cu7I9hWrfO1XTuzjXizdJjLi0
CirdGJ652UeywLRKpQHjhfs+BiHaWgfoVmeuyjmJM8d+r13ad/28RTTB+O+Wv3QE
UjdNk67bimnPSH7KlRROhXXX0YLFfMqMeAWR7gl/U5SIUiA7U3z7e+Bm1P7h9y2A
rMJvTNMKMXhOT9bn9yjgx1PbOmgNyVljXOyUj3AGIwwp78glVYiZ4GaEBLBT85GD
v3D8x4qX4SHZQgJBDCLriE9biNvFF+ICOY20IGMEcYJZeBsea1IzePpe8TsuMdjd
lrWDtUwflMa4gBl17ui8pLC9c/dG9rTiisBZxdA4P/bUHE80XmlINwsS/+Mo1RJg
QDcipkLr9CeAJ+u1E+qVkzSMfv/yerHPV3KVpQbMJsW+2BLyrALNc7oZwxO5VkOf
ZGWruO1//x3XETIF8/f6UfzAUp2/k/ipKYy5KZC+YBGw4a2xMRkrsFzCj/CdK5vu
LKVuksJu/KoKi1k0owGMH/poh+O8UeMf1nkQ0dWP4VxmDDCU/IzqPPRHimx5eIfC
V9R6jiBDXI5utpx+q8q+Vm8IyAS4Rd0W9XO6hS9SBh3dG6LGPGupu3pc0mr5Y4ya
7ZROu2kmBd28PiMs1BXkXlYMG3mVvHUn2cQM9KucbG2rpHlxdoc18Q91KVeEZu1K
m9NPuLRxSHOQTNZ7pTuAA8GjpymapyfF1euXLb+ptpkjbro7r7wjuKcPjf5Jsd7K
/NcHQDlaQBqGwt4xj/5X3paDnoKSKnhqsB9WXcMrIac+sd+klqPtoz3m8GeIRtmD
j9JXRLmUfL4VXU+jK0X3s7h6AyqG5lJ2gRsH/NZ0+9byQLj6AX1e3e2OVmh7ftZ4
8FXLgL0ENnAkpBsPo7CqrTn/snGTLEwdobvt9dvJhKBXvEUJFyvMVmwe+XEgoQtz
hwPJtb4JvvhQehDud3kEWrvNScfVC0GWWMYFiD6sjk4NEuNC+mG+UQVaOocVddG5
gSM8sMeMJz9/omQUwhH1WVIoWl0/A1yRLuyLpK8d45g38slJ/xok4/dWV1Kfdx3+
u1/BzZgqGbYCcnvOSjSV5mHAiXK0/RmfiCRqL0k8TLY6WeYBW6EB0BY3Tzt0dlkz
22Wv3eJJ+UZLsK2CoNHO67B+5Rf+KJJBwNA9Npjm9sm442PP1PuytLPwsMi5BRK7
3lzfiS7V8ck4kG2D0c4dWjoHJc9wgEaIErIxqXwjG2fqJO/CsPi6Mj72Ov9XpHOF
tZCjljfLoOQNWW1fBR9aKPrdD53SBqVx6bjs/J9hSiCQTzUVL3HVmxbXok1UNJDt
SPIWjP6T4lNMehduH8EFTwv7RXwVKAvWNDJq9ztDfAxqJkRIgYHCDxJKcwitH7tq
oaSMOtV59LAhiAR1cTkdM/aePcdFUhMHPmLcbOz7f+HRo3gdUICpywCzAq5FdoOq
RwSQATJZgtLF0W3HL2cpq6bUYvk9ZDQBkzCGD1Ra7i5XGZD+zILowS4xwyElprUU
6ZxtOQeXKMjgMrLqMBE98P0U3osRVGYU71EQdGJyChhPofqjCxc+DgmVmppmv8H4
9cnYgieLOmVuYHO/45txc58KRdPO4HYRmO3kJUxJEenrXeAfln1jIvQJtKYkBVxf
gU6fOfW2hO99zzzA/suTukfm9VykU4p+U6qfi2oxbVndgu4YYH+VBpdSK5KHskcU
JeYlIxu3c8oYyNOZ69jV/9w48ejx85dJLo/AC+dfYmxIk5SzEErdkGQpsqi6bZBl
a5kNSW7o2rpaTh3WBgJYMCp1OpNJYAcvN/2pgeEpg9XhSfQPw1TZSzXLjqhyxyrR
jQgczuWy1LP5ZzNcywRAehfTT8MM/m5Z5iw4Kblw83yEz9qG8kJFWAE9Lq/nODla
hTQR11JFmHErJKcHTzpQ8IbjpJV/zdikyEgsJfT8lvjCqcif/ipgaj6DeBPj6NvX
Ow9BGV46pd9CtpUsyW64Fou5nuBKKuVvAwAany5ZGmOz28zbcnwX0t7ODX/5A6X5
CkHHkU8BmLw1Nv0BCV27y7vMaf/oR1W5TH2MXS8WYObtIxhQ4HoRUZttyO7BwPfN
cXIC2+MJ/7VS8j7t4Tb5cjlWH35LU9OAse/BtrXHJO+CdpOmTOXgAcAcN0b5v9mE
Xm/jlYU1iJcZlBAKwKptlqGcuzfTFDv7uRsVABrBeq033+TrWRKaq5r5xN5fmkxX
MfZNftUmPojPu3TM6fDS0hGBkh9v12uH/sEGp+2TMJQxrd4+y016LrFQds58mXp4
CUWJA0y4EC/F4S2fYzgPRwn2bdUuOvVLrUs7UX3VZzbpdnGAtWUA0DSQrjBGwvkH
lQEAJ4KuQroynzFjQ4bN0J/3E6yMAT8jxDyEF8ThOulob+wDErvcCv02k92WQeCv
Ea7F1k2pfqNmt56bqLgAq/EV+ihVPMaUFHB3qhkEiNN3Yf0AM0gpMETMWHvcPyjZ
1KYupFMvDJVJqgYpIj0ZLvrrPXFyer/+kJY6whtPEsgNmvmh8SAuSUewavWBl84X
6nTJde+/abtEFUWNfK/VUAGXGv9O+hrUZHV6rNMCfcaJUxT/rSHr+bbiFiiwbMIP
34fAkct6/CKIWUd9TlYyWKibi5a+twmC3W6tJxXMUMAUcAbFLO/9/dtiyh+1Vq62
2llyF9YuA6ygGwSGkbSCk+rHp3/m/SEHhbAhC0/r6wkvTokl/ASt2Mkb6YR6gzWd
Vzun9rUpT1qcnizxNy4hlmuytx/nXqYiLhTzTaWS2976n5Tv4CrS2PGxsl03nSml
Kez5xNBKzTxVsJsptF7h5JZ65vQtSuQZ0EHDPvTm4DE4NHIXocN/3Tna7f3aj7hO
cZRuSYcOcbuiYcdlt2agxT+HYbsJMcEfBKSBHvo84dy/PhowKS0081mnFan6O+3R
BCatu0FJXyG2W5hPX/12nxtiFR21Mw9WrEdcQAIb+DBEOSImebnqGBjsSn8cjnEd
LLFFncSlKALUJ8XpnoZXkLktpIiV2T9/Qql8LVt+JPzVJlKmwu8AJOXLpT/W8i9d
b2Sktj2LxxRoTS0Ku+MSvfEGTKBVDcA82Y/xLp55N1WIjL8xbeTs1RbcG/obSVQu
oQdlgNKs1EqvzOhIpyPhJtWQ7onRqwS4zTei9GJ8RTve557/vbne2GeDXZVMIJ0F
cxmvreTeA/mCVg2bt5/L33OVIkdiIMMVsR/Gp0FaUi+XWNXoHwjpUIGQOc7RuTW2
sZlQHZRTjxw1wWe9/xWXOfMZ5TQX9XcnLr0HAS3UaupAwIZD0oyKQdK0n3MfHAhy
Gsz3PvYo0QStYvRPjIdKcTHTSvYNzRxNgBQD9CbzRm/OxD3bWGYFerjQFzcnpTrM
a2BH5twicJB2H1ogDToYZ7Y8V5fb3P0kHPue1iFJLjWpBfDU8/+HVud/n8lJuzQB
cq6BzsEP//UMG9TlIRD3mnsigy5aCxpDFjN+UY3krOC2e7JsDozN0nMYt2F52BQb
edB2fkcUO5larYExRib1sn9Kq3+SP/Rgt9BW4os9W+legncq+FcQPfxNJu4PDoEc
cJQrw0KKyXoHZLgXZ9C4/p92MQI/RhAbRu1/LjeG6ukSpO3pRPe57TKpLhf2jn2c
fRwavQ+kv0ZYh6kRL4Y8/idXWklpE2wvoUuEtidD6WCM4l/sBw8lQrsD3OeEqpCd
29Jj4zQXxALZub5o5r3ediEsS6299gmE3IX8Zyk0MIYLAIgHipDZXtPRkE/bYhhK
BzkwnjrLfMFpZoGcUdOcM1D3LsoEq+QqM+I0elemC40anfJzZpB3KbC0wjmJSu09
oSZBd8L6mKAArnY+g8pnUVnsZGsKG2xXp9OqsevPwCznyY6020icmT8SNegQXjWG
hFZY9JNylRJRVxGtaFqB5qz5QO99Goa0cuVOw8SgiOztIHZyRZCY2fkKDBVwJcHK
Q0vMIl+qKl7V6W65MiTnhrVTUqXl0GwgwsAfyNGBE3RyRo3EF8rK+hYkuU0SwP3L
WnjYDXzIRIPl0XTAdRHeO2nL/wOgPhWqZegIoNkrp5uINdaiBQNyF1BNhtxN7Yzn
hCuqK5SanXY1l4si4xMGMIuFqmyuXHkskK+8GCnNukhC89hFlgv7jiKOMSedlttM
0CYp4dJx6+JvDIfNIWHabpekBjZOH+y+CJccpJ2vI7UckMZaSQTicMN5pLVLLhkH
NZTHlLrEiBR6kEC3NY+jwKkxPpgrAPWNwbM7tV4jJoigVwKVQaZZba6/Nw96ZOky
zwrxNycIqA5S1Bs/KU5IhkEHvuVqdk478HVbJM2neARs01JehKB6cSmWKa9GpYRh
ilmzd/m+6RbBsvBwXZiqmeHuK/DfvkyyodPV2wBtjfNp8GE6gAOJKrZjfvvdxyAR
QEyPScrbq4aaWuwAsxfeFq/KDfhcgsXvkU9QPfYieDWt72nwcXiXGlismskKDoad
6gTnLTxmB6NYpbNNIUAmnOGNAB2X0ugWHC9DkAvSXoXpdpSnFqjmwTwzvYBPuVvp
LgaMpLylWmZXHWW2/U9jJAtPPFrGnl/2X7FJrfJRat89zjou2t7QD6h5CALTOlW1
zE4PNPWJAU4aWznS/pL4XW3l2EV46jCqX3DR3lLNxS1mPWNAs4H8nve/MA0U/UQr
vFJ7xXMboIRYFrjum4zZ/NFiY4916nKz9qyIRGRyke/ryPxv3pmzcaHM3nlqtOqP
KAbE/vjK84N1QYSOVWZdrmFUjLoulr/UitmoOJqu1DMgJm3SAPFfKnXBUWdo+WZk
whTYYhWrOHydq9kaCcRMQbW0yiLssO6uWFi67eswJ7HA6pkfgS9xY186EnAWhcvP
01IJNxs4SDP1tGOLoup2t9ksWJCduNwVQPSXHObFF2csBQWP5XkoEkOOEsBsvWBC
MVKS9P7y0ZWbt+PSPrruMjGfUlS1qeXW3q/iliY3c0Zm91e6TrNAGpWmfGPVCKlf
Ta/CsBKmGdhlaXCRUMapABgPAMb4VmaYoruTX5/hO5/CU9II4blbO9e9Vnlc/+b1
uvKZojk340YH5Y3ZuhDb2Sx5xIbV3BpVf8nHCRQUSkTvrvjF6O80J9xOPZDIloWc
txl3zk7iMdsA3kS39hsCFWaxlJ8t97yreBg8gNooRYZJGt1Vcqp+U0vQ5oVHNU7g
TjcL20ixvJIaFKEcFk+JL0BLLVi/2NHlYr8alY9YAfFsIGNyDGO1C0y/hk+BVdry
JrklJPLY/vd7kMna5YWsSP9Nf+l2HKwS75HidG6i5pB6OvZz2vi1Lb07E0aWdHXc
7bsneySCALBdHjivKcIJEAzUre9wA1oPO8kz8oJTNqEw8ptRFbR9HHHoEt7s8RtS
VKEIOD35MjzRMc9xxewGRJ0Vfaplqv9jnIAxoMMwuDrxO+tNqZZVzcaRy/bAQ53i
a12iJyb0DgRkjBDxu8yg3cIQNs6fHQsxz7a7MDshsDMmAkiHWwF2/4wQJdks32bG
oxqOYfuaBwwuhvpUourOTN3WKfKoyAhLTVo3t6/7rxkiFZtgDs+zrOl2JATZVE6l
l1y8875g2qX8shH4auK/PEJe1dggQyCK05Y0X40t+H6Grln2jkPZyjPsy/q89f4v
UYRcTakX9xrksamwwttQpRMnnjIxVN/zRNnGoAR5RGQNpBP17LkepM3AzRgnZw4C
649z9lWqskZY7cITglJbcaDGi+LHHEvUIIPnOGXYl6EZt3FI8eLwG5RvXTGPcHSw
1rJl3lLgPRhKec/sPcMJSICD0yX/h53p5jufg8ucJAOYqKi2AMLSK0/VrmgcjwLz
cji8D+gYUffWxoZeRBvps0B+1UHtKfFHg05FniPP43cuCdY1DnMVM80WG8Hhrsas
FhzM0kSpn5eRgZYvdUB6xgTvVkUNYD9M/z6lv69t+pWu8igi4BrLPwKHs3u/pkYJ
oROH+uQo91RsP7zTJgoWisAPcCasNApYzS190Cn1HMdQWMDm4Ch8B1lTCF+DtFIi
QwK9PYNVgjYlNXlkaFbEqpDzUyS7HflTBSUqwBRNLPi0ErwBZM5HkpfCOp8wPHb5
tUymLC84+hyMn5Apjc0/BSTz5jM3srwFBSLoyS/dLfijtS3CYx9nbcauL20gOGNK
HlfCAizc+cBiJjPdMjAxqcQKuUGsoya6rqJXq3WSa34ugcWKssV7Jw+4GngLfzEh
siU/rofWy2KYWkeAwZmJYi1aVMqh67YXGDHvwGOKM2lPhI5WY5aLazGu3tKeP1ST
hs0zAMvBNQf8Ryj//VNuRYAa1EIUxCGiro3dekuZNNYJVQfb9B7TKWu9SuFqZmEi
2C/ww4ylZgfVb7+kq6L7IJkXV4Pf9ULx6VYjwL3hCo0Tv55OzgaJSFufiDn+k4vM
xghlpu985QwGjr2tIRgn2W7/IYyFYfHqFshzpQIiPCIfKmJru2x6YmcF3XirIoac
yBGp2xzqJ9CGd7ZiXKD8nFlLSlLTruY3lgwfKWzOW2ms6VzQYznQTBNQvx2VivrK
2gmoUshh0OY516XB4NiJVAOnyxDgvQFxLqkfNr0j/EjSp/tLqW0+d9zd+X1OaszI
gDr/oW4lIDMzuqV+V6QaILLK0GtfRxgEAneyiVyFSr5vBIOmdvLTXgjLiYX//La7
xrV1DIY0MiMmlJ6hVXkg7+PHKWp8eJ6py7R1WwAFVI6IyG9HUwFL6n77MuJsl+9d
d+OEHOrZT3k/TA0roWLPS8UDvTqghvusVSbXAVAPDk7DjS3Ipymx1PjmwJDNaiXp
cHuxf/JpRKTpfNElRiU2z2DCT4eZ2UH8thIP7J2Fde98y0fLv1LtEHtzaiiiFs8O
qIPVBUWHfWKD3blRrALPZ1ZpqtWlSqO047DYutBLlggCais1BVeAhPI1pe1AFywW
svvOgnWGYT5wd9Kq63zG8a2CTa5S4FhLuRPeHsnKqism1VoPlvvzYVpOkehVw8Wl
THCg90mSGmxB4iznIxvPb7t/LYU0oa+RUzHTkMkCicoZVOApuWNBGRw3dVvMTuEx
1x5vvwBtdqF6wJn9dEdhUgmuk6B4b6zh2udfUdV32SSsmquv+jZ3oR4tbzRokTh7
om5DdiD9+e6quuP+fsvK0MUNzl+WkSyllSQIkvxDsJ4rNItz4VqQ43sitm6b8CDe
IQVUBFzfE6IhgThzkNmGfaseKAkMQ3RdJJUH2iLlcZb7iEcxrwjYjGkVhHxI+TB/
4G9sznaVJGvfIcvMEXcWlCG16faMY5+48jm0UZMAVw2dj7rsURgq33xEj+pMxB8C
Aiz11cI6GQquyGcXPrdsbx91mM0bxgG6+W9ziCOPBFC/yr3ObGgt+MsDcfcKAroO
2hsFzz4xdblraUC0tLyVtl2IBfT3YDc0Jsd8bkto46+0jlMAHX/MWmDFqPaDx9Fs
31I9174Xj4tXHqYw/GJgnUm+pe0i6I4rpLeyYWocAAFayJXifph0/C+MJ26o8lVH
5g5pI15VIu4ZRCXUAL9hYeiCw8waqRR94aWGn3YKWgKN1jK4AB8YGs+BguoEWSb5
U+jgfr+of9bKAAVBM9tqxBitD2i9SNAAoXTgDLuqjvWU3nUbwC9UEkitMxI6UGzT
4s+YhM5zQnqz/WMce4COpi78b08ew5kVH+XpEPTEGgm9efl8Iahi8KKnpIMBSz1W
z1Y88LdGzYey6KnZ/i1ec8eCLsN/MAJIo04uuHie2nLtNK4IPvYOAWoXKuJfSmpS
3TUhGGYGC1ke9jWo6Cu+fW7yBegwzz/keZGNlKPCkXdJ6yhKmkPvwp8f7Rbq+Qq4
3rDXywWoYdp0Fk1ETXkgTc8AG+D3NAsp4FCTd2HL9lbpmlb5hTAnWdsDfQ52unuN
yZ454kUaASEy32Ul9qe06B29A5/iIJMxswQhXhSTpl8mlXJssRsN6Vwct/aQD+kP
iEiw/z+bonu/7+ExNSdkreQ/xG0kJkD+FvG4+APdk+wiCVkipUGT3ZS06mCiUEl2
UpNFqTgrV/q9bcpLtl2/5ZmzNtHMQutiHwvUxm02cVA5q2ufq1nL/87JRYq62cEh
pjlDE8CI7Mk3dGGKU9m0Zw31nkO1QUHwLxBJIirFIv5+/1WYeeQkL9HUEI/LXUZF
T2EagpibZgQYBQKBqn0HQGp3FKbsq5rSlfI16t8IuYR+GnjKgD4AgWcP8PsV91oL
elDwHZ2sguvM/FaMcSun1FfB/IB9K+pgxswUGQK/xs5391iRfsT2hhVelarYaByz
0ou11mALv4BSE9ZOSG/afYBzOsUGDVVHrDUIkSnwAupYjojvBwz6uFotXioJOq+A
Qnr5w2qIc5lysPtEdbDlL/0GOwuObvW5AU940DIhA71KqBCeytDE4BXxXs53w7zP
Uw3GMC80WxtaVcbtNEZFuoKkzYQ8KC5MGGLY/hRv2OP3C+DKX6bUETuyKPXp8sl6
0PkHLpdiw/4eBPUcw81u0Wds9AVmQRiaqu4v4ACSe8GLtWApv335FsfrETx0WwMo
tiNSrI2KIJEMZJD5mNx33Jidf1muWTo2wS3IAn3nGS7qCXaogzXRUyPOVU+1uuos
kAAeYNsC0WXqBBwf+NSq0B0ByKpHDtAcYedO6tgtd9auMHyeskwcbPlDlUfiHAZA
Y/mUDylrulid3B0kqLQ5sYBFBi7krC0Mjv5NYSwKUzlFPWiRe7R8iSKBELlskG72
mrrvH8Cj/Zc17aUJsRtg8zJ2g2C/3+X6bU4wosgom4ERluo7QGs42FxeO3muP6Rb
KiVp8z3TER5zKLaMhaVcKWPAkjJg2BL2g1yCVrBb0gr5fNY4l3OaCjICL+NvRcoy
Zb/4Vk5D4vCHDXrLOXE6RTzf5nkTe2XT/+wuCU9nHmtCOkV8LyPgg/mVV2H+nQ3D
zo36FMMZniEcBl7UfaoG/AKPXNmyk6sLcyKrN6NYZ9fIYr8+t4+FvO5v8PVWf0Iv
BHI2QRYZM8p+ikgHTTj92Q/qYpS3/SSXuPhfXzTSOxJKV1p3WNpWDU18lJbGHciY
cUunxQ01f4z8yPx38qrJ8dXzDQo6aMbe4sYk/HdCC8vhvRpNpmmYydGHTATZzV+G
e/PREIxQPHz324Sn98oly99zyEWmd0pZKRlxmSJlJGMT89zfLuyInSNVYFfacnfH
wOSJ06xhcoZYEVk4gaSM4pNV/PJgAo36uU6FROWl6ihDR5RZj65Y8Q13tOxQ0/Jr
0GGRqQ2SsUcsvfFX8ilj15HdyushPY6EKEPjnNAijna5PIxmtlE76bL5dSuC66bC
b/hWuFn3n4NZijKeSo34yNaWZq/tC8HViqQWaD8CYjVrcxLZB5NQpZ2we5tH+fzK
YVS8B6/bWbeNAyV5ZvXCLmxGvajFoIrQJvc7RY5NwQlKVIon4a5CoSvdV/OgtGem
grmiVAuczUZOrLVPRxBxJvpYsRfiNgSVK50oZhlOnylt60fqDhEpCxGT1uwveq0l
k1eBGSS6RZbWnzQEiSodSvWrayv80py9GGczOTWiPCXJ1Ew/FwBJBz0xkjPrFca5
sgQ0Yja4uBwLvWQsyYJG6fFqLyClP3gFvQcD1D8a/QR54641XVfdgGltp5Lg+823
WWLR/j6ZrMVex2hl7XGKbFqujdZryWHTXI8ioSs5Q2pvSceiCZCvfavgF+LwhTMO
XotzQr/z3Q8puQyfEY1RHaJamcCl1zHw8jeCRapGdTnYVHwh/UgtIrCPDwA1rJIO
T3q3KRde9pLMcUM44Pa/SHdL4fAUqvPWXd3g5Pf7KbkI99L/V6SAL8vRo5fOyEfW
trDBC2FdJf4DMOkGBcLj7u7j3mEwfpeyF9Lm0avb2VxQCkR0QoSRsRz1Ybl5skdl
arFj4XEyxNfQaRTSSvgdpY1K/8SB+EsemOgl0FYwrRUrxc7KK1xtw6PCeHAokb9l
t08LgB3inFnjwJREcaz+VVsQfBI00XigvF/ijGcW8ApnNf1gKN4ZZOiO7Q1Cas7m
0qLYHBaTFkpYq4o7vTSkZ9awjwuTtI0A6HMwe/xV5wqp1g4GX82JUSNdlw8l0Zib
bgnIDmePZweTtsEOI9p3FXygjUcv8TiIrWQfr9Vfaj9RyGGLB4Mc4DR5jIABFqhH
Q61JiTLq3n2eAaDug4CTEghMjW8W7tt16qo3bwqHM6jtyM1rrb9A9uY3j/Tz2cei
4H7v/d95dpPledVD+imeGyGqGZexOTI2zywBGmkqLPxUfTLE05frMkdiiaNFhqhK
uCcBOg6El5/8opgjsa1cFCBT+nOdn9O/UztRjt/hT8k8SxbVOS9LTV4LBpVL54mR
TaiGmMxJYcLyyxcaGdreDku/SqfvXFQZJwgcK8kNBX8Y+MssyYO7h2KzwvoZq1HH
Zt3Oxauw9kjGc6uoS3QVVwH8yLnjYJYCYJq1jxGBoPEHoxMxXXTpvEzUfoQEIPHS
9vFFVVYi8IV35w2rKBcRGTvlHwTk/CHBwDZLPrZZHDZtd66e9jDnrSX5gzEecNIn
Z0ethTvDCOnNnvJm1LZVAIOw2sJ+4yYbDPe0W2u10knw+rIOQbNj6EPY+50jiw87
sncmlvaBiU8OFrWC/T3S30h74kda7XRylm8fPG7C8DZnSCzREMIJuESorgaMpTbp
dH0R9ktZmzrLpLp9GcNoTWBkMjVU0d1udUfVm5+2koLfDiQ392ihfdiorb9DRD6V
Y02SCTm2s3yanSmwHfOpnwnH6Qp8h8U1r+VJfL02bYih8+kRZUBppZbq+dMskPNz
uqLhnV0/U+v5gxReSkmj/t3diGQIFtp9Qm04pM75G4K3LmgcWQJOjZEvT6r+Rm15
RIJ5Uvcmznd4ETiKsBfJ3TJV/JW9IhhqJkMm3hBM9hok1/MhsfxkaBPjgreYSBra
7buwMi65rlqPb2p2fPlBfwese8KiBZTkCdzGNNGX9W4QPy9XdzZNeVd8O8C0nsc2
VOU7bGEUDFmZcF/BFsGEetvngSYtmwNQHlMY9dsMpz32qz1u5VraXgA3kEhyfIge
7515j8JsHtjMm6ySlMTF2qzwJQhAd5zf3Dvc3C6/0PRv/6HCVpDkHwoe7+Qarbnj
5h1uB7Mir5jGrQ/GFNanX21oAk/cIfw53DRY05t+VnsSLG6T5JeI4MiJdjnKeCV8
98zjMXomc8a4sZXKkT+s6R5QgKLESsHDlDyPYvKkmV3ZSu3ggy7hwUV6Q3zIj+Eb
JDmLg+DUD17siLcrLzOyWHANOhueQbhfJMY5AtJXCGFC5t4cu+AjM2oKf8+LD5mu
ezsK1XUT7Tb91dF72CCU+4YahtY99/xBJ/mBZrixnMQxLP8z4HsoFUbW2ytAT+OI
bjV4zggEgFp52EQcVdwRN4fn6e/2XszBQZrwzy+ShUkqDdA+REwaLRbtTPffJ8Av
yUswPBVqbEKHbrjpi7eL4MLkO8li4EQpIPD0qKTT+ITMOFmwJYKSM4R2yTD8Nf6E
tE0KUVXIqwlvofTwtVbzxMDIq9ylyuCdelRuyr/OAdj9vRuDHMraoNTL7YzgzuiZ
xxOhbXgJ1/Gwn3rRwSYMmzsttbhpIto5LGoyE3XeQnCrmBXZiHW+iTlWEcAWLppv
f/YxURMYbQO3wHRzeUfLKBhoAjsqubkgyLgsLVE8P3VgEjAhkr1aHftm/jte6PEc
JVolLsjs7RfGi4BwG1PWgQjQXOE9ZDmLGhAQ1w7jq/egcafmN7mwxf80ph8J7Nke
3HBH1zwgYHfRpzKct9UmsAc5MZh6DCRiH7GZMSVK14EriwtyQeuyutyHZhuL5BqV
O9A3ptUWXFP4iX0k0BDd2+MVCyj7+FrY5dToc/+jO+F1FLUqgLRLkTbiaojRALym
rMTsjfS25kTvmjL4cxh0alG5SO4VlZI2Yx5YzMzHkYT7p3rOMOEUDFqQE52UG3+U
vKhyuIUlfoQu4VWiKQMhptFY1FYMWLDEmPRsmNilbtomLTAB2h5frwYdsRxTfiF3
WpD6FFxfuzYa8xS7sozuyoeSvv10PeJc6GXAeKJg09gk+qMFO7yDqj9H9ckPkP6B
fsNTf5gp6FOkr9UuoEYS6ZP7TLqDNAZItgf+QEAIvUcAfxzZrj98ytUGD3l6qfWc
FPAfM6YbQrAeaN+4PUI5U5k5dHaX0cWU2DWkVX6B07oR8oIe8kHlr7j4z26SoJ0h
1kw46PRdCfxmQuIAviU/ftIJPKHXqHgSJRzjYDgMPHf3d6Y0BDDllZwTFwJoJnYX
qutQt+h9NJZGOC9+xo7xiC+sriB4gtol0sz56wD/pkt8nk423er/+1sVgXL1imbk
86ypqKNTSvpE6yPjSyCSFLoeIoAkT/Z/oDs67etR5N1/ar6mTSRmvf++9guNvYpw
WFTyHZkvJe8g2u3DsGrHPnAImDXXV861cJd1Zw6rFBIF8BmYbDvM2gbbqyW6wr8l
I/0xqL4DDLWGiStsv63d9XUi2/LURunNEwRas3be8qeR5HlnyVLjHy7nwfd91408
XLjUPVsDb2o1m69T1GbN8J2fvIJU38Ecq54vU7dGn86AHx7nvob7aMVp31FODnr2
rJdpIHKtBLLMTv8jrJQ2dqeyryLijxvyEUyucXu+wGZllNQMThL3WkzdgceD6HW3
EFSsVocVmDbG/ks3s8os3QPij44gfvcGCPllyYFuTHJJ3CVGikmXuzHqdG7h83Mi
p8c2AzKRAOmyeRIyhC5uyzVpTjqf7wWxZW7txc7YlDz04jyUpi5ZjJ1E3ILQyq2p
5UrkkFzsYB4sHvk6eCVC3aaBgXZBlQEeT4TLhoJG2KucxDQq9wWKIOQve1xkJ69C
ZLOt9XznwWan8jzUv2669UVOLrRrL5NWOU1IDN2XHRSk4FTCQEeAkE4ueknGo39u
Avbs/qdLb817D8O6x8U4vbFnU9wa8BWrkkaRF7Ctl68S+Q2qJ6I88RlQ29TFT2s2
RLeYain778pBh57PuzMuHB/DiE3htNqv++E9TZLQf+Y5mCQt1yuoPEt9AKJsdvzg
Dfx2rPHEyeHWem3FUh3JH+7JVuGv7+yT5vEo08LI9MDz7krRDw5gsedqdS6vLoMI
zPkd6Z/z2TxJe4ar9SAdy1xnIkkkGf2iBNyvp9NSLqQTVDel6XjABGSCVO7I6vff
lLMVnUKc4vdpExKO93+jCG0rNmeffRbq/WUrzeShsDaWQ33y1UV14f2E7qFnIEhT
ZjWisNl7xEOPq17LzJI1aFgn6HUYWjQfK4Vkn/6GObRhJNy3Kiv0ceSsG+FbayqJ
MmFp6ac1rZRZeiuZks/usr6Wb3UWOyKdGTM8Jad77Do7T7oeuMM6GAx1B5jDnwIu
/TWIeujbyX/d7PGEDIVvA+YtxYLtbSBCLwky2t6FP2HvfZZkLhdFl4SldqL0g7my
Kc/4qYzuKQWs7W2lHIi2TGSqpJwB9oR1jKoM/fYHXAPlT7w7+koe4fPw5mcgQQVg
uy1ny0yjBS/MC+F1coGfB3f9/w4vKJdq7vQWZ3KJCboM4CpIgBegU9pQTv2u335R
IwIxkA6W8b5ZguByf3Vj80M9CgZm9nkAYeThZR42vmt5N2UapNqWzLkvS/6zGNbV
CQVKhN12+THuKajuiyXZ2ay/Bd915Uoyps0WgAcKc0hCJjx4DgNKPLpYSdMbpuhV
fQldmrNKI79loxppRKW7/ZGWRjYL5PcV//TE11cpEd4JKrJpSaNimOSW2Mr/LYb+
kQTK9ygtaJ2dCDs0s8FA5Aaft6ywGQJ5mA8PWF5xWv2Qlv/Lgsk2bkmJPOoBXSdU
SzsF7hdsn703/YuHM7jT6HQJKz9rAhUEdnD4zyz89W3H/H3m17jpebz6GMh/mVOo
C6sJw+dgBt+lNTVvokJuO39TbzftyeeQxDaJNh14U51WxZcEqMBgaqmOuZN/l6f1
qUEwMgJEj0piOff3NCnmhz8MDtxUJ3yNs44Zbj+e1qa4Guphx1jdeX11XpMd0me7
x9VmkHZwKO9bFa/xUVyz91aamywSOx8IN1Q5himQlBoG2t+AgIpGelWzmJ/W9wuo
hHjiM4vUX3mexwr68h5y2wjfMCifvd6nef8g8ERMbk6eQuBcZ1P6kc/XOAFfxF8N
WrDgc/CGOxoHfBZe/ZPAmZglaMz8kJNVx7MfkRchHsi78fFRJW6unvtILdQ4fNYW
lnVwnc8fpFt7eMQuUt+xE3hN9/LJz8ZuZfRcbmvVpwWkgAAaGCWZ7NYF2YDDIhgj
hIo9q7k6Y55kLP/gmXxQwHpvnDEV2T+YCytYIA4TQYS+DoRtxZfN8jx0jAJfzzzd
8D0iL3R9NAm348pQ7XwYcGBuni0zPtD62yZY6X7yhii01FvCRfvUqzIWQlqjHkb2
LLtTXAtQZ1XhYx8iNqmdWNSV89c46ow1D3nTmrUmD+undumrc13pZ2aShZVPVVh4
Jc4dL1d/IhA4GKXYy+vV/qYPwZC6Us8yW1Wyk3OOqwsRuZQ9D9taQjRMp9kRUEXl
txOyi2Qfq2HjvbrRzOw2FTOXeYIuBcQbHSiC72FV28nTE/UooA0HCjDVb7VNI+6f
S+eEAlCi7Xhah+VzQme1IlIt3JFhI2Q0uWPFyb7C8DNfwCGWtgjHoMge7CO4SgKn
1tTXWuliQ6Ib2HAB/LpVRc1a/fyai0oyaU3b+5Iey7Ak0DhmK+OgOnp/mpVghcob
WhTKYhEKDvur4SljwdrjxoYgTXcqjic+FR95KSODWdjD0A6JYBruBmI/rMzkfX9K
rjwVq/G5C2QiqsJt3Nx3jIJO8IeEarn8uzuCGsR0QpQ1ZHbyh3y+30Dk+XHFcbx1
DBCBwxomIKlEKeZPuheld2+Yn6k9TR5RTxPdwSVmqu8GgP2rObqTNSFNteUyr4tg
HZgvGKYgtJuGQv6WBzxLhBCsOnPnGttHEh4g1gw6BLSOxR74Mpz/mhQPWdtwencT
1zeiNam9UUnqtK+EddN3/9GOeGhD/Osdef2hZNmcXzeHJC5FRZC7Ez6SZb5oO23W
mONy85jT7Phl0atpYBlheV6zdrd4nRQj6aB4w8rQXdpxivIBpK0R2dDeEO/k031N
K5PtkNwWa3ZXkQ1l0x89DKWKeOxKoRmEaOfc/C+qiq28mYkHULaijGof9ZIk1KpN
wGOwn8/B8Bz+8ry9K9LOv73RT+ewGNzxDcArUIbA9g971tEPpzL52hlZHAXTKlmO
89LF0ByrYPAkKEj6kWYQzXxqc1KQDHfrg9tm4T1VMp5dMPRKkWO/BXrit/2ysKju
2AROfd03qoCfRW1SHaewZxrcCv2x4Xut44H5sAvipdooXQRcZIvymG58Xi08w80/
44yjZq2sTRCnWTgQEU+KQrM05k2MdfigG98DfGjBkR98ubRHS0A61UsezoBGMi3U
yG88ZjapT0XePheAQUMPaUdorAQlg2aPJRgcsURvOyGp3Tx7cq13pA88BEDbP3dL
Y6Z8cIFcCyiHvyDvrTBSTl+5oA3n7RAlZvqBiTgN66ctdSahm5cUEfWS6GpXYxWX
AmIMbtHrL5MVMP12kaWz0e5oJ6IL2hw+EV8oIipjxJ6r74ocvC6enbQtdaO7dkRf
atgea6iP2BIDqdnelMprZBN/A4OaBGcyEZJr407pfESvXtI6kM+7FkTgelxHDiz1
S3LMZxFRcGRoiMb8bDC+YlsHAwDPDyn05M8s9a6sU3/FSKzcHheZ4n2qFFIRAVX6
xlr0gSiyurwl8DkZbA/tELMylWaz7mUm6XEoaGJcCL7TPKkOd/vfDqld5v7B464F
4rGy3DOXrppOYgh14uy1PUKD00BwKum3iBNethd/Ibi5rOURmLJxNPRTpukswnGB
6qfzTk891s1FkApgCSupCBLbmLOk5NhjpDxYCSWLhn92HhLkgIoMXM/J15YnjNAA
BAMtA76pAi5lKPx5GZzCexnYhru5sCn76irVzUmCPhqVVzrwxLy2RG6LuCxJB4TR
3Sc6g8LGtaOmuzEDAP/ox683o+IGtIoSrPelY4s4RMXLdAzKTjYEfxzEQRIiYxaI
qUxVS0cIDRHUpx8RsHljvKZwkSaB+HXJ4535Um7m5QgOmQAiJaR/s14yv6puoZVv
Vxt7RkMGt6839d1VBXPbyaoGNcDXNWbkbdmBa/I1jxjoBVNYAc6STB1qlYoNPC3Z
+2KBeVz8uflatWX27nwAnbz4T/dDuuUFNbjZ8W1PYE5bXY7Q7oqtQ4Lldcl+lwmh
EK7uw8a9c9Gzncd2lMP5lBTIBEDi/n8D3TPLds7r86NHkrhYZKddx+KQpEypD3v6
JbVJNIlJS4iYvB0Vg1SXiI49+ii6T12jtcvm/rGDQMqkKEwjz/zFsQHfrRO/agoE
1iSFNZHt1oEAMkUL5qG1JekVFK1cYtxtQbrt29OvB1ChzX1FkJaSzfgnXTyPAd2l
o8g1EvdzbaM74JbYmV9lyAN/R12oPsNC6I1xH5wr7Xue2DViwTpg/h8A43eBLk6r
Q9U9GMdh7/7f+1FDdPcmNNxGddHRx/Vgrhh4Mgz1jRPyCzMXBdY5k8OBHpIUgkdu
sOs4PqPA5xtWV6UeHYWk53mYFm9gaT/S41R1UE6vP8bR7kkOdI7bYOnSPXxEbNBx
M0K0UvVphkyPuwU10RATz4IVAB/IplLHDVcdwpXxEySCY//giLQpsZfFWnFEgnOa
+z0yAO6eMbt/Fe97yhHQ7UfIh4ylEatqlERSoeg+DXSQ4DFUrsjROsCZHy8h7NcD
dKkbyFNpawPJRneshUJC51MQEpK4mtFtpU6EovKn6oNyixQm5OZdYbwyBCa89PbH
d1rdLFnUWQ5PHdtYmaD3Xu/jriVHFe5eYzOPieMmkPqKEzGkmL9milVWT2XXFTm8
O+cfd7PmC76HTId8y7MgucOZfjvaeeiRLw2GUI3zub77ra41SnGvWg1c44+8/m6r
+cLCB5zjiIdbtYXT2xRezTxDP5ZABsn1xHP3YHfiUBrjT1w0d5J/3UQu8NHwaNrV
YDrLo+49hEIrC6nQ6FaJHLoEfRVUnpSOgJy0p3vBCJypBgoiUoJC4OiLXCv2XDjo
x+GhLH0LAoG2eRGtQ39YvN7xbYFmKqUyHUX87hnduSnhnK7A2cSaCevUe2Ux9L+X
wkYqusAKTIbZl5ANrTakSHUyqLZrIHOu55zNUxgkXHuVOFxetxgL7/9VSFG8zVOY
lvz2XTursUlzhxSZnpmjk9nvej1XQtd2aAljXWk1JbkfTfGTsWVQONuCWdARhZWA
DGA9r51kAwJSQegKreZQ+D426v+ZdcDjW+vcDSDhyp2U5lJUk8/w8SmeHHaJ7kmb
qyKPW1ny9oe0ECD1mRjEhC2nR0VVO1cOwXICa439n/PbL5JzVBQTPcpy/2EN4iKH
Xn39oE/YgeOvsBl1Adrb6hHWIse80S3xbzXpJv3LYYe6gJpqnlqM0bI/bZwVORwz
by4eRMbQTaZ71reUqJXrK6uH9g+CryPv+isCDs5JJkEfozBKz02mq2Zwg3QfognM
ZUzuY5FjfSRZm0hdjWFP4CS3BFOBlnyRkBM9uIbdHTshWikUcjpL0TzQq8hrFCDn
qIcLGzVFLezSRFnBN4m0G8iuUSdmZBpEe95AyyrZUarQuHYqNDs4zhJ/RxSWEcZu
cxDHsb2V/FPrmtQ1IDAG/u+boJh1Vwu/1Dv5PMrGETQLOX64vNiMXdEOme6I0cbS
JuOZZBkVEOmru5NKgvHg9uzgxC2oEAPE7dq2OC2eVxI/lH5ks7xic5+jWPowOpCC
p0PHegJAz2sV2xz56l5jY37JwN0T/jSO/GaYsnPVcxOpJZvXKEpkfuvsUBnciaFT
g40cP/0GIEQU87NT0ylelgoBcTP6LC8m41PG49M5TXjjzKOklPN7a0KDQOz20158
Wg2HjupRljHNPtb+eRQhuIbQrHe9SdrLtaez18KPxhDMM3cPeZCU0lZI9vvkzlpy
VFe/AJ+bMImFz5AvuGwYrv+7gk8kZMh6odgfAjnmiOmLa976PnvIoTjPTxe4uKhm
o4h5Iwp24wynQhtiwNg60gr8hc6+1xbhqB5HX0w+IASLlTVwNCWh5fxTEfK3vNY0
vvaufvkrH2Nd1ktTTG2seJ95l01AvEleAEprgTBdVL6SsTe00aGE4ADnKn8zBePP
mcdzaHcbfVmuNmWIWb/W7cXI16mz4q9C0m60GrDYfNwSJHaxEKC2gv5qqiEfXvEZ
9XeXChHaGdx2lR8ouNBcw6HSlsoGV6GB05W68lyaS1b7Zw271SVTUYfILhj/ILXE
PJnAE3UK93oUu/o8kXcxHlG7utvicDSuYLKaiEZY/yCHpj+nmL1NPbVZHgSE1JGd
2aFALjMMrK1DaUBMbu/yrVbBmrMBjhM3ZCBn/OFz/uYjdj8ZC9lRLC5qa7RY2mH3
T1j5nwg8Cv+meZ9lwFHz1DgtYL2tGcJPgy181E1fzanZmuM8FYAa6cQ0SnEpuutk
jE2B9tzrEJY6GLCJV++QIJ58S4MGUZTeXjvlw/8q8+EtOzQyCLHSql8DDMx8e4+F
ZeEGWU3tW5xjyEOofsRY+AoYkzUM3+xUvmzMJBRjqfCzh+XOogdU5FSbiIh+9gg+
c7XorL3Nxrdh3Vk581uoH2HTiHPkSnKdZFHwEQlf91TZJ/uP6KsmZg6bVS6CIb1k
x0f+nFj4rSqqDXXNn6tpkL483TUB/wilqAajjRRzaFg0+nMQo7x9qv3BDFrCzvkD
aDjCPNMwm1wSAnuSXMicbBSU/WIsOmEsUUfuk267GPCjWadxTSfdZG3XbESQgIvs
steNqZwQHSi7Kd3Yf/WteYx8ZYXMRJguTigGWvdgp+eGHzwAg+WsZBzE7abOzymp
85Y3FQtio1MlFUkyr39cwqbkkf0AJNzF4E5bZgGaDLlFCGw82jId9i6Nc3jrRFel
geKnIENN9XZbLr48tGOJh8X3i1T0nLZABn6hhMRVfOeXAEkIbeuQNYfuJvwv9Ku0
hbHyiqF10+efOfom4Y1QhHGgKT2cWt+MTUBiH931ODF3JsD6NXwftxJ+cg2ySUzk
FwPk2iA7z3T1dd8I/rinjrtiq7RUxg9T0GKMGKryqzNQJBaSB3pSMprrXqFuMOzo
bu0eImsE7HOLsZsgicBBJJeFV5+C6cYwlEVPTeYLIQHoGoUqSEn6CFG/yr7YbAoQ
PxNAcw8OCzH27oCfGYe6TQflAUOA0Te+vvdntCWanmff0qPMpvEqUNkp0cQaFlyd
K7Xs5GWvofpJW3lpCYamLeBvi8sTBR+4SeEUefF8+jmHhovSFdtZ6UxQNK5Eat52
CgqQFKXl5GmDB2KCQoNAr9IeeDOG86jiOUc2sHet9EQhRhxsZ+d3Pj0WeR+F2RpH
49TbG3E8cengqXTePsVC/l30N1iNa6Bk+Xy2bQGIH5UtxOut0ZnZ0IFqRwEyhT7k
crZlEWGwamum05kPMylDH/bkDecyBlMUfVEPcbFlO10KRaf1fdIFM3bypjBFkosh
UaY0qrHQLkVGT1MPl9CbdXg8argmr+Zg7FfOCBWIvYbe64b4hpKoeafsvLGYnN//
9BUdeyR089Cj7RxbaynjN8KQe9BtnSyNyO+QYV2faxBMzUv+Y/VNdY8S36E5pwh4
B/5GIn27GeYPwhoZcTbNQDwY0JerUcSGFPs3pwiNMNBQjhNMwKSxJqfpUm27Rf86
dAUY4M13u5kADK05pZqHVqoLstrMRzb5KWQzQyfRtsCwd7ednVokJcf4VfLK3BFB
rABqG230NbCX7Y8EPWnUmi+276s5mG+erqNg+LIuW6/xUjwZd9GK/CxZrQkCoMWP
AAQuJq3C7E0c9K6p+GvAHCzA8sY0ncNSr35guZz0WvIVKMsGsF4RwlwJHbczEByx
PJ8WPr4Mb1uKuzR3yrN0GFXjTw4bTYU7Hje13RjuI5Pdeu1ux8yhyGyWDBSixic/
lHjRxm9h3dMO4A8jQfSDcziGrlw/1nYC5qLMplBNQJ07FiCrA3SBPiGC4wUyE/tN
Rm7iyGMFxyEio0w2iPvqPC+JRbH33sogMS5UrAKqNQ7o895Tx12IEYWimtdn8urO
WT/9rE0JzZBSB9yWUpnYYrCleGUl804HLtrPgn4x3W7ONSR9woqUIzDWAjZnfICd
veDPI7Zd1jABvY4zMxxANgljQ7ZLzgDJH5OGxb/hE51hTG/WXDqVhKzedR1mKMzt
UhLYILJ5WaH/q0qyIiO4s2imQl7RMEMYacnMD+mvfq5jUeKjgE3+ZwdbJX6Zd0tv
EiJ1J0zBykecSvIIc6zK51hd/SMkZ42AxwMIqCriCdrp9+52dNvJKEPNTkR5Lss3
k+8LMaoaBbedQFYZeciCF9HlXyrSidgBNE5xbbG6Z0IHutNSNX0VhtbqAun21UJO
FzrOYTZLgyVgg6EkSawpRTlXs30t+7swEcrhdUxzDHeBxC/IiZ3gehu4ATq0vcL8
Bs16Q8eWZIuxY7waKR4u7JLQDqvflQZtdXSp66nXTvE1f9oCK2l53e1gpyUJrpvu
JFz4c8wiF6jUkkBnIuUadYiJyyfDW6OzEvMqkqON3LGDYtr2SPMFRAJB51+pRRFH
bGEBwPXpXoGLrBnxi4ObjlbaHIKrSAbHFposLOk4IG49e8Zbqrvx8V1d3n/M3ZjR
z8JkWwHtcp/T8lqL8qo7O4E4APaw8ibJi2Pm5u0X9Os6hfynQiJN5ZJ7WR+7Jz4S
BUOqtxEmF+dx1xc2QkrlNQH4NSe6J8pjMgXipRv2oOS3XgW5Vlhu5GkR49epWk83
ePYUp9kLTbC39YlcH+saCTjPF3ZvX4yJC1xf/wOW/XG+oQUXWtEjtEhkxce+8/Ui
5B/ei20a43PObsA045XST/dhM0n1rbr8SPYyT3SZoUJjLClCFIzIpxqXlxGJcFcS
odIXnLvWaoe0dyLYh681pIFrBz0pzScn6/otAxzcTB/niAlQy8eG7TQiN7UCeEZv
fAn4wYYVi8sASUVX9pCXPol334Tsn8vxwIYcM/70r1KZ1npOe0QSAhohB9IcyH3h
4eACffODlOvpFGvZJTNwvSpAp7jP4gWIbF+uup/wORML+hBbEj8dG7Q3X/+43TBk
Es3dEuN6N2omWK0PLHFtAsQi/ywyZTuzsNhCNElmGdKxL06fvk9CdDfGvXZD3q3b
M8XJXU1XdQBMzL2aeIxMplnWcg5Rsm//DyJWDpohlgtX7+SR4RTlKYi1sKh4wkDN
cR/85xVVIeiPUhqj55nmoDwYt4N8J4+X/896t1mnx9rH4fYRokVHE5mGX80W8MCX
YDu5NZrAh8I5yqO+S48zOsfwDEwsgb825sMsa7N4oClifeIMnW3u3P4j7kpKvAcr
8pjaTdWQdvpB6aFT8fuQWJOo3Ud0oSSX6IzGVciig06EcgvGoTV4XWYbivtN0qeL
5pDP+t5mm3Bke0LgEyfGyeNrIn/AIr89CFdDTqVDhWcDby5kKWABzUWh8MS86Brw
2B/TSp3QUeM/4ET7Xq7g+xLZI50EzsvGsTYA646nFw9mKjxPmMZEXHASh7CDZAzT
jeQ77ExwYTj6n6UnuvqdBZIt+Lau2u6/iBhXCueC4QTNgAunOHJJNfcxyma29gY0
1SjWVkb/moehAgbSSEia6ui+kuZIFceG7vHlMVcJO6J1xksOoIcz0bkyTdudrBCo
raAKfUkE5jTtYvJxMFmyGmgQNCkJPYDaNh7hkcMlcXFhPUvl4+hhQOKOi5igL0wc
dA0wW3mhg7m3zWPMCcN/LL94dvkUILxJow6e1s2adVTPpjlb37rzyp/q1KXaZIyh
R5QfrrrYCe4vEHGfMpT60S8i+ml6mbSTi7xRDfpjMer/7pAybP6Wrlcs1H1cvDIs
gulQf6qa8y1Z0p3Z4HV7DSc0j1eZMYy7y1UMMuz8P4G2UBYOu8cBkvn7KOSmuLrL
bjHsu60LnlI1B4x7fxV6QV5eX3AeDu7oJjAtC4yUUAFT7/ES5OJ7YZCERoV5aGA/
Opyz14GpLBGUbkVvN5aJUyg4Yf4zKf2/8+z4Ak86S9lUFme/j1XVE4ab3W6Kydut
ZMJg4mBZycImTuukDxphvK5/K1p4+fCcJJlx2W1+qXbNGDfRxY+6SLt3/M1D7JPP
q7VK2dQZr4qpbY85UE2Y5qynxsm2zR2Ru0kRL2SK8Ocfw7Wk7+OITi7HS+CL3FZ2
JZzG0TKqoed48jGgqWTeZfx2Qz48bqV2xIch/OkX98F0rkzSZy6z369DZwfZ3xnc
5ErEitcJvLSrlrq6YtBuJca/+w7gkhk+KN1ukUXoXOH6AW9CCJBlUXA/r5tBydFh
W/CdRb7e+Mi5d5bK+DLAGdM6241gsZ/vXKmM+3MzG92mwlWnGvf/2ubJzJtVATS9
EpZmbPxULpC1XetnqcbkLxaHE3LI0h0+/pdkuRikci79uLQNpsPrJaH4qYvhMp8V
0fxqA4lSmitTtmqoj/bx9O7OSc53osiqSwOtFOERHPXxNoEm6C+eR0JJDgwnCmk5
dZv++L0RT9Vn9cVYoaXmPGQgVrLffyaDF9tGBmqwwVoGeAIe5jLGsOhKlN1781E8
PLNuwiRBRMq8r99lggPBSgZRdCC2/CkGl1+utYRZpXixV8wjNyXox/Xh0ly/Jztj
bdbEgW6FwTE9ilVJ8tPsXJpYEkI34thISia6kVYa34YpeKGoiDFnlK1LTP5cCXXj
pG/loXl8fAYdeNnubbMHazJgFrK6lmE+cDYYCU+D60lQUEnds2PJNSKm8/e15Fec
RqjvfG8191+NqOSfJ+pI5NISJUSfBO0qYCc/H0EbBgs8KXZiM3vEKVzoZ+OiYkru
XgHd4CXo0efKPJooP2YTwG3qx65uxcYxMvWcuh5I8cmtAAlkoq6PppUj+kANFQZ8
oaU3cFk1jTOo1h9DgipJhfl07/wMiFXjbJFDcxmN2zCISETUXjEKrfpH95EbGL8J
3Pv/yqdBF7wfOhlSPCpCv+6Nki5HSypTslcHMTPHBT2RymKdGFOMKUiKZuOd58tu
wnJSOGwXXasMNBddwK4KJREd5kxWlqW0qcugmnAN2PYoPWi15hSbDltLN82klu3n
0bb6siwBCRy6ZpofPMbCwUXNdT87htAOrq71i8k5ea0fE30ewxKIkV7qDWi6Eeak
dUEXojVXeOcIUpbrMBu25RQORpxftqh1a7A7mVC8RZxlBazwizkbavN5CS/vUkCO
QCWPhHWjhyekC0rzv199JPdVp4SgIZc/RQnG7W8LPlZJEWyB4WNO1jEOceVPZ+Bl
liESCAH5qMEw30xpW5WKAw78bzfFQZe77OkP2TprzyVF+Yl/j+xahtyS78Bw3bXA
41dhTbIxGNMGQY3CscMLIMhqPjq+MGYaNCpe3DOL4fsTQ/kO1FeSUTLTqQinq6AB
Slv+7P1TcDpUPDNkvhtUivHUpcLdZWHNto95IFJya+bgqWKfWJfC8Ok4DB7Tn42M
jxbgEJWSCcnq9Oc6N8y3tj9IBYVdg6wKJX1zoB9s5Powa3m4QQvmN4JgszrqfulL
jT0WXA5o6DxFFcKFp9TecbCbL63PGvM09mRwDdi/oQI89S1NFE/P8nWnEoGp1YIC
A7bUQvZeZXOsP901BBkQczWEXAMgKH/riHQy4p7wvgqDW2LJv9cUYyNhvudhuzOb
hhVXQ9QXAPsrGMd6kDE9OFzNE6VSYnZ6qyEV0Rmp9n0N+Ny+74ctBhOBej8vm0l3
s9hSRYpulFXrI7ObpkXTJd7Ag+I28H7SemMLuTlOw/Ba4ARghEJbBNgOzPZ84jPT
AOdI9dVM0w1wanOs7ywmDg1F9jr1fDdVluM6aidT//+CJQB/CHI0ypnTtLK6mD68
cet4hr/nd4NrnspX386ffUhOnSnGt4oRjHcNQy8ScKpl0eyWtacbgjBa4txneZq+
/OEkiR5n5Soz5+Dp+Mwx2ewiEoAPfrmriBqJ2lzOuRuX4EEB/sYLiV/TVY3UcH3Z
FKZPtx2iGAly989UU5YvVQ4hU1ZAiBo0TV6lCEjWDoHb8fqMHeNnjRdrc+wCE0uM
v3lMHj7UtLYn5sKVrJEbujE5//HT9HeEun2c7org7sEL3VrnaHI90P+m7diwCCwL
4sMa84lDm30CLoaJkKUdnNDUHnFHivYumD/Ot2EBnrg7FIum94AgE3c3jg4eY+CC
kLzhARUP3BGonVQhbb326qVNdvtF65t2LMTip71bclJGiRBwIAWrz6zEx2zLfgt1
2IdhswEu9UMh3lvNRMrGyCZEDf9YxU0cU67zQIyXomF/HuniBvCS5Mtlk9+bC+Qy
GFihcnZkl+kMfbSfz/4Psg4BVYqqovhBjLaAAGQ7PO6ZNQNJZ/K5MEYlpDni3IAy
+5tGVhHCecKFGxR40lY5sdNwsrupaaY3SWUe0JnDuvKsFXNm9mvegfIg5IL2syg3
b9U0BHHKla85HNDVWhSMkub3De9dObFGVhg6kXOuH6oID62TBQ+gYinLfqbYtCcW
66BQGiMAJGdgkkJPDPEHBhJWPpqIYghUi+SkrUPUCHTSfd8QhCi1PnIXUGoAEzDo
W9fHkoP/HSAFF4ZtxslP30Y0OVPmCYDEnWK4rogp/Z8uYbxvmbzPGkrxEfEn3OzK
vKdhM1mTLVMhiATfyKFJdfKyIPYAYsqXTg//rIIuE69fD7OZ/nNS/qXrM/C46Mxc
kYkjUx/6Vc4oVGpuM4DXbNSmzKl9toiZEF9+eKFtXnTaR5kjf8+ivT3raW7yBaYg
k/JKUpclAn8m5mhBk760csNATi6Hu3V6n5qOEZN9VG8Dy7rZiC7Dhuivay98OTo1
YwWZ5pXSiQ4aeBSw1lRthg6fNAsuJ3/MFWMJcNpCqoezDy5HHQO/Xan+rL7Iq1Q/
6f1J6iJiCoCYj6XSoLKzFpMqjzzL7arEQrQO6KMys115eoiLMdaUBVCASLfnrCh/
UBa9XaG3fEiOfjRn8nPYrk3T2SEIhrRfDw4U5KFlLx4TpW+O0H3zsC/zUodj/4Ib
0XvaeShjIlq181gu+GKo34ytZZdFDHGHLZI447gvebWdvHi3hmPNwW3+3sdb7d9N
y9ywGWhusDP05r0Q+EAanTqZOywwtCprJA+Sjsp0UCBXCdixJmLgcupf7+8B4O62
4jxR3oGX0/IH02DzhSfiBa0YsXOxor7AVINWaehjxA/WDfQodomue1dV5aIv52Bn
jrP/vyCRcRNK5nXAmJRpYdBol1+beCwuRZEDw84NYfAD7elmHeckgQnYr5ofmgUJ
RmiNKARAp0tVDC30vkGk6x/SPqK1P7q30MFtc9ZzN87HHUCxHdeo2S+ucYgN9/3c
HtcNocQvOpcg7lQ4jFs/A6cTl2JBmUMe+QEWhETWlpei7Ll5WvCN0WttTZIDFRRg
ZDXc4UPPCFooJZghCGG1KBCsuHCFOCOsOb50ZIOsBzCZvo1IvU3IH60/R407asjL
7lgB80y/ksZZiLAgcw9Ht+K4BpVpzzktDfcm4I3Anzyc2PtYYmV37+RSxilEoKxY
XC2amgRj92Ph7cHMWjtlQc+wKKJ6x/uMMaRvv8sON2dvMvK+thPwvU2kyr24cWNI
Y0cpRwgF6FE2pU7nxJHhRwQT8TjKjvMA6BdAfyDbIH1/s/Ni38Whky4iu7YDEAAZ
qoGb6DGJ4X0ex4ejIPvXUBEaYgyRV9O7m0bsxd1vrJhHvwE1BOM/04y5e85LMxPh
V65fboUR4QX4dL/KfkUlHo9TmAxklYJeqcQA5ge/MUmsDjV57KMSElKlQD6SqThl
x+hhvVsLmFPBtm/E+2B9OObh4h88UMfKcPXsJv77x0pvz0se9SxtslE46eY2RryW
UTzBv8z4cl1FlQXITbTsooMFWMjpBAXYYIzum4M3n2TTY3zptMbHtvBe/jnzVExo
42i8NOhZ5MQdHBTC0IktxPCuarGLuS5Cwh4Kik9qBUl2JcptJBuSonQ43q9Lb5Lv
UnW+N75X222x0BFCOfVgJNvkn5dpmivpfxC8zAYORAAig+BmPT/J0UvkOSCSQMQ1
iC6TUqIgNn96/k9tv8idaTNsFsYrFJjpz02a7iORI9BskiN9cEkB5ZdX9spthWBB
M64UnhTSfUfX36Jfmypi4iR2GYFl6YlTcXqzW2pdLIzFx1J2pINkMfstqi1sjNge
56G62fFn9l/PxiAbDLzbafdKBOzvY7/dktvkuyzud6EbJlqU6siSI9yt+cvL7AZ+
yKnP5eKx6vO4VJYxglwaqY52EjY+23K/LyPyAC8X6PEu1rS38V0r1mgTfwLKW0bE
gaP8DDfc17QggMlACNIImgl8EIelPmVjrMMM6IIVXMoNotV2NGZkcP+QSy0AXNcF
pswebL1BghHJ1Bho8Xyd6YCMsW0FD37jOonp/qnx1zeDC3xlO1e0cqMspXx1fy2o
XtzNbfn63UguoUKN8o85Y8wBKwyGMGLFI9O6qYzQunJYIrBtOR4aGbDUYxUa7wXu
R+Zvte5K0Z/K+pSQogrFAELTiZvEePOWpBKLU/rj+hLNcp4tYAchUTAqOHIjRGjW
0/r3qZNblQo3ZESVrEGA3H8T3OzylAw0T2KamBnWRy5ztdBY2n2B3F4DmNk1VKlO
bRAn2yMW39wn/aFq3l5bnnZYQw6cdN6H9zbzbm/ui6QS7rtVQ7zjS/xhslpJW6v8
33NFH+MwMuNFZlWkXQ1xLJJbpiVqXnYNgBfyyAN5ugzVa5tlWkZcaoG9PKnYYDip
YmEtjIkHTyDMW12wbWEyVDoVyHyohsMfc44lNQ1dcXHlkStxFFY/mpWQ1/CzhndM
AWguOwZ+WlH6YGXxB/6fHqYpmRc4crHjnVTeIXe7yOftLYMsil+69pkK9oreUroO
dIJR0MAfIV3QvYkN3nPSk4lvvw9rzN9iPe/yUvkgcHgGZTENRLh3uWm1610fGBuh
++s2zdaXoWzwCV5FlMk36hY3SttJHVI09Yu7XpalDslAxH2rf284ceLsUAU1N7tc
Z9ihM1KSw1S1hfB072yb5L2zIwO61kvnii7p70mP3iEcgrLBQLgeXrmb2suRsukv
RJ15q6dGYZR2G0nvgUMlL/0zK8GpeUiBfoczP6NnSKPdq4BTWmHgViHCQZt1i4le
fi5M1DI4rFX7k1x3hSm13Fn+six2S6QKnuJduT6ggPpmBRnmnWSJ0a9sXzt42h1x
pyp6ky56S1PuxoxaX4JFnRRSmaFhHm5y6apeEddrGKhyTmPpeCNQh0jBUiJ5KUrV
YadaIwnUvjsEybleR0y4CpkaQFtC3tzh3Jt2dLen3nTW5lwnA3jBjg8kTJ0pCHCm
xZRGmpLjBDOCViGNr42Tc54Y75LirxeGLbFfbf8wu7A8+YEYJ2CC7B/p1f261jh0
c2s98ia1y5jpXCxQVUaDpp+3cX2rCPd/qQPPu8xelOrpjMlEHXFLwq7gE1uwfTKz
5cr3P/zl307isn7ikT816yCZvOB+fQjwAjJnCzW93hgqx8rl5d+9E/QB+EB3D5zT
I6+dLP4t9/1yymLc+ZW1gbRX9DkxX+iv+FbxOWU09qJF0izPraIBKBBi1qjkfEuf
fXIV9fhwBuXZtamMj5g1pAnMOXlR5BblL1geDiepmqwMp+yiVSp03yJ7dkxcRGj3
0y5w9GbXIjgQKTDRl4yRtk0V0KBCWR1vv/E4xgfK2jFW6cbeRuv9Ekocey5qDWI3
OaPMo1MtLp0nw9a7xom4KYmrDCoPis3cEf5k8jlBKPs8F4/lYHkjs6QnMBxT4gQi
S1CnJwQZhx0en4aGQsBScO1/qW2itdHBKCRAX/EhK62bSvvAAgvgD0nnh9ClWr3F
mioGKySKSl1pFZHQ2PydxvkzZdkJD9od4ppv2ee8rQn0S8PHuARlqAyDK5xxzd9D
K2O4MGk0wyXaBcrhfjywbA17Cfn4YRWBYP6NtHbUDf4UC6cEdrvT9kSHlNtcaxsI
jQNDb0dnJsskRyymmOMz6YTa/U/xVza4KE0XX7p6ekf4rBbrHKYZ24CqRaYYIi22
7ZkxuBiO5SmNFatPj1n9Tc5K7Mnll0/KjxDoFNbf3Hu7hTPYahKDQib742TO98kk
VW2z/2I2as9N7WhK4dSURa1rJjK1lykKem/+ffTrnu7kYhYJK7CD/yNIRIlc4n06
m9RMKQ+vKJ2442SM1CznzQUC6CTpNr5k+orOiFKDhEZRmpm+jJocMZvYfkzc5IC/
Z9I+6ay3WUDRlgzJGFruhacHdn563hCXYrrBK43WMY3sxZcXZXvM5junjJFjABwh
3c63KOX5BhnR5EY+L6p5EyPAKxYkA9EnXLCs2+32GGtOj022XoAs7cNObMG4XrRp
WFs8bid6JWv5jqWT8X1X8PNPNhwaVXu1HftrnMVlKKthNA89emBGVp8ekCWra9o1
USg3+TgU4QMU1tBH03Mp2Jd8uAKleoprEdNpt9A72LCjFucsWigQ97+V29CF0Iqb
wo3HIvQB8FXRe9ywHPurFKQwOMjqWNDzz41sDG75G6h9UNzNmueyIzgWorRPHbtu
gY+iBG4ecR1SWdmn2j8OYRnDwy8gIDVymmPldk+W9hwPtwEuLydGlNvEiV0bqPBX
dYP7gifqQ9jCcrfU/yFwCZlZkKA+gGA6VxOMc+1NSYFZiYxhfrWq5j+Vr0mOgqFW
7CTobTOJxPrO5F8ul7cm7QNalDqf6HIjDxKkWgzPwcKsB8Y4X/uPFLoZgG9ME6iM
lwRR8AIrfoVt7NScRIve2rr4o7ZnAkYzbSoVyOGkb+VM1tGws9Lhfwyy2KwGSDsP
aqe+7r/4LjZYxVPeXSlovyZwhYFm6q7V/DA0dfCzjbsCuMhjnHlQbqLOgI6FHzTr
k8kfG4ytY7rdcx8Ae7n4/cWmG0mPTqu96xW23Ed4C+PwQcBYR2UO5xVPgDPBKiAP
1ADHBkGK+qoVVTnwhgwsrUNzwooKBGbvvar0zDeJGA+ur+h2x28zFfjiiDtxt172
tB4zksLi48fKTxRvu2dhEavk2sLcYqppjht5q8iaZzzmMyq2fGpRH4kb2oucYJsc
khgBC6bP7OZrxEnz6U1SM6eUKMAZawwIQVhAlaFgVw6qWAeJB7oHLCnpjFi6jGQc
m/l5LY/Ro8kOaF19eWaiqRjCDCprNHj6YepPwcv7INrauoiB5Eew5/U0h6vLN44H
eVC8kiaPHDNubaBGDjwJlfn/hyAS+42uw2V/FNOtJYA7i41QWHjHWNT79f/Okvl5
3DUci7wcRbz0sSnrPaXXjv3TGT2y6MhJfvY+PZMCtLUBsFnrwaA48KO2f641xzL1
Xocwwqo59ybw8dqh6qLgk+tm0zvbM+nACJKyl778XE+0OSUZcSVfsgGd4deNi/JN
sKTR1/+3Hm5Jbd66KSwWD8sW/99ehVtsqFijBpS9vird2OoMi7rT9xATfezIW41B
TKRE1+S6CZtFODpQY3qYBXVBuwGWizU39LQUNHy/4t8evmC+H3tpf17lSDXJ7YoH
04msqYJJHfH57S8D7xGmSPUWlM67GVjoBAvssWQtM7uGRBOyLuEGORCT/h9weuya
o0ldgvYbFwoEED+h1OjyrsqNcKJ8N48J3jk9mmcd6gDeCzzja6VyUi3T/DnG/Gua
k3ioemrPx/X2YyaqhgcnJnhB8i9G6/0DZm35BgKY/Ok4l4BWR8q5EuxL2LRd8kzw
vMyVQkVAqA+00up4GuX+IW0P7pR9MqkUeVFI0CKAKn+QI7ywhIaMgrmMRc3FlA9D
XWRyzOAjSaIskP14ecE/exPonMxtFng+FDf5rgmz+KhzqCn4JRX1mUkRKD4NCmJA
J0Sa5MRM+TD7yYwunK0TlrtLpd7o9mXX+rMgcsiDXbh59fxT1pm0M8A5WsJVcV7j
VQZ4B86zEc55fOClGWKOCyPoLRb/duQZ6PwE1A68M4Kk3z+wa/uvQnCvDc3ie8xe
0b8WAe9n6Ql+x3QmGzjyqe2xgH0GK1TjOL9RDPrZjwEe8cOpgLdTPQbMH9qj5aGx
EAfWKODRQCzcc3D28QG6uUDDrzKYcjsbmHdV8FH1zcumwD5FMZU+kh1X4kpXZQLf
F9xRka1O/JASKDa4TG5lTElcPrThkeO/OKLcIj87Hp4puCaHSqB7Ic6rNE6L9Ltd
WbPccEqbgtL3ymnRnhPNVcbe95Ahnl8SPi4t4Cti4HIex4nQcoC8G5FNkJtjfoL+
3OHiLbmoSe76P4VRIj3Oxb3VjsUmYL3PreDOgy5+lcDXw72zB97edjRJcxUXqk39
rk64AAJuOiCtiXULp6PeqH17EQBGpm2fMPvJDWsDvkaK7TLIuxRsSfpps0BTEMf7
SsojDQkNzo4V+uYBGb5wh7TfuAhwJVwIwoNOsR7j26VWudZ8UwvZ+zHPPRKYdMVN
XASQltxds4Fx+HjcNKmC/0bEr8KYTOdtCTHKZRFNg+DGVZpF9dvhpBEo4oFg5SBu
8KY1NjjLx2A0AFCSRiAyBgfGCTIr19zMLXgARnSkSNUfJSQUNRUQlfuWPGTJsbDX
m0xw2tGk4E6zo/bRc1prZ1c7S84UKQ9uyHJvJvs9C2SrsZxeclF/gz9angLvixez
BLOQnw02t8PQt/sfgN03ayCvOoLtO1DzjXAcxeaNoRBC3OlPrM4JavV2H23vB0Ly
BL3CbU+BVDqpolQXxwuDd/RV/n1xyvsVhcjTbWZT+aAwhUPwYmicwDP7sgmJz4xA
DKLdTENZ8EdmeWsWO0GXL2hJ5fSJNCnZgAWlNbsT4qMtc4hOabkkrBjRjECVWCFr
du3dlpm7QkCtPAmOfZ1cBkJZQJ85mZBSilHPi++WgN3EjTgzs4yelkX/952+LXXh
6lq3g3rLGT2iZijiDS7kP+E42OrL7dp2snbGrgK0BFKPfMsqZLhwA3wnQpqk2YZT
lWElI0riClWrtRh4G/R2fQFKWjfUzRMaTtAKeu9PK7t1rYiGs/dq+J4+KEt7YH7X
jZfc/rjeJzY0N+Ty2cSxu9S0fXFGymaS5s+d4Zw1D+85G/tnfLzf/GcJjPAgytO0
KH64dyldBgT0gPLJp2MyhAihwyc2JZ2uvuwdK2Vac1+8JVJGZPE3cyRE4pXdEAeu
Qvvme66MIxBiy3BTLi36+ZfLphfaB0FY/ItS/upSVBdNic8nqD1tkj4xNHZBCl6D
8czbjCVin+eII2K0B+TqnZeFPCcpQ2OBjS6x2aLXCw5kpKSti0HUpES+IlZTc3Qq
aYDxkkJyQjoPH7bmQ07PQ1vUCLlQZKmvlqO7i9byw0dzn/wY5HRAXzUWGCpkXG7K
QY1VqjWY8K6cuige/5k0D1Xr8kTCTgMdolg2NAO1b+bFn594ThevmMM20xeWKyip
1MnfKLeiTuJmnGU7v/wMWp1SqhU2QPfBP+4AVoQhN2kPgvxx8w1WUGZ4C+srEP98
r8Dp/uemhfD+XLVAtpnqazphDav74PsflGRMwVy1w4VvRjS0MKH0Qy/VeFZEBkOI
yx5jZ0J284H0eDtpS+OzZPyXm86b/Wqt3aDfaM3pMRDVoCYtM+h2JBaLK7D1a14d
Phz4L5oyoHDOxVTKvDBvMZZtO4Tz9sg/Q0MK+ayDQ/UlxYwJKVgI9fhrUrtzrJ4w
zGVtBoQWVZVhOwHl/s3wyEK9De2CnmiT+QTTz2a9gqijvysTtMYpdc/8+nFX/kl4
xo/u1+ItvkwAHFzBbW/4MWM8MOYyJXExz9g45q45yU2ZVLPHcTgSGzu+A4lICbw6
Ze7+89w4kqCe+eiJAQBp/swIHRFvCGm6MCgVpU4PZQfWL9ur5G2LE3i/P0QJiaMS
UqSh3MY0PAjNRwo1t5Aq+od+Bm/twrReMUe8RKhLDxAO2iur5RH05JTHr+5udaS6
Pz3YRLcF8PVB8J+SkkMcI0Ftqq1HEe1jXpxU0hS/k6Z7ZkQAHfNMiaxhQgduZrEb
GZD9FdrqkGHf9x2VnQvY55Dg0AAMojq1D01uFEBErbQrQqt8NgyckKZYP0QmSv8S
gO8NwH0Kt8rLyM88n7Ckf6nkmpS41BTJTdKIsTO/V7+to+6GJ7H4EDUtV3AMKKY3
s7KjqVEuELFV6FEMR6TrDI3lbelj4rI+bNUC5BKbjXAV3m43VBvEJk9QjE0WJf3l
E9Vtm9J7q9c/3/YwWF/2B3R8hBEXptoGcqe6476wj0hX6uYRFv28dqHwieRJrGbU
rfhI+frG7UoWBBSuA3QSc+ZvMkeZ11jTilQyJ/H+4C2qbsI/HlPiyE+JfOq4Iosm
wuiJESDMku/q61UYNkbrqiqhy9rB0cowohiHJBl4CfyqBEEN5P2OjPi+RTp9vYHn
Eks0h7PRDZYGTKma49+tHLtO8RX9DLIfNqw19mml6StYa8Fft4BJj+QDkEDA9boe
WUS4zP7rEkOL9fiiENe9T2RUAXVFOox8n8OBSkWuqPOL87s+RTFPRAEmlddNqiPA
nibUrSotW656Y2uOMaNrt6FlpYfvr2QKbraRXjtpQedzL55VSzP5+1uV+FN3WFIk
Mg6aK5HUhoDISQ+xLTTSt+UgkSjZrxZ2tZPUoz4GkAqKCSg7V5BmRqiUkNi8wsUP
Kzzra2Wqzxy14nsiz4FQPzR2n3ZcTBg6RJV63EowKmea9AjSzF+OJ/2tusCDY0Ck
XLO2NV3r3Rk7Y4MMDg19h2VnuhrJvR48MkcJCJztKAmWWP8sO1ZDCBZDac/lXAe4
AKGWMDP6X71hwGGEbCXAaYZgxNOvvD0peISXoAHfLpxFupomdxhhCicZFY1N1llj
1gbwBDJG2VYzW5QkeHsJaDrgELvPqKjitJU/WgTiPfvFk4f4gyzxEHNDhX3U4aMw
IaFN40Wc2p3k2uAck9xlJ3fC/8XexFAQuqxxKJ1y9EJ8O/1dxZUM1yEpVcOoncPC
xqKOf4AAOooB5ynrEwzvFJDdRMw0FCf/BALHzP1caMMsGtzMKxSNC7eKCwCck2xB
2yoBlODhNOq7Zgkc2SaiFL2b03vK8rFHPGsg79rHVfydN1u0iVwdLGanVpVSq6aV
Y17czYy8OYwOtxdwZt+KNZTLzQU5RFchbwT2bw8e0OMv1M55SrtNa79LXGRczYW+
KC3N/7G8E+gaVO3CwJx8zjmYZiusnG1bOvuoO487qWW39+BSA8dQTOdCAbLVS1S8
1rEAuf27aSIdsKfQFFGy3HXXUZfz58SITvgvV8G6O7otGXnuLBTnVFKpYD+xcBFW
KdrrM5Y34oa78lqidkM4sgocZOz0RgRoJBiPuNAkwQJP6hY3OdP5/DXFY8RAOucs
4YzMMKLiYN+yrXSxbI0ydrp/hGfS5fRxzBQ0w5xLm4yt+o63USeCw3HREirGOaMX
4PpLdn3hIp/d3FeUGiSEgSSKRPm3+SPepcuYLcIblUIpLHA/npoTZkt0KVqK8MFk
PfKWN8YBgOMl1Ifl6y5zTGyAU8ZyPUZAG0QvLoBzyJfM3NKYt946LAW0PHpqnDD2
8OtkSOxbvYIgieMDD0uAAO8ZidYeeTUF28q/1UWE53RGQbtiwe+3auMe1Tsfl5pH
aJgfrRssRAJcC8mLWqGQ+lr4XnGAYHQfeURJKtEJo06rDtQdv+RvUSjWq24kVyGf
YKN00+9DKFFV5nQ/7esj+qqPoIVF3MQhbXIYa5++QacalPqqFkaQNEhbFXhb+tIX
79XSzcqDsFsCPnMqttynWtmAJEkVQ+BCvGRbCpBmhiekT2+r01OzR3lBgoRL3/8p
foaDXKyurXJhCDYPm24hbwK2wmnXic81VRlthp7esh+yr2kOiwjVjXbwRJgEDLc0
tMXsZpKm/Nc9cR5Lo5OhotNXrLXOQPmIqaEKD18pCF6FfqUrhI6L/9it1G6qPgXJ
TCFRUQYFLGN7mippGQeP9pYULReGNzNglg5b2WlLf8bB1EOH+fo4zC3tHqeXJA1e
lYf22dyZ5IXTV7XMLZjW0vogURQlBPlN0SSclg4emkpqqZIE5tdFCNqLS8hZXnHa
2ZBHfIJvbZJaW260U9YVFi/NQ8gPAOw1QtHQ4cmPUXorkP2pQEtEVA9KIChqtutP
RGFN9mKLCbzsBGdXqGuBDjnD2byBEjVtxHylem+n35a9ueszO2b6bYo7e3O4titG
p7+RhX0ygU4g5hG/SFMqRXCpKbQ2UQZo6JzB+7xd+Zv8h7OqzM8N1lMfm6PkUQQc
TA9z3U1L5D0hlkCqPX5uO6qepybRKqqNTGxL6ngrGMomebBiIYQ/akCGns+L0zU4
XqvZuBoiWZeKHXzxzlqVo/nMRsqqXrkk7OG7QWH/ayaJGiIaR7YRWmBzmpMx02i8
lBZVBXOu/Goco44zDrZ3zVy3oW7qvaM1uBSX/7TcqapYrVBYXm/F+wrRWvWTI+KJ
sKuIK48KEf4AjOndbdC4tp8wXzoz0bWPegQCW7Wl6WmwnIvt6DfdyGPJGT7hh2vj
/5JYen34miIckn55WccGkNukXEJsLvWp+0SbU6kbU9kw7yNXN0sW6AE0UFGVI4jL
DLasfY/kmsn6JgOkDdm4EEvoTRiAGrm4L3wKWHYhQ/m6hYjs/+mRKOvPGa9rxh6J
RMbc7MpAVHDsHOFcD1fR3YNxCT8+l4Hl8iQ0xinOAtJ18+oe04BlfcoooDzdgr38
W9gtn4rmIQoYD8y6yKwZ9IRoLM3KlQos7CZcTBe9w4nmhrvAVxBezFooTaIyWnHL
OrmJ6/kW99EH91v0N8Dvtkq640Ldlw4Fdobl+T1xFG8cau5rtxq4rpdxp1J7YZLB
opUxrxedNoXXVE05K6vBnYJVJXHr/iDGdBzvxlaZhZz5CSpwXx/PdXgCtB4qjoCr
xhhObHcdN4wLAxyR6kWBoxmEInOm9o+g7Gd28vI3P0mzj9yuYmr9JzG9KsvRR4pF
htHc2UNqkUnyz9z9iUxGT2g4OvXfo1buGphwzzpxNvqsTDyFC810T27YkeDJxknE
ssWJY3le7TpysmQoHBWHZuEWSu3PXKI26/UMBPT3/p+CC6ppsK0MMXaW2wm1A7O+
PfBw1Fp/3vwSeW1XFLUFGoZDWwthsPKWbJig7cFGJ0dhK386V/HA/PrGVL6B2kDS
YNVP5hUxn+Pd0/HpstUnBRCNEY7pDTZhFOpBNbsMdBwBd76HHe9tA/qBwwUk2zNA
BgFu+EyHmp97KMMHn8K1OFP7bZtzsJKXFdQpzuZeNTSA/azIaLkbk4LOtd/JXgLy
NWtVNr8u+4ZoSRX1goNC1X9+43qEmW25iweIsle/3VXi6s13oUdBbT55taEccK7Z
zwORxD6F2xjVND9Xodr8Fx3IN/RMON+Jt3gy7hxbAivgC0pf4OqZoczYliTtscwu
2rBXGrNX8zJzxrRV/zpYG8yVeF8C0p+B8tbbcweZkzOOUySa7lmrgRIXP7cNyKII
UbRn63Uko7bxmkfcE7FMSDnlCtFidCV8+dyjE4uu1Q1ycmvuJwoVh70NLlq9JnV+
Lo+XVxXMvgRUQn69DAh867tRv7RCPz88W20XuaUmAaIB5Dpb4Q73P8Rhxr8io68o
ElUx2azg71aK/LO1qDnHzUojLIG6hUBAa3yNJA9KghaRFtSJKaqsiFK4itY04C2c
LEZjBEwDwrE/InQcfA36vzbWGbWRpJaFzJPt2MXIv0Sb87r35v+2TRkRSrIqecZY
WgEILc/WbWI6rsq1zccxNaqjMktOQDawXlSw0DQbqMbcsp/dP7AABSHiN1umHL/2
eQw2q//5chyZMIFI61/u7OljTamiFRUV5hn9iQYfnpPk+ZucH2Nia2kPIC/OcjuQ
xWRT5gt3EsJCuL781ZIWuIAWOUK8SwLl2j2Yli/5yIhLfrC1xUL0U62ttHAJbWfL
V9OIN6IRlWZLw1xromEGTq0RUfZ7juLewZpVSDD04Ftbc58jULeC5VlIP8OlsKOe
Mri8xe3MtUJ6+dBULZmSNUreH3vs6u5O7jiMqFcrlogs1cVb8QmaWyXJNAjbPoBq
t1/KL+K2mDPR/p2DRnB+pCrsrTrvamJ66mX1s7+axVPu/LOSoCZErHbOY0BRW6h7
bBcpZs0I/a3aI8/k9c/S75K/kb76dFssLWpNPxfYN9OMy9yh4Nlkm2sL0Gq8I8pL
dVfhm9UdMQq9RTFwYFh57Q2J0G+PPCde1En6MJloytlb8qM8sgkDsZOVkfgVOKkm
k564IDEJuu072zrwn5muUxfksrxud6QwdXxaNAXJPpAAno+f2LwFlM/73tNRQmRW
IpnV8wiRazOSs2fgVUFCrIY5pZwLXHa50hIN8+nkS2J8lSsqlr1UtoZVNCj9yuc0
LzVuyx1XdJlyd1E5UpvXsz2R7mwNAucAuE8vi6bMgtzG3Zxf5iBxVoUZq1S/Aula
RUTCD/K1UajZgZJ6K5ygKeJCXLyQAsj+JskiNkvUTUHgqMuMeDVPQd7QSxlqN9lC
NlFO747TqdW4/VAOjxCtMnV/sCJ0EK10Kd0lZES9UsQqOttgmc6LdfNpDSD/+rwJ
4Rl6V7fz/dyVSpVQZQcxiZJSYykUuPCvhMM+amqLFv7Digyljk+ADHiTe7dh9/Ev
DzxuZtgcW9YMU3p/HV3Qd40Ab6R2bnFt1Y8zvOsRVbU0fRGJ95P5Heqw5VpoY35k
LwiFGy8iBDAFhgF4c2St7pOPl67HZ+ZX2dcY8XvcfxA7ymTQcIQSuww56ld9TFKp
KviQdArCFsRCptZ2Ixr8S5zDQRpXTLhUAY+OsOGXLbHNi8sZ2s0L3A9ASqoEWh+G
XjNA/iuhDfk+CqNaVUk0j4pKvuCDDUdHBCE+GtSCXyvc2pVg0xtLIw5uJLTBtBhJ
myLd3aHUNlJ82MvgC408GPnt5+20XlhsthrlzFAtepUeHhbjSGaqExVxRtSYOTGY
SVoGIzinHSL1oauAM+Qwx+noEphH7ekPw3Cj8N52GmPepnIO0pI5nDy4eNGfXlBf
qSZQo8hcVSc95L/7IJhZlzZTEYh7oOvYd0vg6kqnK8gneMU2TwmkJVkCClC4E9G0
pS6ujKjGjKF3w4PNUTXnUTyu9JI175NRFqCLXsUiYJxqtqkTFW369DSTeFLp5AaU
JUUu63prh+BGN0JCkEfeStNFexfzUXbq9SvT6V++nTSqK/2EvhpgJX2X3bhihNVx
mnicovr3rqkM4Ez+U+EtbD/rQV6+zcDK733LN0ZyUbfWwOTYwNxZU1T+h+7l/J45
2cmvCGNa+N1Oj666k9QOYsOT09hE3MfYthCHsKoKDLh+xB3Xdw6y3o8VWRSRaE4s
lvmaHjloW3SPKDu5tSec0siuU5NGhTdNsIvqT48JG/UJS8va57mcAJisqfwJraRP
byV16Sr5F/47pGrehSXXw+QW/BCQ6pVmogf5F0OoKe8mUK67y533VWo8AgrQP03R
br0svfkMfZKWkBBiN3G1i8yXJFVgBFHPLL62RVxRDty0xOf+OPToJ3LyTQfVhBN4
jLaH3DjvlD3El+wyG09vKcZW5dsY1QYfBjDmBtyrXm7J1iCdWdxvGEfHQ+6OMWLt
snZUsKGG2OWPVaMjGhJHZRESKJDT3sOeF7HP8YhNcjBu8sDgptGkEcX0mLYCvbJq
NcPjmPPU+E9ytvQTv/gzTwnYhRodcCz9kfS0VqUDPa3GkfekBohR+bHkItXnYNjT
/1yJVWq4uXFOXSyS8uBye2gN8EoVwECxnZ8PJIPPkh1Csy8EQ8oxD/VG/v25O6Om
Axor28scmLZM0fNzrfG5moXY+WKHH0MTdO3KZW2xhc5IYD1QnknxHYAY0VvsUn0L
wN4ojl+xVs09kof6VxqZg5hOVi9v2No5tAAEtPKqMcHrV+/Jd5KLI+eRnZZxjyKb
K6ruE6n79QVrgDWeVLoDtS5R3hlerRwkKmJuW5+rOqmTSrVzkpI1EVzK1aF6U2aY
xjQc7/kJsU8b+WxRMerj4Tc4RLNCf+cTA5dgtEPw2Us4y4VuwZK/AzWVu2U+zB1R
x/WoHF2e3J553Bsyvvs5qorK8ofFq3ZaosOJPH+FRUzSEa/3pN7jb4SoF347uSXJ
rSOncg4xHgadJmuTpnkxE+e71WeqNfC5OJ18HVeKMyoiKhf9gTbZTeX5fd1MaxIM
Fp26GZBfYveAay5eZCo0LHiOCUSnUmjDtHc31ykv6Vge615g5bTyLly/Jz824vRb
8tYaaO2NuygUOJnJ2qjK5c2D6UwPYt/QUqS4t6rlYLYXLe7fb4vHW6aFBqyDjye+
0taVRdSz7u75mKgMz/kMfp8tpnDhtk5WvV+frrjPvlkelPyTi2x3fhsDC0ENqYRq
EzxUZSdePwS7H2SlXjr7c2uuiKQoQyCtNNhsaYrsWoHzYzyhaaBwub4+kKiEN9gU
MpiqQ5F++YA48tdr0BQLpSxqOp5BTfGjPl7EXVCWNQM6B2sqmHSrtzD8DdyeM4uF
Cm++eHmyKDcBgu1xVhb55dgROa2i03tvCNGTv94UapWfxYnAbWV20L8F/x7DGxsP
OLgKGBBzFSp53tdSLp/xm0SZKYoe9DYR5RPIwJJi5mnYb8C/SWlwagFrxE366bEC
BPZTGv24dEHEGPqgTQBG+sG4c3gsCnObAE4aSZnriWrAGg54m9U5kWBku38DCzIE
fLnxfdtxIaGiZE/rN4LLWCLk0mHWgNTU8xU+BeFEtB5P5ktq4JvFNNpKfPJ3lc8j
ZU2x+uK3cwyixLZR3P9DBKpiXKz+JGhezI9eyObY4LE05Mof2RAOkzDZDw9zIceD
53jmT9JzjBfgxEL0J0mHAyARvi3cG+I8T+LnZI4qXAckJ3bWhVC1k4eQFM+cAPAi
gV71mJI7gck9DuHuvxaGGYezicfNgJ8dwgmjw5JWMzONoN8nR48WRG796nTOrxAq
C7d3F2rhVK3rg6dFs0+Q+JmuCVjLzSCn4qV2VBshl0u5gbcYhesOir4Ke69bBu8Y
zQg1cUXzCLPCbPsUbmmEjEAUzyn2juvsaeBWxcP1Abay8JZRqQw+xsCcXicmm5SO
CCib8vSYF942/DiaBjvqD1Fk0i3ROIzW2CKlYXc1S9vOl7AOvwr35PwwPYxSyyxJ
NwSnCZzRyRWBEKQT4EIVS1Mi/BYh5RiSGT6gzjUifBN50IX/M/lOXUtYQ827N6Rg
fFp0u7kW44vLEpVoNceMsIAAiv5yVRKu1okNVOhWvP0VWEpgUMO5rHM5jWp0f3qO
bKPQoVuSFjngjeZrzuloKSit6bjrbGLiHJkzbBg9n66Txf9Zsl3MQAMTxDl8JewW
ky3CUj8ElKE2Xvogg7asPa+5DMU+gH/+cmfQJejF6k4MIVrlfhWHTp/I2D6++w7w
IajYXuO3LpHhq5gOs4S9LV0dqWh1ZPZACJNpNgZx89VEHkbcpDXnoxYQDOnhKtvr
CRQnGpoA5ywUxkI1/4Rqd1dKLjeQjBHKZnAjMmiHZ5a+eZFTN0OtROdIv5kRgu3q
IBdA1vn7slKxNas00Ky1mifFqsPhuTCG+jfDS2UxjXE8QvPJ5M58nz/elqmKBR3D
J8jO//Qae5hFbJfRbyd5YGNlMsRjfh9ld2xTbYx3RX1xLdvrZsHfjFDfjGc9F7LX
2sSaY11qAjxwgnMMAUzXl31mq0T+IrI/0qkRgWNcYV1wKMCmGf+dXwGI7gZ9cghd
Wjcm+5/fU4exUfqPTZhG2FToKsK9A1SNz2Yv4AZoHhxSHkQh1pHAjCJjE8ZSZAje
tXt1kyDIY7W0BMWzt1CyTWbc4bA42lr2VWITh+lxFouEcX2kPdW4SDauQ/tYR8UJ
jDUl0EC80S9FKN29GHJe6Q70WWvs52tFmpVBPH70zKUJI0f33fymSPyGIhW6nXr8
wOXHLQLqKpsTEs7xQWWj7eJzEdput1OtU7JWyjh9aqZweuW3O/huu18Lbl/3H04/
VfMfOhyeEcnvlP8GvjDxQEWNegFPrqqKIfIg7YgF9jGbUG6DDWrakARnfi+xbW9I
9ztCeRb/kN5mNo3qufjKy3WPGV4weTP6rmJWZslgHyUlDCLWu9hWZOoX6CVmW2R2
9asZxB2obAZ4bYvBNNFLKWzL4FPI8ONw1OLYBB4UuAMTGW6CWNU5K4OmNjJGJPqc
T45z+NxlmNPMj5dhZ01x4xyLuSeorcMtAmuKW0Xz5mGio7cJ7gbdJASRuKgKgnf0
o1hWpVvQL65a9AXRU1X7ORSUpiKnNqhTWPcYRqZfRDGPvw2cOIaG6UINIGYRYU3L
ZI8MpgzRYNRbZIF/48KGkxijOyulCDWrCTSSUyKfxvl1ggouPRERw33KPaZBoxDu
lb+BozwnmbaDiv0jGubY0uO0zFrsQowg9Mfvk9oVvZSbuInf7OidVHqto40ZOzN5
HaSV7Hzp3nrsPW1WVVDsZ8wswdDIGzADdaHD4LfeF02xXRh7JdWQ7DCWxiH1ftCc
pNHrFzPaEeDxsys4IDr3/ZfpHpmo8y6aZadZ7CwHlGcfhT8TWmKfDTD3FYNNuQx9
P0NhwI1aHHjlVpTgjQiywpQPaa1yI/dfuuj+g8sZUA3Q4jSrA6Am0sgLS/CslGfK
h2IRdJjcOPJcdsV/2ymuiAV5N+HGuOFS0f1aGOjJYCDHBnDZVxDaLqX6Nitmzmb0
xxxhoCIwCzkoY0tAMs3hikZ4frYRzKY9drohWWImSk+tJo2JmZ0HPFLmZg7EHhoB
OryxkZigNY85NlFgxDet0kZqW6RWucYRAwF82ESjTmDOrWnxqlRAtJkTDkWdQnx7
0++GR6WpOxOvBuavta2dLRR2SK2Utg97efl6nhDThGBSk/4jzIQKk/6VugEIaYE9
5V2Q2VN7ThZq6eAQrbpj4VEBw+zcF8WVZJx1qoFr5qeKNfVd/q/RaPY8ObwHmLem
eYa6p8vZWlK3NJ8uLu1/aZnzY28WGjrF86PxXVgs3KOFWlHUohpiozz+0Qt9H5y7
eBd0mXE1kHONrpseMcBuWdsBAd8h7sa2fpIxRahIG7GLjREGCOTceWjf/OYHm5bT
pQyRndc+x9LJ5PRscrk9p8ZAMdlLWJj70LniLMTMmM5+TVS6mfK7oxsY+dREr+Xj
HwiAKxjlY0L0htQvzA37jxCfc0kKkyBeEKwMarYFy2+k2G7h8wSGcn2uGABCqTZa
OemHRcJsS1RGp39QJKzDUKjt/ARSY+5BPl3oOESGmJnMBfdTjwYqY6JbnhGyAH7m
PEX7ny4z+gmtFJ7AqFfIiDEU7dt7V5aDBd6RcNTbhVzSCPV1nzWVPN7KuYqBu0SW
JsByl63MhoMNpBsX+mxWSvKvQmsN0w486tGeqxGZNwDGRolw95AZq5DQktPC//hQ
MV8Fwi/8LTGiAfRQ63AHJZoZEqru7kAee85VMe5TNM3tgcFOWlwhtDsdtTY3psVs
xgAiKObKt+vAOphQSLFigPG7tuuomENQ+37LiY1Wj21WCsLkCiUXtKQCX/RKao2I
UaD/ewebKpzeAqYTBtmKNQ/GjieJqBJ5yGfHfcWU3wHN0m/WaLLyX/bsZDedfA5M
RSxbz8oYoNnND6PmAQQteuU+2SX218GuuO7ZMtkXw1lCFYghefMI1Jx5+fwAuHa9
n27pGv/i0rUvH/ywphfe+U6rDnhgCxOCN8qzfMxXxpTlDG/vwwr27VVmm99PMs2f
M8xXyxX8XOp81mqr6QQug75r3qqqvv2wDXBFrScuKCIRaDnUQ05kUqmPyBOy+a/k
58xnzi5xyfHIL3l99++FTA4qYlyGmMMfm8k/dwxNkrXgzdfCrvw1+0kmmtP4ZyYf
KPSC3OCBiPije430NFbqssuslvFS8Ch8TqNS+Wd3VHmIOeVyNHNZGbLIWLc8aGkv
P0UymaDfDnUSWeBEOzh+Mu1NG0pMKw0zIZKKZi9T64GwQ/o3HvQkxbsBb/UwditX
2p9gJuMwcORQiWnvgfCvdX0qeIn5FXHAhmTOWBlpZp1sgepv4qQBBuOyR4UvA4gq
8x7vz36YSwrfofYn0U3bzq4O6yTeES2Mua4G7K0ucFlvUxTLUenKR0k0TQwgUcSz
a7y+50TzktYQd/p+Gd1ToRXx/RD4niPyczv3yer5MsV92G6t1zxYDNtwKvhkEwww
eEuFg4WHnhdAKAxKQpMkQFbARGOZhPq4cDP24ZhOKgmoKTdbkVoB9qIb/icLC7qP
8ZT71tzfF7gutz1jOKLvpVS8gjZRkR08ClMZnz0A1ClBNqpGm76nVuC1CtKbHVp6
wec0CcmrYJGAw8NE2KGTfojlnvn56KFpTd1q14jskQ5x7iblfMPTm54LzrYqXBhh
JPwjdyBCS8Y3qPMpXkMpQE5cbNqmf1Vw5aifLF/KVpF92YGGLrisvbliV4d8clIC
pirLfLhdmiULGFqkCpq/5XoscQx9Go/FMrkcQUF4XFmUqCchtlaX84bIDZrAizhq
c01NpF104DQLwl+Ci8RbfbYPoPXBdezBmfBiuwbYNBx7hbFGpthovFeH7+YKC77m
1/QEfO8mOj6fdHwsSKYh/TaG1IK/TQCzipQSytAuLFJtBJUITRtchyYDEhX6oaEY
Dy+v/lb9M3ViHudxHHzhtbiszV8NETr+JzP5F+wcP6PkNLB89mnfzrpWW7ZtcLrg
kEWvPid/o3jP+rx+z1hfBGAHvHQz1H9QE756m4XlBN0KQ4r+Jax2NkSVVIWcVSJY
QHIIvO1jMBOV3zREjT7fSOmYnUaaHMYuGYdnZMwN+nhdY5DgmQodjjvSMNi+Dc1d
RMPWq99OcJPIDZrMkhnJYYvUw2JdqmZeS3QcImwNoHyIJSInikY07saN/RrgoVrt
7o+eJ12zAzUYyIwe6pE46Rw4xYiq4K1Da9R4oQC6SDze9BhYsCVT7xJjkvuvOD40
sam1121sBj26UUV5nNd8JBY8qDf9wO9yv/JSl2Wb2EC2dkp/SaGkMyqaU4sNWiOo
kKw7rQaYFUYbdAakFwYKozL2YzKBCosoRFf0Lcnyvmx8qR8RxnVXnKKopecOWkZ1
wo3+39RVuz6sSESVzmLi7TpR/LhKeKYtMjaT/TXPfP7VGqZcrEfzo8ZPVweWT8yM
GMhIQkr1KaUBWgqI87z2nmrCK/kED3KZ9uQQiXoW48JTfJefcYXYTpCEEoroMYOu
NzrAwJ6cIF+2GvDKC7p/H5/hnAWMXq4gDaBurFSE5fxTHM0hkEAProkesUXH080O
omb3usllquup3hO2g8qrN1lT0BQMVJo5hMBLg1MnA8vfz93BIsCAQw4yoCeSA/Mv
UdPo6r/D5VX5JY+o4xOipFReDMddYKU3ToPLRD2aR/ST0xRW8+C6qsJmy07knqeb
WD/MrdneKtKfSCORmlTJJFivHXvXX6FnQGo4+JsSSMXn/0uPq5bEu+XAPXW19cv0
yt8x/iFo8fiL5pMMJpTSoJ/dX7DkYbfK8LDDyL7Qbyh7vql284eRUqYzrTcZIBWY
mgWrA3vaNNIjG76cabLeYCIV1Yj36ShERcLUhSuNJsjjKhd0vxZZpOu3PEc9BzFH
90wqPXnNddXsIC8ouoaZDBuyTqmLfjt6Vl/PYcgrH8dT5eK+oisYzpKFfdNDFrRC
jukKM+wX7iPKkDvR+Bz1KolApXqVafZBXQeOYe6ACCW0rn+rEDMXLz0YT0UQtp/X
eig8FCusFcTEjdvgYHtBi9BRCqg7a1wZZtp3j7LJ6C075qItVEMu61CxdxB10M7l
Kz/WU7GH8sqcDR0qhdUL07/l+mKzfFZzjHvKhdbSViE9M5LLXpigRKGSPTo4RzxZ
G3geqUC7DPVPoWSzXmayh0/7zMQ6zUaYWHhDvfkdYxdciZuedq3qP/eE13U+X2xb
5Z9zVdo6tIRCeNefr01OZem7ToiTy8LE2MoQXe39JMGze/wz2Lox0RNoBay3fYMH
eRSX9DDe/UFuzoPtdvpOyGhLLpxJ4oQOP9U1rGMecXPG9yPEepTUeafcLe7VO9cn
D2skNwPRXRU+91Mq9Tz0rc0jJImZiojuXGXVNN3wP22fY3hGsD8ojxOyVJHIogzz
XaNghdG4NR7KtPHMeA/c6KQe8LMb+vLDZ7MTTgT0OQ46R95RMr0dPIIsE3A4pDIH
57ZR0uNNNot3JomZB6IbUCpDhwxKd0bPiC8V0HYGS+RK0p9DBZLU/xcaxoK7rm89
WI0JFXRj78avi0dM0eiEPGnRqbjfXrL2T5IJNeTIkNAAuNkfpn/rZuHce1rfhxhK
kGxZf2Kml4c6tyyzX8zZEQuVgVZavadfH9w6vJ9uIsfcKZByNSxzG1DyLSJI52Y2
3II2icFadix+gZDsZXM7tcUclfJMLcWcW+/9JZQW/2ue1n98vhZ1y6mAq12+KEek
578DLgUH/k26V3y5C3Ny4jgAc1KpB35K7XX5454dNIk6itrcWIrcjnFULlP8bljH
PxxF+f3S38YkcUWbR0kzaiftfMg/5+r5dshCjuvklbWx4BWw/JNPNTiSIN0t8l7i
r8egtdK/ufcJElgHU8Pbi9CwrWuRrWLNt38WlB5B0QKX4O0Qc/iTmJQVahtfcDuF
uDk/dsIEUTxBMd4AbfCnayINg3tSxGxmGznYZjVV1zWdfw0UWkuTGfBRmL8UDQtd
ftj/YdtpwAgkhF9c6gmfwfhX9ouO6SYy5F7/8Ck88MSqVritgCs3duFdeYzU2tVe
zJRimw8BmUGFq768+wxFJMCLI6R7bHEbP4RFr8Fpono7LbLyG5DEr4Q4370xBY/w
mGNJqTgQDoxZWpRRZTMJ9d732+8SQpd2Wq+a7M4ykGZen3kJWdEMYj6+CfbgRUTB
yNKuS12p2kaJYVaJTLc3nbOtIOjg6tTEQDT4ir4Drp+vOrIadA+KKxKz5lBT4IOX
ifvpdTf6XvWlZh/LFLsHVPrQa5QJPeR4cn4SzwkVAOFspXhNfLYy8gbAD+h7qcbC
tqjXXNWlV3PF8NgZxHkRZfZfr+WAvDszLq9xneQ+g9fj1Wc8vYIgumrmHwvlU5YI
AUSJ/Ot3fgSBPSz28zgYqLuTGj8FTqfZqJUIVMaHqIB/PI4HzHX92MbZHtdajwsk
3p6bANo4eGCDlDgDnPuLeJf6it6NuF3q6JnpXmoxBzd14vJYevF6NN1BoAYWqDsD
pb8xfaz/JKBPL9sy+YD6lTS1Kl73VX32F1GHcTsExsBZw+I9OPUPHYcApNc3nIdV
4Eg46DR54gURvw9owANzbmCXvfFg97NyxcIhbI2gsfMMChicSGwQESKrFmv7Y0xf
8EkHKw4q9rhLIT/KUAN42Pc6kQr4OTe6V7/qs1WchFU7WT2wFX6MjvJWPBomY35L
41yfGk4biP5Dm1zMigFepFCySTzG8NsGWyaeR2kwM6J5X/5NOtNEnyIZy6o8R7Gz
CZutSFBqnB17ONHZUT7qkV/dME8y00koZ0k0TZJAa3Yj8SzHTaagjeImPu/FhE5U
H++BGlUijflnAJJAnYp86eEl7PHOYrW392KDpG3c+e27S2fIX4JLLSewCHUzdVIK
VLXOVUL8eviMGNFsnrHcNKnb5QCzhAV0p/AnPGWIoLc8551+vTf4XGchkTfjeEmi
Bb1qXD5x0Y3ONr9bspEg7T9EJ3f8Ui1GzcS5JO0eC4s6Wu1PlrHwGcbdZxt5kRaH
fZ0RaCFBXCnOjp43luoMzL+SfgZ4Gb5oYHtpD07GrWIb4T3vM3tdWvrjqAagj2b/
lRB0TYo1lP4I9j/YtoN72WVx/D0sg31xNKvjc1heIZJ0YCwMeV6rGFy6Qd20BQft
vbslLa/JV3HbaGAEvQXrt8RbNeNCAH7C+4SJjjPedLDBok2Wd70/luvGqRc/X/qN
MFpSbvfs2kInmyjD7XizvHLry8WpH4FqRIdN1nkExSG+HG9zxBNWahwuIbpo1Ll7
YYUIFzMg/PCAFNk47HXvnwsQuE2im8NVh95aFx9SVZpKf1xhqfyO7XnvKp1TfpN6
bHOWZe6jtiKHT01f03WWJkaDH6CMI47vI/CE98IjWh+g1JLlTNhVoE8KwpWW+f2k
u/6sIf/wjl2jaBbcLw0LMPY6xTGPYJGxp3CM4WiDLgPms225NLXc/Mi3taK3Qw43
MHSCPnnmj5NgEShuShqk9Ccxn92ebA920Xl+X2brFgMpA7UzbU8UL3YeIqTS6a2O
nbv4WVyBWXABdET9p5vQmmo6f6jm8pVx0HE9MGM0W2TPf80beNHA+2r44uBvsnsQ
ztbM3hxJJOIg+0etdsCKw9H7RoHTGu0htW/EwOx5+OnaryfwuKc6P36gBj0VuOnG
BSVvLPM3EnRntvvSFV64nkRIWYUsziu1KRUaKhbs1b7b+5QDcA+N6Q42lN/Qtx1a
ZSdfMNNDEIdEWyitNOo/UI1QWKqbuCx6MxYggL9qJC0EFaj/TgX3SSEiwrET9xzN
AQFhHn6rxbfBT9OviOnzXprEIcf+vgip7Z+Ud51RGzdnTzg61OXRi3HuQyh9XZy/
wcA/mBD1DZeK3UWu1SyjCoiJCrqWFbUkU7tLwZ30Ke1tfK+U1qWZ86d5ClcDDeY0
c/HGV+/TGLy6xfnOZLIARo11dIyIO5eoZyzZhaBBNKBXmT1VEUbKBuzTlJ9IrQkm
i5KjbuPYErl8M5iuWfrLyvGKy/0J5XCqaQetzxzGNNRdBxeCWn4AzVtPjAng8LXS
+v8gDiHRt13x8foLsZv+kcrO2tc0KYh5mnE1qGqOVETwK0ncpEDE4GSMzXsnePkA
jGhiHIZWRIzjLUq9sbpIqI6WW0gkhxjiurIPya6B85Qkb9cgF4vXkrD+8WtbJSAO
E+FVTkfXavj6qt4TnOw8Co00iERiDsPnTDxN81wTzA4MuPIuXTcM1E8JE+PJVAgU
jRukCBw1KoxC3XmY1Vmvv1WIdSNgNxZNeS7qsiy26Tvkv6ppTkJOGkFbg8J9Vjel
2qayIK0kqKz8xsrfo0opsWXQNenN1ZFu508ZU/nK9nm81GOiBvsrtB8ARIjP4f0P
W2FiOprukVIvu0sQa8ZYAeHodol9VTx8ehreeyiJdEXBccEzy1iXiKgDzLJZVx10
QO24SWRQJehXHovSS0ZCxjFLezRgCn4k6gK+wm21qton4wqwSyAney9YzrBEuzaV
OGBIP0+OrB4B+eAR/+GnOvkVJgeWwU4h/MVTGb+yhJKObauZKv9T6D5l2yhFKU/q
F01QO7p/V36DYfGZc6iEAWpLheAh2UUySav5HqqDY9cm8Ngs0rvcgqAskpmsEDmV
jEshMASSAHpjmGQNFJguUyhdzYKoDXNNCntRx6op20USdRiB6yCwj8winyIIGHZD
kdMVNE/lemufHw/GZZjElRA8PLIJngXnJdVxNKHmVZXOqi+1VqClb5Wt3MhBMNYW
tuKAUYzZJZ47+gs+J6hSNgvlEqMzzFDKcEUJ+0v9gSDPJQav9xuF1FR3SFnH+39g
U7HeDaMIjqtfW3WXVi25rqV5u9PEtLDM0N5qEyCSrXu4b25tZIYq7F9FUDHHYR15
HLjctqtNHVxmcMN6Btz3+e/0iO3eYCNvZRH4AQLueYJk6HMLWoOc/KOj+nI1YZLZ
qWeeEHo1vPmCGfO4dtt+8Q5raaj5E6uOO/u25vI5cBOGVhSoGZC1WtGONU+2EW/m
tlMb1AX+m8j8jwuoRvdFn6+ygh/21bilo45RzB1tl8xkmCvdW3DewEW6GeQy5ru2
nNYapOdpSarAy8rH4knqf48WWxgpS8TX29tZzlJhinGI9LZTKe7fscF41M0pvl2p
XplkPUbtTGRGe5qUEjJQN+n1xaok7CpJ4QC9GDc5QcfqwUuXoNsDs6ylkjVf3uub
+NrgkaQKA/IwkaZspzpMPSHQDZGtZFe85im9nJTrPGh4N8tYD8MJ9BeR3KG5cFih
DATT0GsObEb4MuP9HeTaM1GzYJsq3/pgr8gnwFJSF8eNAP41DT37KnORJTM+++L9
ywgoEwR6JP938Sci+/VCzCprXH4xliNqL4/1NYhZTRb3McsnDW/VUrUixbWNjm5/
WsMel8uYXleSkkpZ9B4C+trEWpM3SxcLRKSsqNQTatga2io03Avk3suJeWowmyKO
5px6RyCGt3rX8PGkt6w+K1OIHWKewoNkvugkiGIrhbO+hJlbf0dGFetXXZNOlmfp
iOrLkoDHggzSaUvED5I1vQdMmBknyKy+FnWLvaYR9Kjqjt9CMRJMWv/ECI4T3wA9
5rUUVYKitvexsYvC1lIkUCHJtnkkCl+fepsLyJoTdBUOW0P1XyWL0hvN3RaiZGLs
t+z6r9hraN3VFdpVah+yR7D/zhmHuSVYoxYH1uQYlsQRH1KLNb8rQaBVVhpOsl9W
5hEnOFpSwQINtVZ1qXoZqCgFUNPXk4Nr6J8u/ptGsCBpPhXMkKTZ7eWZoiKHTL7x
MtH3DDNNuJh+Wou72tDJnrzHnkQMdkeu8u+stG8kr8kGEaWh41k73V6yoYv9YPYN
JhNNXFIRG3yab7PYujjbK5khMZU6Id7QwAhrh4nASsnPaQFEzlHarz0hSulzfUnN
LTE2Hty060sskqeoMMGbTexYrGueHGkSms18WHppphjBtdb/rEd75uLd/F/+PXlP
3RMmHhgJu8R6oExfmtwkBfu6TpvQIqZHb/NCltPFUh97M5G6DbQkqiGzNnEDNCJw
CyeIfdq6FEiGsoEfPgBcVcQJUqbylWvelHyOm9L4t+KjXbV8G0i6EQzMUfg7LUsI
8MSelYZYH/jhGBtTZ9CS8Zn5yE8cx8HnbvgeTLmlUgE6qwGxMgZQMBAihwrTQzKx
MY1v45QTgJGCIjh+juFiiOboIqnaoQK+jjNfySswnQKMLaGP4utSlXVN+Ak1GE/w
dtHI1yDtDiocsCMVrlmDWIXndQkOY2iz8OQLWQyVJcFMXkXLjFtwRjMVPfSCcEwV
0gWvBwxcuL6FXj4pZKbBhCC6Rz4diFZvuBPSahoEiKc5b3kg8bH0/aLqhzj3+gvu
pZpfH50e7qvaQ5y8CmpPNip5KWzgIMKQjv/Qlce+9INn7zTvGXBpN0K6Ag3oR/EZ
ucvS2OdbcPD9Gdmt09Z6DiYc3rxM2DH02gmmbfcVmAz6CLhLYJP78DpkG3QHBD/j
YdtWMm+K36w7YHFivNCDAowDM6C828nOK3yy24rvxNwnkO8aRxlx9z38MlAYysuJ
N/vsZ47Rn0OZBjHlyswI93rTLNnK/Za3AN4wku9rF54i4RF/AwnxcItVCDrmeYE8
0OugvzwzM64Z0aEyCSry/t1q8ClDlGQZLcKDHSatTC+dLqgEgQBzuuzxiOk6DDHG
MLqpzqhthSAmh4svovcI1XvkKm3cqPAouztHXX+HruiC+jx06JqFs3G7jtbLt08F
ik+OBC9grfbrelZAgt4bT4SVcyxfBjSjCvGpibVBLt035qsJSMgKDOqREJAEUpe3
JCu1e3JAAKwCWQY8hsW7ophklrNq9PXs2Gyhj2W59PvSOORKfxFeKPkV4GyAVkIf
j3Nn+EPKUi/IiPWBzjYH7gDEqT3SXZUNiU/zxExc0i0dRNaTPeE+CGKPo6zHcRdt
f8tdTHg7fp9mZh/Z769b8Yvi463WVI+doSdeaPwEioupVP0Ck0PAOzf1vzzUzO3G
3dF9q0EdkmBiWWSNdnfPM4+hsNtxGtnACqcPfKs/hHpPjDqfZJaKvTe39/iVpGDJ
NQlIBJcRUU1aC2OjUMVzjA90iTG5FhrW7L+BMY0W6AmlawLha/WnuQO6Mp2Y+kXo
wgIE1XhKr4xICnd5EiHRwpO4Rq5i0TY4Xdt3UKSU5I4G60LX7GStDOI7w0dcz6FA
Vb5+7+X2yVby16dARIZl3GnsaB5g2lwlfrcRv/jUUk4tMbNBmtLewzCHzejLQQ7a
O36MbcYlN24vsYQFzjMBAR+h2wQisq5NCUxnmAxDzQ5hsTNVn7gvC+WW4saWzMKF
kuj7FE1wJ1U7s+x3elKQ4HLb21VeOMazAIEH4gkH0iqeLN43X5RPtY5O87AC/nva
PQJgl1Ib0o1wgBq9AdNagHAUkfygId8cp0UL5ueI+iHN3SICguPxpAh1SKUOZkXc
U0YZwVx+cqvtoYi9Jl9NhWUrkN9rAZzgWU6oJ88VJJgfJyNEn6brsMoYj+a4EP/L
sb8lfSiRRQzNkeASk75JGQt02lCg9iHgNrLCZcFGAhPLsh5kN4hEHTcAsPGROzHL
RSeebT9Gfa+6WzA+v28BgJjaB/33805QkY32A5NvF6YpoZw6DqnBlIGC7l4gMP2V
BD1Uo9LvU8HDfZ1bYvu9S6HeaUTvjw4IFnuO4yvKbA9OAPdO54zEX7R8ZFO8LaEM
rtfYtC0H9rVCA8iJ0jtyXxGPpmBal3X6loOLhQMoK7nVxuILtiuHhRXbG85xQVro
t6byRpcx/qWO3sAJq8rP71cA24Jc2sap2Hk4HTBxDqnZPghpIjRezhAQlYEdSEWU
s1UHiUyunzNxo72ffB0oSR7GHuJ4Uo+dEKAPmKUY+zXC2CEJJd/UDLh8iOvnGEYe
IGWQoVpPiZ1TZqIr/K4+WFq1ZLEkRMcf0O/uSrHKKTWw27dvcEjTR0EohGyxeUid
Y2okl6aTB96u0U7O1s0k+DyvYD09VhVwG4x858eReCeS7xISx969INiJJRqorwLd
xZcgRJOg+P7FPI5zKV4NzKR+rl7Cot7VCKS30XU/shq3cNnT0ByJhzglfNAsdhPb
cMrKjsaZ1lCZhxPvgRvJj69cocTn4U1LyrZqp7nimTjdqTJnf7X19Ptk59AH25Sn
KcDc6Ix1yqsIVoDCsMMDTsz0aQ418C6CJDS7jgXIBk2suz4DgL4bdAotYZhsADzO
c1avWbK03PisLLuMi9kgrRNs6xU/rxbsGOvSwvYodCuH87cV7FfvhxRzFqsmMowg
N2DyELHOC/NRohFWGRbgqQQV3Iuqh6iQNtrtNNlFbi8NdjHhoNiYkBQJogqW2jc9
7f3e/mImZTusYPT8kFCVJR3ujacdtLAP6kv+WRGgzIYqVz4NGghxqzJFhBYipbtc
hLVpe9kaubl9Z3ka0DCFpnWGfsNDIY7jX5OO0wuFenerT+Wckj70ECsmgA0hlO7F
502y+kFXRllCylbh0MhXwzc+C3HMDCCZFUaXxuj8tsh7I5KQNrCmakQFQSzb7WDA
yLrxEozB6aIf8Eg6suOU3961A3zbMxvQG/BQfcOyJ8fOy4EO+2sO/d9ggBruO/dv
j01QU/Bn3OhHcv2RBDqddo6AF1jZ94l5B9DP56ZuABUjd17QrXI9MVA4vSjJ4Jht
4Y+0k4Fvqme36zwSS54Cw5TOJRN81+CfGHoQ2XI16hYHYL6nJjjsdohvyM5UMupY
+AXLPGBSQEBwQk4ixOpHdoBPNV/GwDjl3/EfWZL0g1MPat7YymFOxd7w+CiMvQtN
tM9GH+185ck/CUI/DIVizQqxqwhpRmG0vKjm3aV7nN6QrH13JLv76zFjIdYDXs+t
gWQ6xpfGSf4G2esLbHwjWnM8X4ZZkUNwZy5qm0iYBwXd3JKgMYhFPuwlNd+MKQ2m
MzMf7adfoUkP4OdeuDIJdRBeLikUp/JDAzbtzgWmPYFAdB7p1j0C27k1CkcARmof
ZvbYodRf0dJInZqJHMzOW7yCw3LwrTZJHusNuPLT67fUnPMMUkb9iQmvPbtQT1+8
fyHsaJhpzLB24krB8VWeMQO1msPdqFQL9YQaNvCViZG3EaKeHG0yUzqTPWPyBI7H
cez0Rb9WqYzz9rlU6r2UBEj39G1NnoYziRwsCezSJeWrpeHEM8TVoAJI4VihRxjv
qgFFQWO72JpoVHHfICh1y/17ZsA+Wjpl5OCC6+8ctKLWXMRO/GLxfv8QlI98MpnJ
HtTUtWyXPzXyv62v+vfK6tbUPMoSjallkXfrV6Riyodv2WHgfJD/ud/4vNuMw9hU
aIOqAkSjyGlJgwidgvxwMZT65G/59bQEirS64udeCrjL69ylluBcHBb73Mswo0Vm
nAQiDt93ZkvDulVrhxzUG0eucoCFZ5aqm48vxMOKGCfyzKaEZMeZCdyLO7SXUMpN
hW5KjaeiqUaCyN4pFP5gqG1r8JumQOUDb5TGYdUSTye7rAolnSPbWEMOnwFFLC0M
6zX4GTdRzNnp8lgNm1nnXpydyBXuahJq3fNTl84KmubXUxlr7iBWr+utN3e2NRua
b4RFG8P21YiGeMwC8lhZm5wz9hy2YEI9+IklvTe/g9o+F+lPp2WIhp3qZbWJF0U1
AqnWTY4tzk7uDPZmZgbLzLu4oMFn7fh+hhTu+Q+TcMIdnKeR5/ifgEsBQJYSUPJh
OpI2KpqiRQQ1N3Wz5zg6cHiDkl3eObbbt89JsVDvO9SXkaldwjPbWYy7U/rDmxZ0
AMX1udQwHkdbLIUtfFTqh9CDOmv95i+MZTHVS9d0OfJqclwCakaA16geaxjm02Hj
GRhRrmm0DGdWlN46+9JUSR+/F759uOI2sZ1n7z3JSE4aU/H2qiKz2LZIvqV7s8z8
rWwvpqdh0O/4nEMcpxIEm/7ZjPAjPvMMqQF3uCwoDNomCgZb5+vlcFDYZTtuOFiE
50oLS+F0rXh06D036WOgPtMV4aOidU/4Xwhg1YbmBNInHjPK/bzU/L94nmDqxYeS
oaCPm8bjwxxYbKG1gmwRHbmIoY0LaMzIT3tJmVVWldRDBWkmgrkc/MsIux0NFejF
rpNtIHuemPsAFObq2Ww4FnYW9MNebv2CFiWS13rTE3bSzxh4cv5yr5cL1C6f5yPp
YSe2042XhHNGkAoLa8rpF5XKm3mTW5UpQH5DRTohqzuvIbHMOM+F3E9HKbpSt3oK
eSx4k+pL+Lnhk+nRBIY9KKKACjmWwAOzOvYqOlDZBzWjWnx508ARL6Jv+2b+iYLe
h238JuTNxrvafJzlz5PN4k61PUxCJewvNy+5onTlTJ3Imb/HPIvtSr8DP6xAveQK
Vhsi/gtbBKtrCd8Nj3kwCQVUgIXx+5Bd78ZR/X+zQ86v6D3bldO8b+iPFqxkb4Wv
43ruAyJv9R3ep62kmKBbZx+K4HYfPQx5ZtM1Cxh8EfvkTaOqqhH2vSvQJ7n1C05e
RGOMd0BqMeLS6HSF3hG8UCqQjBQyCgd4fEVkp18LILIkJDR/oysYiDTFIJ3Qu0Od
Q88vMMiYsO/e7wqRzQ32HK7zLHsCKWi3uLRU7nlG2g2f1IJvBl+5Fn76F063sMIb
SjCkvZtlMpO6Y5efLA+PbgiXH5ErtjpvxtbnDxV3t3hYCxes2Pf25QXoC5thfdUs
H5yG24eRbWS7BJKJE7vkTWVtusyYFCWRgVDg1JQ27MDPRjpUVYHUemFGA/STseGM
XcW7mna+a01340xPGgSZVLu5A2s8d+zJ0ZKsIa8UuLLS6kzmhpVGyB0K4gSfPs9l
gQ5srAodAjPWRrJ1w9x7c2G2hnxwIoXEBJiHPb8aYz4AhjCtD54XdrAgEW73hlYq
Kqi/LNbe+JLLacIr2TrFKvtsFmie7V74Zn8jTc3LnGfaQdTIs+OJyR2L0j+YEU9T
EEW6EmzOvEXHcr7sGaO6Ms46vAQVET2k7sKI8KWJxTVHFw+KZw0QP9wKc4DmsL3R
S6vO9m9oe9Q3JbF+Bvk9SEEsQ3QlURW7b07f97bpFBam+/zBnlmJM9RkEHWWROUy
jL4znUXzJZBZNLRwCFBfL5nQFlz0mTHmxjW39xSnLIJ20eG2Unfzuxpe/CEbz7Tk
orz72fRYi3yoE9SP0DNEyj7xcormg7aiFK36uhpYXN56ZSJ77mKBQLka6s2Lxrpd
9zrTAlps85ruLFD9g92C3j/hM992JLwMIS9v22T8Em0SCuUea2WEF9FT66+0T7wV
Cz+NP1YcsE5ZSPIL+Y9SGeNnE4FR7k+97rWk835/TOqrVw2hhQrPSZtvHRqo2tXv
dyji6bmB+tJ2YzEePJ/CWugG0QWxBhSjNGwmU7vqrdWm0v0gE3NnugsaDsUOX77k
xGYp3SZj2UXeHDvL2mmgm9YmXXQytWyWtMFvo8rR7MNcW1l0wqK6UVYSyBNsfkNb
qk8f86HXaj3MRbCMVfCJPsUyJwUzGpZVK40jG/jBD+ap2i3+KqoBUctN691rVarn
cD19b7sANw5/x0MsYWQOWSnlYq+n3E7B+SxwmCZcFh1FUyx1xKBbfdvTH4dXxDFR
bl9JF6CwLy1XEZ+X/Rcvl9039Zbue0uRmuhQyMJqHVpKVfOG+Jm7b4TU7qdzzXuE
kd4T2Hui3NoDLZZoMLifeKFfFE6qhwLI8yNpcxry3iRlIT43MlMnlRviJ8xdOqEr
Zes6xt+lGxmGjjLOt5tr2SyR35dLpMmePN6Eswt+TqAhBi/kp5zwVR+8LBibuSdN
HzwYGNNuyriI57UOHaNkSF6smL0/ihXRQE1rsoJmPORMP6utb2WClKQGskpxFfxS
nBw7dPPn3j4BvSWWaRvmi6BFzLAJ+AOpnIQoZYAbKM5Dsv3vd+lNpoZLg8reCgh9
Qq2HuIL8ogOCFdB5Uv1Fg528bJ6AKfupJZ1koIRq/NVSj8B+hMPdwJvwWCOd7ZIT
5tvcoka08x/NWvhCMDxaiUxReWC2aoqlBFyN205CgVPdkABGBIjHeRrSRU4WumTR
9PX5iSBLQqSnZdU3KVqPDTMeiWVAa9ykL3OZPHMAoHk4cIInNtIoUdsPNvA+OxPG
184SP1wqXsOUnprSk2QfHwF6hzCiDkm4m/7B3fgqLAdpFq7b+pAzQ/09xkmGo8aH
exlaIXDxRnHUIqnWN04y2LrahixcCeAiAKfiIfHNlaZ8WHxHqUpCO0JWyJJAF/6X
zCKjWsfSvd9DSVk/qpQIz+K06FcRLdRfY6qjrUB7tatNtl7T1PAKFRzH9kKvJTvV
gDh5DYxboEoGldS0rD2HuC45UTPkLqPzuRQ1Ld+hTbcT4OAjtTJri8/heb+kdyp3
uavoT60xDTckncWCsfcCU4dlXBTXMp1Z8Xc6F32M5jLVIduLbcXlyioRKmRzae1j
6cq0NadW9TSbRuPudp3Z2dictIVyCXz5S+XOeb9tOH+1HNeKfhEDLp+XtGi/A0mT
vwmBr0hfL4Bu1b3xhcLrYTNeARXMzbxFwXJQi/63r19HiQIHVCvfVIym/qUE1By7
oJWxqQ+z2ZG4V6O99Sgvw0qjDuchYfantZfEs+kTlW4LVFsfrW8kFzAP94yQYcP6
NIR3hFHg8wTgGnQQMJl805iCpJ/exVajUNQodspFkaKK77ZiIc34wVpe6HqWsW2h
0IyRD+Zhc7YzHPyS1qMFFJpMo6T0jKJIacRF0yBNgckcM/hg5/aH/ZV932gIIXnR
X2zn8KpLTX+1s1S1ZZSsZA/lms9VzBf0rkGPx4s1FXgOANFZk4qL5W8lhBNg1DFp
0JPO/jRYYlJBI16njgI29dqHXNQ+nNRYGHNlW9zdvxIdBeTBQqeIQIJCratYJm8+
1/KY4DGToX+meVntqPh1lycinMXhR/qhhpkG2f/eNcvZlStJkTJ47u01juzqdpZv
V1eobgwM5fV4YCOiBEdOgF3yFeZEJol+riaAFcO3OLDaGlD7p1fOAUd7IRK8ba5Z
iIJasvHOuwqx8pCLH+bPPiBMuudEBPM1mVZcg6dN9Sbikj5zKMHSSEVuHqafHXvN
KI2oLjS2RiD0iQzG4CsR7yRbqHrdAKhGPyjzPjse/FM7pEQj2Y9GAKAsJQ0j655W
B+8ZXmYQwO7uMwNw4NFXLDZxN7Xsu07Z5mFKJGAQeIknTmYvKmChZlR/Ji9djmXC
FXbIs7YE8AfWqnq5gb/P7a8ebzOO48KqwNA0C3HVDf0i4DEA9xLWigM2KtVHROKi
pLiA2jskPT4+zQE6/RF8aR+BiTLGtt8ynWajUVsaTn7a0g2iN5ITAlusXTmlBMmU
mQR7sgc4DRJWX2MGqp515PEyv5hEy0yTq0d3jrK3dqriJcGthlaPf8zZ0aG4zZqX
APqwxB5etAUpCcyeCalnfmXw+mooguUSuSY1XGEuv5f0COyCUjkklRCJNEQMTFgp
sFu3xhZLr5WSg5gIPh+R9H3wFrOQ5yuapJplF3NgHLaq+TdcW6nNe9vY9NXU2/YO
yh0o1gB/brCK7LTSN77wIljZbXjrRTOKdGwzt13ISN6sNgRB0zvwigC4hBC4yA8v
3dysZz9EthDmQ6z2e6zZwmM52RY2OSca3KqLx7sytb49gLWZg/TDXvbmdxyjeMyi
Wr8EBfK4Y+HI77hvC5O/St8hWY+9+VXAKdeH7oWl5tY1qBMoPSh9DsJ0tE5CKddC
ppUMNoVuJJeuMkZOJuKunhNyD6L/XmrokvuJVif0ZD7Utj/Kr0xYyYbCxLpQtx+k
It0kb1Qee9Ve9QOjycvof1KzZCfMdipltmTGZyFO+8s1YZYcPaPmSpXYIVWzvKj2
jEpMhqOCZ8voNvjKjo4CtxJIHjLPMm0qFTzC4w3t8+Q0fqhPTKiJ0/LrcNRBjcNR
ueNeiAg5B8yJIMObPsy9JsAKLSpuIPx/sdlGCiE6GHALbhS4zhaSNBkKou6I2HE9
i/8QSt55I3mADOKntC70TvtcigbSZY/otoKkA46FEETpyPYjY8VK3+QX5/wIln4P
Hk69Dm2EvXmkMgZZDI1oTx6ylHlDY5Xy9q1CxCscpvc71ty17Tsi6WBDIwx7rG7O
BeeKBFFwUFE5+y54NpVc/38aBcGvNFiHcvjlCeSO4qv5b3Hha3ArB9nnOtro7xaT
Q0qss1bOTRddE6bEfhRvSjPZ9rGPxiWZec4lHEWCgslG/GFb0rHuqOJASwJ4E0Qe
b8t31EzNlDjnEXJm/jUIMMkckBqtHNcORJ9XEJGKflPbEfSgYuyitwY4ArQRouGh
Kv1xOVVSKmuGQa8duln1sCEJaESr0miLeh4Bkn4kYWLewdGgb1TI0ZuTvaQjCZaR
rJWCWZvQLspFoRx3t4DJNn4Kf0kpD8viAS178C4DwPENf96BE4O+SGEVXH15DdlP
dLP56n3GwBK6Q5uIOSa735HJDtBPz4y5sRgjlx0BRt5DSJ39Q6pb5+b8jpfJvyin
HnJJ1SOnLoYA27gimF9AJcKvBN7X+OYnJDlNEHfCRk+n+QWadyqyorKVn/G+2LtZ
MYA4wAkqpyTdsUPZA4VXp9xsACbddCFOnFsKF5WarP0Ob60px4O0CUzkU7KcMJ88
eO72lfBhY1Q2wsRtjOj+1SPQmiIQy7dZ60TLGA8IpNWObz19rMbYcl6eHjGmUh7d
znAIexUQhp1AaYNEkdrviPDQVPAJgZprzubwMVhoWEZ0CrYJn2VeZYsGS8w9As1u
Qv7rHBgYm81Zt4Suq4cs2SPFOjf2N5WDeLnnjkmPF5fbnH8gNJCaPOIL9gDlHotH
duGExLBnAN2ReuyWzneSHHSqIkjhPICo7017tuZ6J/9P7aKcnFiakBX1TXh6KuY7
AOb38goh4cGK5fT0wHI0cAn03SD2sLQGlFP2ia6HkP2yEnef997MMbaC7eHtVrYf
OJlVrTaY0lXS14ciIV2KR0ENB4vnnyFe7yvgdMvxFZ2jMh2EDMzDidfViLglQPmB
zFdOeVa8QiVp2xpt+hm1jb5z1NbQeFZZmimMQ0uw0ftHpingrd9ssyGHnbpS5zk8
8q3wKdC/vWLL0GJH5vfOLOWEJBWUG/lcG7oBVvEiFLugVug/cAWPrelqSSwqL2F7
ZDsJT9553iKSvU4KtuIUB6pSWpDd6sT7CfsBkNf9Ebb2Unh/SZVEi3o8iCp/pekz
hXpP4iNXelhCHTNSZys8QX3RXaRvRuAomDZUB0F16UVOhjeToA3SwjRHpHwayyqR
qRttc6EiF2d6dk0bwr+doDu+8KsCDJBHsnhfaqYh0wkCGYtDCg9kNx+2b7OZJN/j
TbS4xgsc5gukfHr+tDbM1Cl8u6+bhaonCVjan2yS3j/Q0nYiTTfr0xa2NS9JS1Cx
rFfw66Sy/ZBNYJnBNYMrPW+YFyoL4gbO+/T/B1Je5rFuJMfGH2Y6USyYMuwOTgJS
+sUGDmZqQbKATAEcpwkAo2jiW5SZNTMgj/3U0th9IUxnuE5LLHT+6UDq30mOZXl0
WhFgmRedDo4zvb3L5aszVO3Cp4kMBy9rTwwCHM40kzwxngaCAle3OfwsXGxWlOnd
KLoufRoXG2W5Qy/9NR4pKq4y7SuaItYdbhk4lKGYUcOEpgv3lCdO7FEvsPh0J1t4
NDBujJZJmMbJ+TZTAOV0M5P0tQFdqnhhOm7z8vcgWbs7Zh9K93wFQNlfFzMyE4x/
z2k1nwn+PtpFIYmupKPH8b+9o2oBkftl2dnpG+q/tOIQwJtXUf0Rs1bnFCyC9BF3
3Prvm2PCX7kohEWsOamgnNXAIAikXjMKTNPR0Wl7duXanZR/vc15KoHw2vjc2Yma
bu7UyIAszOfw5MFgzh8oOGK3k+/IGnf0nV9r7tBGl4HOk0epSAzqstwDA/7xh7K6
8lNZrS1xG7sxp5AJWnT5b1ed6TT4LoZQTE07JToq1V9qKVgqEJEGCylM8Qrfnilj
LPbR+5WpzUY+hhpv/OPxJ5u+q7d0CEyX9Gjisp5JhyVkOXaiqxHQECOkQ1hyWlCY
dQE8WDb/DqmweoK7z2YqIWOagi8sv7qIONvfVGO4bjhaSIl9p/S6QhD3tG1XmWPL
IOh+k/zt8buEeoT56UEY5ZwdO5koVPRs0/dL1XJ4VVx/pAiJt6kyV0k+9JlOw3Qs
IhNbqQH4F5ICXzqNbU68f5NMA0ZxxvCEKTKObSlCkUxb6TcEYN4zO7IWHZbh2meZ
ygWuP1yerXAJvhvmlXnJx9vBl/HZsKf53z3PGCZLp5eHd7Z2C41iqKtVf/NR5yMF
NXwKgbMrSCjJP7Zx+DcJ7I1/Fu1aYY9J+1TXWpS/0BWJgDDHGVpml3yoblndGNld
m+SdpvSvkla0GaLa3S2rcaxwnzFBiEZqBnAXC7t/DzMaMe6o7hMMr8cKB1af47y2
npzb9DMMrpWRfN1HFzfMz+zJ3wEU4iXZyKAyCj2eFYjsmCCMQANMKpvU5VXVLGwl
k+xwDkUkxsSxdlIH2URQRcyVxMTTcp5TgmWhZ0AZ7qXdNg/M4AyoG7ocfJAXCRbM
DvdC3wsxfT9P8zi+f5zXdgcoRduf2u54h+paNPxGgn686HxqxnyiRBXx1wW8UNKN
eGVRrmk8MLlSDtdomwgYJO5Ct5K1UCLRc5I2E9cPbeNiEce5+LUYuTCd5pmzMTEW
WHBcE41UaXrIj77v6LjeHCGNdFcN53KpTmPS80DdCwK6OvYuyG7VD02T/su6M0RC
Qz+O2RCPVSWTLv2g0okizpXTYUAumc0ra9eiGPWaBSRXDyuVSc6rdAh+4WGqncqc
BT6+C/37+SgyfzcA+whQ0uIzlJoHdFoiqB8V0Er36+dFUdo9Tlx/QXIgd/K6Wdx2
XKju1GfBdqz0hQ5vwFSCZi1P9dA9M0AtbL+MJaHzKSCRqkGc8qXnkpP8JFbwL6NJ
PRGzWbtunMQ083RRwDTrsrpJs7OonJJtDKi5c6jrgrupEZCTQNrJpPqVLrppqzv1
SDxrlHag9JkfJcukJfTYwIMnpAuBcsOx8hi9waEafROwSUtZ5t04FgejrVpqhM52
tr8sWxpyyAZ6CJfE0ugGhpuXCxVfUI/c7o/w46OREU6BnMAGnHNPkX6c3tHg3mIX
Rob8bfykPj4fXnEqgmC6oJKwGnkfivqVnvRbmCY2VBpUNc+8mmzf7aBZraj3HJQV
r6uZb2ns62f2bqidNABuAcqVa+ITTIBLSU1eQSTnMhmrEhOBUgiYdOzt6QfI2nRb
BcAbe4ZKJSVQ9rAJxmnLp6QOhyoEnp+5JKvr8NVSvVXxmT+QOJlgtAo5q7MED4fJ
hfdAVEv2J30Oai0K9Af1Jb2LL/VeJgvv/ZSxRCsiUTa8STKMacUnoGx5uZViPj8H
xy0ZKhQWQqlq4RKnOFKRRqizVIVLzQj2tKPkDdVvn+lvdYS1WFW63AruRPMk0FZp
/DxEddKM6e4lzCBOoaf6mkRABCgyA1JaAN/ODtB+Q4mLFnnPoZaduJMryqL4J1J3
+bwEneBPSvbVvXD3q27jhdDXEP/NGIF56eemEFIleb30qdt1oqD3C9Rl02cTqR+F
ESgEbYyvwgkcedOXrwWiyhL+t2RyxMAnAF5IMRFAaECO2EOqmJG0nfg6ZhIYgiyq
vvZM+vivLw5Ii9r8lrtfDPWbNoPsmZ0Kj7cwZQ2hJKfCrou5JVGCL3JSCDc96J/O
EHVXGA4VQqowa+ZngzJ7iif7NLcZvSm0KUo6Ey7f1peGfOPZYKOIV3MGIIV13a5u
RerUzu8oqh+9Vz2GNjGQMhkEiCQ7upJStHp5FqlYMTSmVu/BdnIdV1gAFOlDaucN
DzqApTX9qmvWudAX+yeB+8s77n3dpbrFp4vKJ3PVxLkjpcgy0Ebry6XXhPNogPrt
8G1ltau9T2HvDwtFx+DOEatzzx+GkeySfn+WNfNWB2YSYDd8dsalTlGF90Zt45QB
UBco/AUavy073fShj9R3Oqq3Mj+vjsr0wl4Em8fy2OuYUilwaMW3QVf3tyPtiK8a
UDHR9j/+pZR0BxnaXa0hY/HRr8VnQF0zmT391lmcjFHSKIh0SH0bNvyhbza1+P2Q
1GU2gMQKpeBy3CUBy8cFygbmDKDQC5PWimJN0l2RGd7tv6j0s9KxAEVS03gS6w5r
NCgSLsFJdWX5mnYD6eZyrYjuBvFGMHNMoAFwPlzxOblIPAsnBqdsZy81oHM+glwI
S5BxeGLcWj3y1IaUE7d5w6HcUREE5NsIY42565gT3g/eXzkjM58gW0WmEKnfVHB2
fz9lKuJxcstrt/nvsIOQPNAX380W64iAypVsz+i4l5OEgsOxkyDJo4cjwKALburR
DInB1UWQ9RZ1a8yPj/l7TQu748meFHsc5tUMtyQzU1r5IrHuw5mdIZbhDU6EYsrC
uTkzay757+xIQfdgEUZ99xEdO3sB/aulIoas1hw+DmAjXWsraYDuJdObCB22qD+o
Rw/cxn37HNJpoFfvaI/QCfLTFZfTEUx+D04SepOVMoPA3MIvOY3VJPYjhh3Y4Sbt
qmfeBj1bwKgAm/0tOihG/TrBcSdksoItNXMtGiH8kgYjxfYpKCaM/0a/RVbD8JXX
MBqgAO1Hbz26wMGjhPQcuZkjy+c1NPRylEpw99LZIUt9u98ElLs5OPkkU1uLsDsy
NQ2o21W51gs7a3SctVNQVDYlS2SnVEfQFC+Ze11/zwNxrI02y7aFr1TSIHsAYNFq
MLC2hTr9GnF1Yqod1xwLJ956V63+J7SDhlU9j+/rodgzjqjtuQRoToUjyS23jV45
/sLPJoNFzCL4Dwgm1Y/YIMw2muY5zll4bWrYWHZOrp1VfKb5VlxlWFKhWxOX4ijx
5jNDx9ZGwk4YZSqjmd/EAyG5nhdlPLdRihdYaIKbu9g1J1NjIzbB5CRRxRlA+38i
1SltXd2gWoKZTEIXqxEQOntsqEGBjxjpnU7AcwFxtDu7xaxi435BD8vpTl+SNA4+
pzHDzyne4/2bFor5jXtUuQKbcZ/z+80NfAjp7VTaEWSxcliE2KHaRQ+3p3X+GySy
XnpQ4vshkvaKLb+40FgUbojJbwXGYTYaOvbs0LNvhQhdw2UMGRMiIlh/Xh+KJYCT
a5ZWxBZsTjqmm9Dy5NncMlWeVcwYZfKxqD8U0tJw6HEIlOxn6lCIS/MKcCr1qgXN
snU0G78WPW39Ot5onEAd1CmXugNme8OD9WHxTXHVU8V4uhvux8DzdIbXVBGXEJZP
FTXQ5dc89Np6kpCztsNXKE/PHwm+/kKdXrTRlrWkFzzTiF5xlG7e+np4Fl0Qig3c
hDEC5aGO4HgF/M9qAUDH3s+tz/0n79wJIVDVKFyGDA1VOmPpgNIg83EgytGPun8T
CluDNZ9i8Ey0bh2uqNdMUoOgxT+HFFbH/oAFZfCdnCDn4Ua13hExjMSAX66JaR5K
n6VQ4qr7AkdRdrT7jTxYuYjodDWhR+64RknBMF6YdYsEOGdEIPakgm0h9gmOjdGa
NDAk7le7MynY7qHIkJDlQ7Q1EKMH5ni+OIwfbeWYZpHO3WOVykPuPEk3Fksp2kQT
xTMbwgcd7VybF9FuDS+OPbHQdtlu9U+QyiovBY8angc0oCZ2BRx110Ld+X43j7Oc
ddMhiMtJs1P2ojCtxGtjA+joUndk3lAMFTSairUqPcurFqbvOc7BpsGhzcx4TL/W
k0IwlQgOl+rGlkJmGvmpW5gP/GAOSWF/ngC7Rf0n84/JLQil5JrRw94ewCl8Giea
67gTbQK6LuobZG75s7oNkX74/kew3a/gd5/g0LbmzFkT18hr7j8aOgfatSoHKNVq
8kFTWr1krMWBeuH+5uG834dM4XzB8rn4uzH0TOhCd7uzuaK58ox2s2wJbarBZiqu
h7Z03LXrtOS8L/O7xHJWd6dyyAszg36yicgRN0T+UBGxPWqslhXEERj/aESJDDy4
8IjjlaxI6xKfJt6Ju5lePFwc447yiXn/hXGu2oV4SlOcPZLodl1ON1wWoFoFTRfk
Z15j18zx0t7V9dk76DFy2rCQOsDl6Zf7y4bo00QbK4gTRwHipMVpcfayqWsq8OHe
a8IloWHEzkMWStPZ6E81LnSRGht3bpwIlaMT+DpKMLQkSe2Zkv6hmYAcBoe1dBRL
ZmTQYMtoi09S+Bs+8+u0PYzFoT2gWBaMITMgND7n14TGrpxI6CD6BeY/B5rB49x5
bB4nwS3UMqayhu1S130dxwhntdZp+Ekf3eHMkeDcWxZ03IC+WOY9Pz/UOKo/TBby
QLVMcnbu5l6dHv1VPZsjK2ccdHBhq9ZegqVUsmIX2DsagsPOLyQm880B5LSO3bHR
5Zt9cCxBjROryESVdaXX7HqKV4aRdUiC4Oq56w/mALBeyroPPNnuN2lMOUdtsbUu
GzWOtuUBQHZJNP8lkSoadj5Ez3lF3s6ddcpgCF9n9atWAGRGbchNRE73aPRCG9IJ
IJZZXUV57i8NFXpMG5wguytOp3EtcWuvJQO9WtzpOf7OkNq8lH7kabJoQb9hvKCP
EgkMgykUJzzu88++hBfv2OVbq+6dH5QkjA2KPQ3CUu6iq6n5IignMqpc2qtomLKe
eyPnGM6OTTJzNkHpMk6/nqBHT+Ma+kYaYoc6HC6StJDwUSF9SlcX+/GecpO4s10Y
2zzC/lLKfocucxFONgTSHo9vfMivBrHY/mLybMg4kl55hnhXH1FiV9n32u39a9KD
Eg8iUBVLsJgsTac4hHAzuhpTtPhCWlkGLinI1OLwF+R91MtYhEQUfD7hoD2z3cvD
c85DH1+4qwYinmnQoMwRlHyXp8//SrlvqWQDebDBtEA9A045Kxfn8u4HMPFnMIAS
heZwxcEpDM9qKUj5F8AYcO3S70x/x+gKtKAAmuzODXu8bHH004JffzjSMEMYBeVy
xdlfYtlx0KcgnRyXEpR01IiwmRpatKP8XEZMmP60gurUifEOEdrJ+xpqPgendIpx
reBI85WY7ayM8hiPXYwGatecUm+uSQscZ2fbuXiqRTKZ5u4Yh4Hb7h+5Zk6O4ffq
m767cCEDp+6dT13ivH7E1/i8cC2VghCyOyIFpEI8AvZSTBA/SHoiwPuwLaaSjvAK
Cy9ZKaI2SZ8O67RZyCW7erpPHGPzcgfhShxfkR/x5LW9ECaiCKNycydbDtYR0VXi
c74veteybZHjXF+NBRLLaeGujsPMod3uqgGFANabmjFcZb++h0hWgzk04rh2CsVH
Ohq1am95E7ubVuczXInxCFMxZVPPF7fCBxCvscRj2AGX8lM7qu9tbYAUnH6wLDK2
785vp0m54Qh7dTq8R13yV+hXaox5IZ1OJfGYiGHf7A0FrRWIIrkEIXTeg3RZf5iU
d3tD0Hk065Dw1T3qT2rA7bowlLHcOSkItQztqJdf66GZWJtgqyWeP6aD8GMNd7Ri
dUVhBOu5dZqTCsJntymgiQbEfrVfUYoAMO15r41QO8gU6lwJ975C0tcV0tkYRgbp
Hz9WVILQ/Y3g4ecxU9WabFY1zyg4eoniDzRU/lOf4n/NPfNSc70m+ipZzOaeOW9G
zI7qdmK+uOmvUSa0WppSW9k4HlBB1/6bdyy5srosRAxTT0vhmXJFbh5M2tL2B4cs
+9obysNfDWJjC0Jgm+7cPzv7s4uypK4z8InOSFu8ZRyV513et+SB1gA5iLDrU4lN
Hkj4/G8hya/1T0YGIJcQ4GQFvfskds/vTpIljeGoot6k41Wcc+kT4HB8pfQT/Tl3
f7vsyRJ3k4PRs9GJKoMZL0iB5CAwXwywqSVR6BOd/YaRZWyvLgt3EavesRyAg/PJ
3e+cZApVeUhi0C/JvA4sjvEqprdyU+Wq2fEHLQs7sLZIaSynNeN0ZetRmfbdcQk7
9aW8BsIRJE1ZjVCzGvhl2nP7YOyFVAoLLaMavLRUwy1Iy7ETbbavDMCHOHA2aDqW
IWSTG+rCnBAQfKq6Z601TAZk7TcPL6yPLeUWXZ09GJqc4ekkGZh5YU4g3XoVWqPT
Vyrx0jv0TNhyswr+3+U8gYp6pFhlCzmSkhKi7pDSHfD7aSkLJ57YzD50cmdnSKif
i0i2BqThyFA18UkkPU/7TReGpSV/j0A28gjvv6kt3X0XkO0W05mY1LJVdGZUwz73
M0xmlPwF7ADryyStV2DX6iN2PDVsgHS+Iix4JAt5rL3Wf5+Dg9N7HjMlDv56jJal
RWnSoVY86Q6U7IR3OvPLQ8V1S2MOhah1PWwXUVFhICqiEcZAZFzF+PHkabGbKJHl
pmQB5buebhaRqlnBuQGSjT8FgRvkuBnC0bkXYMQkEcl3YXejy2pq66KRXsZodtVU
gvvn8JvVqdAwPOWQpNfZuo4KoM7kAfsCUbtaAa9bgb/Jf11dUZnX6vFAheAPV4Ab
CTgsIoR4bbgLh0FPQ9t1eQkdbNZWUwSzbY2aOUZPC8O+6DSZf7f8EFL/pLlT9QBF
LDMtfEjMjuOKgKNePaPt4aT8UGamOB9X31M9h0gWFhcN6z9AdokYlhh5ZHCW8JV2
04wfKpcOTXKKZo+CtU1iT4L3AWcZlAxz6RI8/MnCtQzRrmD/+nvS/3AwJn1n917e
7JaddMXMHgQQyQQhgE80JSi4hg+s6EwhZihlOXe0vC4LhnKmpTTsgkzaxMJkfhZS
TkRVbI9QV/SavOWuOfwjr1ajZyXG8/+ofYITPUJ22N6WZtbQ+UMYAgVSWjwEVmMF
jZOSghyo3ez7FSMZOWfa27Se1cDltvs6ucCmwX/AiDizHqJNCKt2b1Uy3yvdE5h9
72HGYpaBrXGd6ikRH0zLEHoyoSHINbHe3VXWT3O9gvVQdUGQBQaAw2T5BtCX4nn0
6aUVpHTNS4tJD0RQo1ZCjX0Kc/PdfA4vAT1T1qoO7t86f5ZG9EYVEISwdQOjKspE
s4ZWL2Y8hTinPVnROlStjk9xwHPjAbLCheSfLcwEPOoFU4yy086UTdOcnqs9CM9G
TNF3hc38Ifg37lSso/109TWbSWbrwY1zZp2N/aulthtupN1mGZa8Kk4m6wIUDu3V
ljZQ3x3RL+TfHVEzPfvZNjvAAO4ZWCnKp+nyrx96pbeqfk45BnOAR56T0HYik717
wUiAz1ZehWfj31O5XnyowtQdx1ecOYav0rK6trcdmZY8RL8UQmHm+PsNre8YfN+q
H3SNbCm/sY27IFVKFqOg7LSL3fhiKCMzbtKadt9i9ZgGMzRu9z7pGlctdyJfkHBl
n+B5tvpqoZCCkjvZzuG0mtYp0Xea4vXAs0tm7lfJoac9LIVq1U4ic8JyPAZe7Rjf
gN8EpKQO8A2QPyZ5Mn/sSuBsU5qfzwDuiSwynR0eOLgAM6HI0NzTpLCBs2NQhA1+
yoElyGDt9PwYwzdxSWrROu4npqvqi0iNpJWWaA3fx5fdyIUQFjHaHEJkOKoS7InR
CJshOzprDqqcTfG4EjFfasdfVIgcQqpPWz+2UEgkua0Cue4XA0SyGmCV8H5JiIg8
6BOKV3T2f4Y+93TR81FlranAyySfruZBbBP7Zelv7/FlTwXJFzujgn3brkmLot1q
Cuo3drasK7bU2F8XM+jUD5rGFY7rBGWYyZ5XlkFaJb/eMlXM3sRhi7M0tWzuXIXe
0yxKHSFPiFwAF63r7nHOPg2PQK7w+Joo/1JQcTmVi/VI3Lbqcy90evjK85dFus6+
71v/x+RAP5ebWYz0uuUihoJY6FM2ZuZKKEtGe1vgnMvoJhFp6SRlNZVkK+JxIcBo
RTK072u+LJB8J41TkPgg/nd5BHBaa93VgEFpk83aKsE91XkjJcLhz1aN5bT0qo7+
KfCyrLwmYhLmeQsn/8UDn9LtuG71VTrlmucdaQXIm+RAfWRyveTRW8uV6r1vswP/
/CsDftEKpKSlpfe9qS+6b1g2fCRg+jcKQo6w1xdUXgSZWU8jR8VXcClRgiwcPtT1
ug0j2iZ7mYaJJidOBMaCnxwfsfEx8OTqQVr5/kUnsk7Q2AmDX5MQXDTzvCOdLIWh
e2f35L6pcWNxHnHo6iJjDk8ids6jeYJcKgjyGcsFPBmoMYfuv727govSOyc3W7zp
yPtZZVCHsP1r5U6LSyHKRU8dsmem71xIQ+4Hhj7jlletwrqAO2w2vQYpYNjxU4Fs
fizgt08p7d4YFp3wA+4RpgPO4VtG4hfL7TfegfCWrHw+BTQ0a7Z3XhwoN73U4up2
uPVON3RcxV7KG2A/IOYTsj5FjvaFbnsXPl4AL6XAFUpf6N/gYr0e16iWClIP4qrc
bwZ2kLmKatjJwSbXLIQo9B2Aq+v+srX7qeLO+CDmnOurBSivQg3hpy+prH/+1FTA
CeSzHDjEUbScYTD/Zh5Lsw2/pOEalKp7acl6BCwujRRvhk+J1pTSNEXL+e38Hz22
v0LRidZi3Zq6kzrYKzjeLPYOwVX+gls2FlPzLB+DUkXXmIFffAYFnsxsLUK0Hp+W
IZN/IOSgRSM1hfsWj8fn6oLW00wkySAVJfh1/2I60w+L0bdHXX1FWBSFe35MBa8Z
69v3AxlgVWcRP3Wp9k3xf3LCOV7zYQojjqpro9y6Ve3HYE8GjN5wpEFcWZLk6ZT0
GI58Q6yrez+vACwfkyaSXF+gxylFx5rC9JcEZiaMJZHAF0vePOV7+hzmW6SXCGUx
4kDwp1Gp2OctQiF8gKB0hoJ95l9LntMpAIOFXdodNm8EUkYL5z0fkHP0zofAQ/uF
nqw77gurGiYunoBMh7bSrXsVzZeo3K2WxbfQvMorAypvA4vOTF7+4L6lD2CYdXLD
+Q3t3i9iVWwfURy5YwwKMSRJByOKzkhhEfY2IZdbtW4WflJ2ZgBYijw3qhx/GHiY
bl6O0iFYUBcnqxn2leDYctJMM1MMPJh7hN3FrEDVlov1B7ImuGppdYRL6qxX6AlR
WzbY66Q0tXCF50T8eP5Jk0pfS6zf26FD8KGMLGPGVRlKdsjiP6WKvOJDyMdf32N7
6P5h6glRY9k98mYfRfGj6SDJiWF4KWUTbm1D3GSETPlNJeZ3OMgRaPew9T9egZBx
/ZhDO20yggGy2V3sAy5pxgDy8dDIWRVifp4gcNSiFKQLyV2+4iv6Rl9qiA3b49gK
FIGlFRAstx9SigfxwItEEAY+mqR/jp2B4uf13KxdAPFhWtd2VO0azIcZzTzHSX98
By4tTrFd6ac6/lPCbkTqdSlEpyL7OmtZqPOSaR89VQwvvfuJCqFYsxsHEW9H3FFk
Jx4yhJsxA+vLGfTEPdeZIu6ThCfm/xWWHMsbtEnFI5tghUmL91DncDOp/qy5VriZ
zm/f6Krds6e2H306Fm3dFLVe/GqVqtjFQwPoEBuQ3jtT5jDIMaNbcFjb0cUbdqHb
nLH+0lQ+oEcGCL1vuIhwThcBWj7RbZh9BEkIoPN6Rup6fBl34PGl7KwpIJAn6vFh
l4ylc1OJOLgYnittMGn1kdcIog5+nh+2e3pn8BkREpMPNFDbzwnAHkNRNF3o6DA0
xzTko55HlgucSq0kY0zUioFbAe/F7ZyrI7vmG+zlRppkK/HOBMJVQyrsDUsW12TD
DU+fPp/I/AZaB8ns9JRMWHY5bqfNBQccI+vxKVXTZ8c/vh6KTA2oyLMBafvP9DI1
emU72v6ecgXlRvleiva+zFEO06No7RtB7XVy6aLfeOb7JdN+BJYPX21oQqb3n0wR
R4Ps+ReFvfW1lnkjviiGwMc7I9KX7+5lbWNWAnqr4icZ1wIeAzqMsHpieRzHon56
REGON0G90/HGQJVTeje+lCXxltfIbKSwtAGGTxtGTccqOul5lxFNKjue/qiuzLxB
4becRWx7GIxhUUOEJZr9oMRZgEJHgZMXB1Eiuq74Lc12u5Xay9roOGyDgC87fuW8
IqoyBB/O3vw6Lp2umiEq63MW2Tel0Q9tfaNQp0p9QvBwDSFNef5HA0nR9OoIClGz
MzsMHSi3HvCvM1fUqyVe5ZzYxJ+0oRmaLNzuiOLsrmLpAz3X41X80adCB5yJJMad
2dgHJuZr1Fg9C9uRv546rUmKYHx8BoAchCbd5R7BCu3AmWErtousIEGFaWlNRbOJ
yY95lY7dBqjjumF1BQFttMJXs/rQrApjckJ72Y5qPURKBDeQ2BYxDGpjkJGRUvNr
Ym+MUtAcjn40Ni5E7u52+LGYBkT9NEF4Q1LXaVDypP6U0LIIiY4tYwhAg07U4yzH
JQ+TC9v3A91Srmp3GMEhn5aXDIGIVPB/iTc8h5J7H5PDiX1V95oJEzslX9I4WzIA
Yvi4ni08vkF+HUxivS6RCsPQ66nJpOt9bfp9JLWlK126srqmxYk/W2Bo6S2B7jwP
RjKOWQiSeydLspfymPQBtdOKbhWOCa7pZfeGkUZYTcOgtQ718EEzsq+rs1Xv8h18
TQ4gF5+knnHK521YyjsYar1IOtG2EiDMnJuqdDm1G5+xUz8B+6rlB5KN/iQ++Aon
5EB+QD2vtJrIIflbA+1WCTjiqeTuCob6hLS6zMYATsoIdFo4mDvn5LvODAOPpNy8
eXwCplq1lG7YwSUIGc/s6d+qJebMNx784yDLwN3oaKO6i9gux1g4ijyXxiGZMwKn
SrKeDvUjGvLtLOPlJBPff3RI+y3hRa6dFd3I0sKSCbjiSLR4zCETxqaTcffnDQZD
8WiD7MAA4pXNQHA7DikahcpNdb+IAHy3roMRTRg9LpkkZ7PZiSR2YrqRaKMxy6XI
TG1AeD8toK67PKLqNNgERGInL50hwkUN9wS9Vxzr48cDNyS/emz6thmjzKkAUz+N
P+ZulyCJg8u0lULRoizUcRGPNoHocb417bv2YMQD/R7bAF64GofL/L2Tb0vvMw2L
/1iGQDznWX5ayIzU/xZNC9YNFR9jSfmup8ijyL6Lra8E4s7ytydCpdDczeGSQr4X
nSjdOrsvoBHQ/CoVVdHkk7ewl2DBjC9MNj7bpkSmWKC/fy/asXlwK8EixN47Cflo
QU/4FtHH8UO5D0rQIp6ty8QP4CWCfqjfZv3DJyHb9qy1zDJz6nHgj8Fo7veZtU6Q
3nIJHUtisFHl66M+iShwWVfrlc9VRTVDDqGtbH057n+sHOgpAYbGvkWqnHX8Hvo4
nLNNTdwAYv8Fn4jWwxy55c11C3SImjTHvSi5cazDUKZdh8hPginDZCO8Tw+VleGi
2ZFNFWePdokywWrvIdpAR36nIbXrOm7kD9S829NTfULSWiaZmgDHEBtG9hPnASb9
8Pc9BlXZjiHcCwShWl1wpZXSESWpIS1yzCqwCtK+PolBCBCtkiLJmPl+7NRtCXAa
GWlORsSusHSSKxRF/fAJxwbs/XIAZ8oX396Vn9Gm2aPgoZC9dM2RAKLcFpLZLrvd
mEnk1N58jOa60vzDRtwxvYWlI7T9BrXos3fHl+FwXhHXkjTA2wL4A1w6pKvx4eLN
Dv4A6XYyiWhLRMy5t7WlwPayUxyJOt1nt0ad9+/phWDBPOGErzA+zXGPZAGc2gCI
bh+BfDmUd2W1k8DiTGgtWhu/Qa0QMwftRRhRv6nUizYwuuHBL8br+dSSiHPGvTrE
gF/VqY25qubL1MMtMSrSOs/cpBo6u66dPJxEQym2xODgvSxI/GfgawQYftAplb3o
hBkDEpxD9mxBXFRwMCxcA5We7SnMxP9r5eM4Pcuj33cd4vZTnJcd8mld++G32xiF
C1MoJGlswnftHyuYC2+IWOLOYycQVE8IdPabpqteyGdYEuW88jM2iRJ6zUfwXd/z
By7VjlwEp/qhMJQbs2hJFVuyO9lb+Pl+snwRCLPlboKohKFR2MZ5cpsnMLl435YO
0mwLRUoU42PXQG6FGDzXBfo+Rt5WNlgpyd5w08N9q7g3m9aRz+xFAsewktbI7S/o
aSYhATDRmJxEalRASBcnHwimaWu7j+TLFwUqZ+be7rsupHpOK+PoIL1TiQi5NS6V
IT/bct1EGM9FZIwRtrGz9tvd9VkMlzSObnq6La2X6LtA0x3Iw0iFy+d02ZtZbP9S
jelutiE9v2Fe5Oz9TTd7P2CJhrAbQ79bRm0Nisibih3BSMkksSQe/PTmXs1Bpuw9
Eo3ZmAPtgFOgkiqP3rjOp3KHWx7QJ+0OEbW9RvQNAV3G21SuWuzQZP5CqfCMxgwP
IAjF12EMa4GMY+/xQvoubDvnOQc//7vwf4AGcmnlD0/ca/qTzlK/X2U0dt4TFSkR
g5PUT9adFTfW8AHGa+PAyWFEGGqJ/uEX4Fa4Dqi7IcKZBOZZ2Ap/vzbfp39qg0bc
GUK1DO9oDVIg2RMGDTUV9Gl2JPw8b1KvQgNv+OrqlssrFrKeSOqe7vTB72rrqy7b
qgWWrsNEIXsGHSe8InhD/crmZJZCWYzUwznWZGkmZnQG3Tkcd83jKsJr23MgclIn
priGc2a4vWQWdLylm+EkZRjkgrAlQUE05UyRmT4hHnRhq8GSkvbJwta89Qoy4goC
ksH5f4RDLYZZIwoQ+OU3krO7G10zA4smK/wR8Lfp0mXART49S08xmPyJTBKTpubS
s+/jJA96auCNwO2i0LcPW8+nMMpcig1xyfBEa8BgzW8lo4wqe0Tx8zeUEi/r3lot
mjmfzNV/6K5WUsj5TnnaUHUClHiAoFWZEWcPKz8nVpTyUjNQzcP4gCrpaebOJoWu
VRWtki5V3FxxM/CwPcIBlt6JAShwRBr1SFsBAkWn4fGJ0FVrt/ohcAF5ezcmsppT
ykua1Og5vjtUQ9UeOy9o/fcOoz9C45EgblVBaDWzR5rysVdQNuv6Pts/6/hbt/hV
Oay7XPxippAehsr73jqCSptzSgwTxwyUMeVaNhvrAXcYhxlyCh939fHrR2PPVBV7
5N7txol5XxFiafbxGk5iUBFHJfFHtYwAdgOVCxIm9JrMei7CtuygySIoVrm4cGJx
wF57mlQAgScez21sanVMKegXAKgt48IfpKQG6Vu9BuTYo0u+5ZUftmffTfYe5J/x
oeUQCHXwJW0qCWMc6Q/sW4v2KdE6Zbd8TTtQ7cf3fRCB5DCkkkkW7Yiuo6DN9PYQ
pF43MdhGyXzPwrFIvPoXC53k5wIjwejTgO1xKXrqOaFYsjxWtSS390AqlIMDkD6p
lftO02v8vRm95+e6KgvoS/8ZxJ2WEs56FriGP6Ev6NE7X2Zn8nd7P7l+/e53F2+z
veUTBuPud6YWGbvmZnVyKrpdlaHI1BAlxxhHgD1SZyyBlO4aXen+9sUGkcD6V9Kl
60OSYXWdheCEMzjXNBNdx2iRqSbfMlyu7adBAEVKyJR7kW95+eJE5PPoukf9HsjR
u7uJ+0nf6sLKClauJljJW3EHh3z8wy2R+AiGwUiPUlBD0bS2JKB/Qbs7qRP5lleQ
6PAzpgwG0HgqqBGipcT5NaQ5Mv2iqo2fqnrOygZOa1fADqFVEIccJYfK+1kI/SGm
leFYG9Rbz+FTo4N+GEwRK6XR9h8/c3jYGy/va/C1piE8nKt+tMDW9+2P+sx4rotE
Rmw4xr8mNk1f3b9q+wnHw4jR/eWhxx290dgQFmBNhPnTLU9D2Apqt7K7jsBHI12z
7GIJ/fjA5zgzTVWM0TZahU25UUtOPZTXdnK+wf1Wgnwec+eTAF8u1Y2LnCZr+nFE
IKRXy/yt4jbLuLJIm797dmlP3b9EdKWHs8ABUwq1wk7M5mG5wSryMw41ak6wPLHi
SSwh5xfuIvef9htHahakle+pB39DlOD1VlZURfGYzfpWvkpPGKcHJ7sMhlSJIYAF
DceKPt2/k2/C0THQPZ45KyEHX5EC208sNz4PO0U7vNjpsX1OKH8GOpxbZsz/yWjg
voNcosSEepXTU30cpBpLYoHe/i4LP1OPiRrtZubC8VrKtpq1hOmCSCxP89UJE3/j
ZsVgClOGkK9Msb/2i9p1d8zhAaOcJnkVb6ETrfWVGVvj76ANmjOwo/bOe5SPv3i5
au/R9TYgsA9BAbGkzjN5JM4+Qg8vw2smsD9kmKhb+2EjiqcRYU4QJA0fughjULp1
PyXaXnVy7UvhODIq8as5Tie51D/BiorbSGI1BnHtsQndVhBNmkpFoMbpmb2hmVZZ
8vAXzu7bpO2nt9knIIBkS/o6UJCTDTVXSyur5AO/Xykvugez4zGC8Xth39Az2HE+
jVZPeNQERPE5Bm/XjT8ajjrNVV9krInoZvmIROZtFVoKQVsXtxZw+JZ7b9IetIGQ
3Sc4eGtqEwcXM6mA+1MGfZaxoDuNBdoZTejKob5bh4yNHR4wbQG6Fk7CTCHpSbPh
tAUG9Eu4Pp0ygJ9JYSPwIdGkEAoBiFQdMdDJ+YxXp9O+epA9AiJ9+2MQU2yYX7ge
3+C90sOU2fkWRJPaoiRIEBJ2rD8NJv+4gT6Ag8FsPpP2AHypVU9UGoB40kfYxYRQ
5DYCCseKlhOEJiDz6EBkhOO7No4DOb87yBOQ4WfEbnxcJIQb5JSpTuFUkI1dw/xq
pgMNq0ClUC3Pq8IHsbh2NXUhADdKCzMmYmHDmS7EfptMreiezpDT4UMr6rkk/SKm
DFzhSEAzVIoSHxxwp5U2ezMM2tALDkYKXmuIGkCudIwS2eab3RtKecq5LexFiTee
hFFJ5aFabLD6KgoW7emvuKBEFIIiCw1MGnawpJVjD55LGyMSFzR/Uxar55YDm0Oz
siDPF3ApwwHufAKnihCPPLaK+5aqL0v0DuBzYe+DLKn/e4MfgPQ1ErDFvQzbYDyB
qXBLfCRg53VSF6TBvc9W6O9qy4ncwX2pxm8cyVmK9Bc0LN/KVBQ9NS341GXspJTg
9NZx3PoCX5RUC0cfdR6WndapdG3RWqIWA0Pd0fgPUCKEenuDE5xWApzz4DfP50Qo
S/BIwJnRL46Fx32Nwf6ItWcuSifUMPf4xuqgZxDabhAVwCw5QuO1+n0oV1Wd0vj2
aAzRp08Y7wspRVmxwiiORcEXztE/7xbv9ViQ88aqXAmnHwSFjscN/ph1UFeaEdm9
f46AXOOOpTjMP52RvMAwpcMfWoK/zRGcxnFpB3OBkS9B/kazDMAdfSUutntXupMW
KBbTr3GD8eCEtpqARPaH/eS14tlJJaCi5ZBtZrIjrO4eiC7eXeBTtvfmmoJvP3Qx
MIEMqLKrbBnICP/gRQ+L5PzrkdyYpohq/vSP8OEkKU2IN2kpj3hT5vtR1VmBKZ0e
reVN1TVYlR4nS3W691QwS4pOUUg0zhnZ75oWVVEcnwuP071o5M8D81eiBulCvOg8
FLLR1NQAJDR+Y7Ztylky7g990DHRsTqF/ZWbWifmAarM9KxnD/h2Y3gAMOAhoOqM
U4XmiaoZdtsafhuqbM4KjxM7xpT1A8VoWekg9xdORhMJd4tGaY1tsi5qA2t71HTe
g1ZJ2ZV2tSFyVvtqWip2S1KKIBwiEgXyfhbVR6TF1Y1S3BuHvgmzsEj6dVm5F3DH
Sv9yrYZMoAVGsvQcFABbai264Wf+r4RZFT9XKY485duwQLx0xV4MrauN0fTfCVn4
Mur/h3VXdM0HDjPNLlP/Zjz/NzhJ/JbT4ckisLPH9NpQIh2pdw/a0v2FX3n8ZR+V
SnKEZwwB/ba4Ab2uiwbh2K91xqOC7pKzi2y+Shsu5bKn1R9DbSZWW6lwibpNJ0km
B03ZLO3rgrVm3zcOKXUK6ssnpVDT9FNnP7XMNvOIneFiYZHMUUIUh/5ON7gdC9l3
jHJ4mGtGShAmHN0V+o6dFqY/rcDtpXyPJVu1Tfeyk3FTQN2r6kRnLq58QiOXmQBb
R2vOxiiwaR6fDkMB7Tfzi0dA0k/98ohYEAb8aWiJ3rMk4OsyCTN/Xh8roaFVL91f
vKFMZ2iuh7aPReeY2YhtwW3DXh7JlwulQtzZVr93Xt6WTPQsEXOScGyDooDimhFd
0bBJJMmtF7p/B3gRMjknn0chdjG12MV6CCpzCIuzi+0677j7+oXnL6wUmq2aLT9e
eO8+0sVflBc3vUv0USTcbAwCUv+wsb6tGfKbj5dmI9isyFUm+klmVHmW3qyu2hjK
hJV5ojmdCpSeIxuV6mEf5OXhv3KJL2ntHRz2xEOJV7lbCU30pHjgJg7uUHj/KQiR
FM9zF4+EOQCOtTbY9DNNEwxr5VOp3kWpmBZncrbOOh6uThrKwhTwyzust4hFBMF2
pogg//VMaG1mU7r3qdeaSpCb+B8CER6pejmczekxSCvpUcnHqh3g39QBPJeUyjlw
tl3I+0qz7w9CbERSauOsVTd9eI5LLn1L4uRKeY96642wmLa0Qdkh4L/BBat6QxKP
Uh/x6LE2dqAdeM1yCPcQlAm6KLw8RfzJ+Okq1D9RqkAdo62QMo4DuosEkayGA37x
u8GjOSI3OcudN6z6A4q0L9PiMdPOLjgY/XvzeSqxOiakEgxLRnmWE7GZ4JDxHJpE
3N7xaD7ppS21IsuCGqy4wajYSeGgeZJH65ARDHw8qzA97v2PM+hF/K8jWTrFZz6B
PsZgO8YARhM8iiFXUFtWr6OMfnvWvW2paAWBrifAzAQ9IgHN57jRADBrisqE+ntO
qiaVy8I46D3k8shLeDGxwrRIgfPP4wCieqa/Yiyr6bG1QkJQLFgEbg9huWjqg4pX
oSzkor1bcpjlXaZ3v5F3oDmMszb5t9p+oy9E+yRFuY5BGX3Rt8b3DgR/WbfAYl/f
CCLXZf+G4CubNG4/bb8g1TUv4rmVK10BzMpJ4Q2LIwxRTzWq6wEMmTa5P2v5UMDD
9bQm2G1N5Mi2dEbxTd6PlyjsZLSP+RAkjQ49bNTbw+0EpmZWAVOobpXxd8GGByXa
mc7nBulkNSAOqD/Gg5u4Ano9RPoRM161+YbNxEBALrosSvaUsfm5gITAYwCU7ivN
TqnNEUVKzCzY50ydvMbZmQ8aLNDx3X7ee4SpyfcVB3ZeRKSZK8K38vzf6NMbSajq
1N2mL6KWlLjN3fGFBCklkXb9x7TX7Km8Er920GGzaPG6FGlAAL1wLhFftUwwtADP
RCccMuYX6mbRTnN7V3zcN/Ny/i1GPbs6bOzi+bnXn5vtbgQ+nRR75DxR/O4a8lEV
+thFMQ1o6amH+OVOLicsuJDDVqbaJK1yOb8vzKSMlPzYR4B2M2V/T/BgAn9l9Alf
n+KCtLD54qSGTbS25sW38bckwlflZg5DDG+uAZ9UObImcz+aZuKMYoT1Bocf8a5q
1U0lOjx/FpF1qBOmzsoLXX/uO8MHF7ZPqjjHq8kVZTV/XyllGATJuk7JGbY5uC3a
BR2/Mu6dHl5wBOoOmVjXwErhOQmJnXQNPPqwmUxzN2UlmchbAtu0GRlM/osek2jQ
aZ8TqXe0woX0Ql2zHSqzbse3eiCYJdSBMUe0YhJRtB/mep6Pbgmhp7b60gs74NBb
BW26wVly9XuHo8ZPubyW4R2rLYhoyCH6bdrpNc1YsrL19lf9ibnDMOK/WAeWr/t2
ya2hTltTNOUBqUzr+0fBPP23RQaqp/2O95OgCF96awd+GyGRfup4mrxF8IZ44/4y
TXdU4ywubFtArG8o3kYG6x826zYGYuu687QLtnwFSbZ8DSjiWEPsDHCu7yChKUcH
K8EC2YrHIhams2kkwOA/5Ks2o4gakxWR/KOF3V9Nk7Piz/kDBF45TQn/fmas6xDj
ZWb74LRP+aMqeFRmAyp/PReQ22JIExkEHTJXPG59Nxm+p7CouVAvTcyFFLsvXeba
FWZcrT2EkVYG0hePsLoykWNxl723zuDZnkDYssOyidfQxlaUlY0XTYYD+LKUEYXv
rPlfsia6bCZshab2XCxkKmQmlNAJ/JUrvme4DGXUx+1x+EsZ4jC1arjboqf1/GcO
NKAOXNw1xKJsxy90Q0fU8aUwL3ebxsZwsxAB3vr5kPhUDBccosad5t43f3SjUabc
aYK3sUPnaRTxg+7W1iyA/LZDlobVXZsiVWK/eIenI22Q8ha0fErvYbzHDmYXfFE0
LeVGPDnyRmL1NVkUfThWJtJ/jnpkxrQcCV5ESeNqiCS2e8guc5hIucoEP8a8SMvZ
tt1aGJvrR+vUsY4CdU3sIkk8VrzHYkHbsnmjnMSRYECheGHZjcwB3XjGBd5ZOqXa
sWBFaRBjR2O+a5gOvhjPT3YikfZ88b53+Sng0PJied2tYhIed8+PuoCV+h/VQuRo
iuu7u58vAXDJHf7pD//k9W6dQPcT2HVrhnCNXKaQ3gfF1iaeo3+hBbJmZTGm0gMR
/edGFyYUIrsbDsR/lTfBzdyVe91NR70fpEfPNadnH8OXhWDjFOOw56UVt4PvBp0c
hHykwmtyjcGNdBu0mAhx7zRKrz/p6Z/Fk+NNJMehSiWwnjoIBNS+LpRefcTl5jrQ
R5UWuNRWaNWlDCC2oUyXplpArdg28dZrPzMZgzK/YwUIxia/ac82Vj81gRMeHfzK
U5idPSxs+Q3ecq15zT6GJOWoqeR3b75MXkvU1QmLDPvM0RAk5IN8M00hBoMRbC+4
SBri53ww1P9isdf0FtpU4LNx92infJXsLxWff2BTOdb0XyAZ9p3QwwwtffbyPt5T
F+ChXcnd6CubXKRfplYDLLUtkiajOWQPVLyekI+mXFeT/n6+DcEHqqouTGOwgo/F
ZRsR/CZgI4obW5FJx6eQArNny6S4Hmu1jJB8dJ7TwRfGF28fi5UtPKfihY+M9zzF
4Jrb/GYJ7djRDV4biYvpK7qpY1IRl/0ft1OVFtzgnq3DLHpJh9jks2n8X5zALnjl
JTpvufSmyrDCTG3L9Q/l+dyB8Wu0hn7ZaKtxKhFDZoSiYD91NO2ZbZ3NtL5RbCWd
rn2JunwP8UpHBkHUefl9T8kfxfZtVeH2iarNtu+Jl+xl2badOxm9x1GEO/kgVawY
/nMIJj2qg7jLMAcWLscZL09hLRwEJhh0tS9y5ytMJCK2RIOj1YZz0UI2HEo/KSzw
naIMhHJydTWZWyfJQLBFahUHymZhnfbhVhjQjd5qhKqkh1mDt60D62dvlnD5gdXD
WY1h/IAEtfuIFEXpjietskwtqSsr/YXP3LlB3IzXVN+9P35W2qlrrLHSKFOfx0o4
Y3Qg/uYjk8i221eHtvXgTrg5iDgD/1a3Qu0uWvsb5Xtf2YazyvKd4sxdf2gdlKXO
Wl6GPAdj/ZgPKA5PJeyPiP4mPJGqNcVrlcnEvel+s1OvaFvN++GtY2jwRxf+smI9
E0wRioO+bDMSoEKygtjYSfCCqrX0zSSaAc290k8jbDkgup80Jz3L0I1d5qgA/GzO
58n800ksbNJKO34BfLYNB1I2Ol213fthD3b8sKw4ZV9zEJJZqVY8IVARvacMCEsa
w99IoOvWkzdAgqBTYE18N5RHcHCbzRQcK0sVBoSsO0zdvls03/44f2DKoscdw7Hm
uHsr26R3c4G6lxU8mVkqWd5+w/KHWR6OcLRyUbRui2f3f4XAkXNK6fTFueS0GMBs
DgPmyPWDl5cIW+vR1bN2FXe3NHMDC6gBaWdkdh8sPGyG6r6FqYPdRgrzDRlOM/ZI
B01ovVNw920yTlrtlOLFMu48QAx2jN5K4tCiNebpJfjlggDpBeHSC7xMLvOCnY81
W7JBuxPCRbMmZt+gOqVwRi+TACNullyD58HYna9vT6BrT5a7NvZ2gpqteouBiXe1
zk4zvNOnRapynOZfRXYrOaiJfAVBRDb44SzbDui5GTpyhHtI68WfoYTffmpE9QVy
YwNTYIK1IjjreiAPD6NKzPflooJnDK4q3l6JKhZAj6A6HlpyRvaSYUMLC2kd5AeB
qr8VYFnSwI9RgupgzWS62rUZIUcOoh3N3uVrz737ReMH6+Inc74E75Ao6ITm3f4h
cHN3uptnT85OxQh7y1hN+9ZGMqzsVK2e9fKYFwr9Fa3yiNBR28i3qEO0ck654S0/
QNcneZp55JnT533CLEcNhq2v0YzSF2dKt/bvVdFuAnHENmpZ154SmtEao/chAtPL
WD3hGCWcBFmA9LUGtjcw8/1dlEXKuXtHpOQRGQNC+FhkVNInxDOr8QfnUcrhoj8B
zQNCsp6ODfx831WKFj3i5BgvkUreGXA0IiOPifehFosARwA8W+RWurkqSYGV00Hy
K2y33ZZ1OpBswibe19/k6k15ujWA0ck0c3zmxF+lw+S191eR+GCfPUTJ1X/zABxg
WHGmlZLnfOnTYOlwxLDAMu5NEtcujU29270BqNu0Pt5eSApmwUW2LyvfolSihe2k
umVp+kkHXCvbpyVRbaPJBpD80ivxB3iK592KEnS6C5SARsBEQIdJhxpwa4IeS9mj
4sUYdjtvC6wru8kRj87wMvZ3z+9SYMweImR4zTpugYSyinh5pENxZqsY5lStESM4
KqcSscXa1/WKBAUf6Lhw4DF4TmEGNRi9ZEoN6gI4E0q43tFwSDr9wbWjy1CCW2me
LHXYtEUU6lDnrz6iO8YUscboh0PlQMdMtfFRzBvLmwHb+edMDG/U1tR3pvjv9Q+v
3jNdnGhkI9Ys9mlNOxDmSUJ4LUjo/9oijMrXQRI46V0KWw2J01R+il2t95XgwYK+
wpmu8bI32HI1AydKoCpfhnIDVBPeigdRcvUIcIUxpVnNSUS0ggJs1WSz5J+ABEkt
DimIh/ywehc03haS7IxwIHQ/FJRZ9Dv31AYjht0j+2KLa6A+KLYNf+tyJmMmw1js
1btR0cwsK9gUSy2yQpEqH2AxJWvGLO7GEhXlxtuFVxU3GPlsiCchwneBMV66Qy6e
lbqTculbY1nILGfVp743uPAO024wtXNpRSkUwZVuSGsQfi4YQT5REeKNFrBxAZ4L
+q4wbs1CCJvBzGDLsF3CYNRpf1owaZ/EAHN46Dy5H8Dq4eyYyW7OCZp3hOE9eU82
RnU3nLz1nKE84IkWQ3Un9IfcT4bdAxKj29IdB9Xab/Y92LvtuwPHiyBZXbPtfm9A
0VEYe5Lg3iBNdLu+78z3Z7fzQW22od0wtaIRvM0Aqbz852kss27rV6J1OBWbASvg
KnUJc4ZVNfXXGEYCJyUjuu+ELJqOcOqgRfrbgof5kx68ke6U5zPBqv5gwV3Oo83U
7emJcqYk2A1RzP09u5vjCq3WYFWeT2m7vhHq1udbPw4SAyM7ACrEEf3XzTclYeWy
wpM0DjqILzjdEJ7htrO9M4+nxphINHIhWm6WSNJlroxZSYfMrFEuRT1z7+TeES6E
5v1UrUamHNw2NPNMDQLHXNvOIt60pcKbouGdUcmaKj7oLq4lD01v5KABJzIzwYXc
aG8XbMHwKW7gPGm7FMy52HXM/Vu7f9RgiQBtg91CN8UWtU4+AgVpRROBdigoEGdD
ubn2okEscMBYSWWn15v2eOT9BY/5ywylp5jMkHMWwbGGVfspomN0uqRu6+HnDauB
/Y6G9oOZQY/wOYIWuNMDPsby5tPTEoQO4TuG4kO/Z6Zug2YJEvwU1mYer7P7GBUe
h7pt5ogP/Xd7jLvxLlrE/Qv+oF3R0xzP89u3eknZ4aMFPcaXvqgZWrHPEC/aC4vP
iXOMS//3DFObmESTrxjqne3jJAkvWOMq625JhxGOSEa4mEWJ4jmhYM+qkANyfqHn
pnjeUbS5MNh+66j6F0ZY9DdxRq26QmFFLvxG3/oNE0YR2EQINJKOK5fEqdc9tXO4
mk/u5F8nDJm0dgGAnb4c9875nvzn+lMtSnMcLnDLEP/bz3GrPB1GVYBR77ySi36p
dCXub6+/rfGHgJ8YiqAXllu4cukoxujUQYp4Lxf3McM0Jwq8Ukzsuc3du+Jd7Z9T
GZhKWVV/u/B1T68Q5PWqZRPcBpdBw/ub+gjhO6JPeKe/rmtN0gCyTKmByQogRJtD
Ub6QWvCItP+Hwifmx/fp6B6McLHZw4HS5aRYTmLPYt3aeu2nZweHyFmQRlssMoBl
ZjBPdzewE0g1BsFGRp0Rg13+kGf1INB3osVx9iguJ/5W2mI9mEdWQgOuMqoMRGpY
P8z3LMewCHEcDINloFL8DFIde3zhWf3iKdHlfVhBmFAz/jKgS+29/9Ov+CTC01Je
VLOUD2C5RTNSDBxaZ5h01CFoag+Oe035DXeNJczzxP+9P+WMZJ/2xuNlhFrgUExm
aqchruHd3XUzwacKP9hO/3BbR2CpPfHrtyxbmQHn90JB4s4OOK3FLWtly70sVdNc
nANuTg/LC/T4tF6kg6JkRw0yjBJGpujC+Pjav9YGOJgx08mfEoSkQarGbV/E9ipE
zzKNOY+7D6L0yWqJ1puN+wWRukmj/dch4qeoW31Teyy8Q5gVP+JTF5Io35p6d50d
izxunFnTdPEAn5RLB2Si4Yx5Q9h46WmdYHj1eAyNCkyW7Djo7qE5ABkZLdg57nlK
RoHwbbDBQjz6u7nzcTid1G0Ls9tFswFcoq/oqBk29sKTzauJ3zMKkmWKX8epTGax
Lrxeu4u3CImVtgfeuGI7jXsAgRGfMKEJkyjGvSOQHPPNLF3Dqfz+tZNg+EW6hOlK
dm4MWJ0cUJw8rp8elPfVnficXTRDlO8T/iWeMRri49zANyJYN8TDBvZfSJhcUKBo
UMFlQT59jWMjWejMTCISRDIUoUZ3va3bT7IE4Zy9CCLkDmzSRh+mPlroiEyW3cH5
dJhsh9GS5h1FR53XjJ8sEm++XK8N+mqK90nVZoGfUcvsy8EOj1TW64duRKvTyjT2
xTvu4UUDZptGWbXLtSdlvKE8Q1boq4iBRNoAZRuJBGiCz9iTWhL6YNIavJChprJZ
c7yP3+KzD+d8iQzt/D4pYKEOAW4DQHIncjQL0C1OZUReEZSR3WcwT5XBcndr1Fch
lAPKLnjx7KeVHGr5xbocs888O6kskDym+g2H47CuH0szAdalGmTJVUZ03DIH5q8E
oTswAsx5YdvnZxpBjSWa/Lj4M5GeX1KAByOBAXcxiVBg7V+o7nROwEh00DpzHA+A
P3QRtLUfmUYhMvswwjqU4F+6ZefGFq6sn2Zzl7vMr0XQUKXYuHoaw2mB2EYh49b8
8u/N0l1mGWKfo1cWGe76YAfAPHo49FOgWA4PWHZ1Ur0z3TRTB9iG1UXbb8bD4ohm
x7vGA45mFF4D43kzd9tR/FiQ/ENsNHpV7OKJh5r9/0B1+gedMJhgbctqeMI1cg/4
cGtsl7K+2kFFVXh+hGiv9AFvNiCQa0s4et1NyOf3RGytPfKzgzEnUiavJmWI0V9t
+TAqWjVq1tcDTJKfm6XBphPvwaXDztpMuImZYhggVzAdb6WTuKtQZ77havBuDh/q
DAOCF+dSziu1eDyse5KvsVvoYKfvgoLGkSKzqS9Km1QuP1wzjpk3jrtekjD59Pqe
0TzOjdeu+XjXHsE+Jipbi0hw1i1BJAT+eQffOFPnYCcOR1+MxvnJQ9U2SO5Ha8cx
GBzH63XgykNyS5g2RKslr8vDdVprliAE6eLh/n4CNF1X5IIiPKmySxnW7pl9gvIj
ofqS/O6ymqSkIxyuFTlLqr9brtOPthb/Wy1Tcamb0tIX34QO91aSQb6jqIoQ58/2
i7qEIaNC2jJPRvV82NPfNhJxMr/dhhJe2UWsjowDfF3CupYzYZP8giVXGgtJ+Tvq
9FfAeX9Ggc9vzGbHwSMybgjNq9ipqGPShChuKu9E5VhtzQn0WTaQ+mdcruwV8B0X
+Z12W3SRbhIQzNv/cO9HhBIIGeXwedFeNToBHfrhL6Wc1bPPUyuOwiVM4pA5lCRH
ePziUrXwKvPZuH2iz5Fyj6tN4gElm2gMtZzoGuE2y3YuebZmtqjQj5Vgya7QKVYE
7fBAdSQQd04PpZcbr5EFxniK5SNuEDNMnIXj8nWB2cm3yxE7sqVrBTqAlej5Cq7V
O9UDeMc8nvo1vWoSu3PsBc4h3+X136XabQCb0t3anvgEj3yqNQvHUf5plbouFpa9
DoU0ST5KHCEDVLXsjvvPouV7JtpfXYFsWWKceDFBC552t5YrlBvEdr/X5+DQ8nC6
oAbk//HHaExxdt9AZmidbPrHkIp215nevhclgAObs/jjuK2qUv0ovulf6+BXlFCE
Jr6Bs2zKEwz8lOzJm9mv7Rx/6ZNYUh1Px8WRxhniJMLco9K812x1wIItFeGkqKHY
1l3+XZJGl8PceKg1uoByqR1uKfwNRIVtuw9QCTcxuc8dI9YneUKRdFRMM23EsLPH
b8WR8adv77Qxjww6ADP1W44mIy4FCazDc63hR2pE6k/9D3BgSNGMV7ZfafpbVndI
nMwFEXxzsgBS58QIMsrSgxh23eVyMtfyblDrMHNMNWfvwwo7PbGadK2/TMOaFWe7
eGMrDtQFCZOaghpEy1PZbXaZ8euB5jcbOYDJJyi9gGjCFDYjLf+UxP1v9+XGI/ts
aaXF3RvismGYtXcPlMkXMCNpU3vdcfI6FE/mY9Iqd+A0hScr50BF81c8CDvw0mvU
ZUHBvNlsNs6f5dYg9vtmO5GvfayR6iUU7eizZCbr/NCPiGbHh2CQMYkFvIhi9gXL
eojjh8boUdYVr7xNDLymV9gCp6K52lM7nNY2xJBv/3kw5QW0g8M3+f97KBlvHuN7
+J9VCa4smHNvk5vW7njZhlTU5OYYVXHn+dFbtCPpdyzu8GlZJPKOy0DIH7Fm5i2O
Bwcfab/Sjj+71Gco3zxHHCGEHhDNm6Ky4M5oZym65d/E3q/QTAvVhr95cB+/rCxW
djtcqzEwgBnyx9pgrghVnSYdubdlI+W7dn4OYZvDMnpu45TQ9MmPbLfuXT/d68fz
yiMZhT/vzp9VjIefF24ns1Jdu3zy43DAeuAXpg/G2spUJmSh/DHOkDcDRXeCQSwL
QJhp/Jb6rKxzunaCddlxIe/TitznbKAgx75cHtr2mvhcarDF1q1bj68luVa04YBa
wqHsPzQpKFHouZqS6rZAfxiduYZoD0vebudGsRbDE/l9OpGNVCOtif03swIPnDBs
pWaknd0i8BUSdvxLY6p2LFZKT2TGA0m3Y7g63rnRC9rLc9sl2meNrF9nifGVDWlG
9XuwmN/LR1sDZrdmpH9b4jp3p79zTDCP6YDD//ss1LyEQaVrpVvOsXLKaqPYyM2f
ufm6HYO3vdM4t9LOz2I6OttdTHQx1WoXOcGu5sTxTC1SbJO9Zrn9IoLVE/E/mbAh
4S/7o4gYxpET5ShYJZV8HVB3aGLTFjQjXF2Sy5qb4PEcFApp3ZbR/iIJWij6GHHn
by6kc8yVoJ7sLJ9LAaO9obSnEwnVh0rL2Y8FDip2fI+32ZOOljlnKnp2+FXFwdNr
db/6EiJOZCv5k+t7zTo+ZJSZQZpGZLodVyEPtTbkYvlJQsItXQ5XNInau076xdsu
GP03Nqws1tf2f1WvQWsWVRmdKss59S+UcuaRHnnqy/bqSIBoPHQjIqddKC0A3Z9T
dxcoBNPCA0mQvWS8zckZLb9y6vzmzB1gEgkDQFYxxrPk3wMFZj0EhKvrYfAdQNCW
eSuyTgM3e7uCRHjv60JItzKrPGjPOIwI+i/QX6+gwzIwforJBQU53c1PJZNST1WQ
iFeNMXLjVxeGefK49o3d36jjLJCT60r7mZjbBdfKKPU1k1mWn2fa2kWyV0AJf+jG
Zo2dMCBwfJAijP0QoR5EbsRw2wxbhYUG/LMu15atjsGf+OK6/Z+Z8AYXe/UtRYRs
McbiwMr5H3R3vSSHR5lVVfjSGpjfmjw10wTQYCsGbSUzWXWdjMTvLNRA47fV+7UI
E4k1Bu/8/+2rwT3d1nvMhBNFz2WCUDUn/Jsg1wnhGWswknRHGLDeQu6MwfdKvbbn
anm3EvahwtbKcM0fiDLNF6NkAcIhyogSTFpIMEl8JO9A+JXteSE6ONfbTeAgvoM2
JN9bwIbON+3giuufLWGgvwVDlWT3p0fY7juoO6m+bS2+WWAw156qTRWlAJWHl82b
FUchGJ42IHyG85ndpqR+nhXTCESRniFy619LQKHeDHavbU8MUPdsjgf9daZHU1xI
Y2BwIf3srYstcdp9Ufvo6iMGlhpUWWFp8wyQ4hIH/fAOTNyh22+GycztIBP7xIg2
dPXvZKddHhT8Ggrp//ehUpm1gR9nGSgenlfhZ4tFOQCFG2NWwoGG3PTs4hheOoW5
+Yodt97JlFJs162HequpopfSpKoRvC1vnnCXOXAauBkmm4HPwk0vV5qz2OKAj52F
znx4WmvGcY1dMBHvpafC/rr+84sVXqsUe2w2P+aHI/wasbYg9ejJJTy4sQhEXL1o
utdZlnUF7zb8v6wpUFNNaQqAzJFJKF3ghJy+rd9D1QpURGIG6QAMm1slOvvs0vde
Hsa0N+CFbq0dgVVVHrFy/Zj4ywgCDwpQB6oNATRpj0yFWSkhiEm8H91cdxApHj9o
SfEhrRI3qU6uOAtPv8RGCK6yeEAfsnbHMPDilqUEtcZj5KIC6I4nJc3tAXhTAsaf
ycNOK7dzMvx+a93eat6WkdCWYg5bQxRy82urljMFIAgM6DLrAPXw7vQJqjy66Qtv
d8G+ncRnXh6zvLnLIAlMKZ3ogxp/mg2g3eWIkNMxC3LSlCXMFbRTFEPOKvSo7a7X
BGAopt2BAAQ6KWn3II1Ds56Ua474RyLO2qoJmHipnuJWXEaR74BZBCaOYTmQVSqO
nH2zKrqMiRbgSs1rZJBHwSB4fEa9t10BZt5d3dMHrMhm+W9l2D02L2Ccjvzk6oub
V3TG83EALpKVqIvH1VXi5l0N8d+yqAbMP/+i5XqwPdHR0/9dxt++KwbYNkZWkQLD
kDJq83LUv8d/zXzGpd5ph02PHkfsPCMCzQxlCrjFjKLBTdh6VfJGyx7HZYgnuWLO
NKFJkYE02+e31rBLM+3OLAykhlhkdUxyAv4F4okLOclDEh6fbpLDdS0If5G5lmAE
/TSjPFBqc0fWc4ZoO52Kr5Wkp/JUpaR7r61qmYTo/E7FkxbmccOw86XNafy7CFie
9BVbgtS59oSif3P+nF1Si0V37V4lg3LzQSvaCIpsWSZguELhV4rLSpFitlh3rVxr
w58GYYokG225Iusk+zzP1R+phZZNGw9UEBPlGpoXwyn1onW/iWOameGVEFA4LnOh
5741SXyPmToQyQHNbp+eLl+70K243LzuwJf3mWOmgfL7gGUfHbcfvH7sGR9KLOgu
fSwymaUnUcknGe4t3eE7kjoiOgs1cINNBg+1txCzxRCDu+5X8c+xYrPL0n8H5ChF
9tR42AflJiJXNUtKth26P0M3Z7WXGLafVqHw0rQTjNoI7VzPZ589N1e7aBrCQFNj
A2WD1J1D7VZdJJOYHJhhm0hLBAUzxFiAQzyMIs59Sa4f5PWw03M6ZbxOyJGZZ/SN
C9E4OnXxJffXYltqdAvudL70GHFdKDqECsie8+tB9RMXfNCcKhp6H3YH9Tri/dz8
EeXT/3W6D2SHHvLsBWrqlSI3VD5APL6a2F1da/Ufq1LdyIZVEJKRN/Mn6gSpy+na
3X7IWOCbBQQgCb1NP7ukDHHp57drQw0kMZa/MK1UsO+9j2B39UQBo7wVCrX7JR5k
ESAbI+/6RvIdjUVgkzAVCKPMoZkL7EuE98cSKDBLNQQfkpI5M3hpHKxSlTu2rqA/
hehggVCCWuGMOiIeOOo9RTnEpEvziE07z+TTr+r9qEMdRI2V8RiY2g55+oYwR+4V
bzLTbZDL6RnXEvNC3ZDCf2Sy/+qOEw1svXPbEgjFKF9ivCePDymQpiOm9AEV6qMR
6JhBOJsHl53WJG4hCpPcXSt6NDvA+HrxHBkFR2V4OYps26DGNZn19sEvLKEyqdQx
vHwoPRl1riIQkogA5aHKrp1vR7eQFzNgszI4mAbe/pTHvrCrBCx8WmqF1iGZ7sX9
zKm5Xy+NFPUMeTp1LcfZoXVuxvyihVKj6Fbe2ZCjVR7p9EW9WVbPKeoDBr2Jrtad
3ji4QcTglGY3czQ1fFMSpEh9IiVG4SN6iGRKcH7bVnAnzgmptHITQHsavihXUvCv
16T7lvMcS4BV7b6/jdhSRzIA1XV6VZne3QRaZTkzgqF/bmhY/sCk43TmXjxyJlu8
WIoZqJbWb5NbDebgvCy8/R3Z0HRC/yC+XE+RHuRnLDeGplAk/J0Ao1juSE4sWTsI
6+0K2w6NUpdBTd/jUNy9K7P/YkMs08CkCmTku7fuzJmb+E9BWtGh3m94EYmcSp+b
dDl2ym4jTiomBuF5vVFmj6GiWTEoyXdhC9p4N3KsAAACKLSGlTIQqoCkJhLti3Vq
SH8zddMHTGM4e3kzQdtOj4dZxXc+RLdBwA9u7E9DjAz+FkYjemi5sskhLPBqGa1a
tyMVf0lUWCdwApfpZkqIiasZnP/YgiKu43BAW5Mt4UtgkvU640WwFy3LfTUWiB6Z
gMED4ZSD8BSDKY8TsJm3tUlQhxNQ1eOy/6q9VTw5cnPXvyly2xuvvMRCKXtXiR4b
h3EzJNL3CKQ7xTS2XgRx4ZUXgdF8sUG3zMipktZ5blpmHNsmKjB26Ao6Ejoph9+3
53XxOV0aj7vnpYJEXLTfwMzWS4JEYCo48L4Li5KQN16P0XDzuIA50LCzRu4gNpDL
gA/GfGD2c1yN01tdD6ecKl6/9WkZslD7TdMAo9rO2qJnEavRKCj2vA2+hoaT0Ma1
ilGjTbGTDUoqZd6cLR+Py0Vd1+0490NzPZ5glmActSB2YN1scXCYUvpxfGIkzJtt
Wg/IeEnOVrRWtjtDCoFg+X1qsC8ZdJQPuXjmkXFT93BvgAza40hQRL39+BIMoqgQ
J6C0Cy5DRlYhkAPti604KJLvv5/u/E1556Xu56CHTyIkcwGmWlW3GaduhapLz5Wg
aoWKxylYqNIY4VrYHljbX4jXgqe7wQtWWUIUz3me2KIGIuKaFhbgY0C3wlVwphio
U4k1SDaAgRnf1q4aVu0CCZwotn9oYAU/x9hyhuFCE8wyc95PNa+FATqA4h6l+1eV
uMYu00eHRTN58pDM1J+xliG4iLlP/5cOHELPL0yPeOMhZx9tQJh6emwjW/23aI7C
KfPAmgL+juu6fHGY0jzNJmRn7/t/d8ZB+Q6sqNlc+j2d5QTGFIN/xDeBeFTW3aHk
t1kqPw0VW3mmQeQlQbVkjlBfU3iK8DvD47yFASvjaJyxLOj2Gp0wjvGS0Fsy/ILR
FWbjgx7pphFeRdGzjeLcUPezXumTUI8DKHxdHCM3ES+0oQYAim20iptdn2aKSdjb
RYI9HJ5d5Zk5N8MUlc/hQgCAfknz33hBASJ1Y/jOuoMpHcRDtxHyZCfNtHVmvAuE
OW9kpGvApZUf5w7Ym/k7A3PXGjKDUwxi+M8YPPpHnSUpvv0jzvezDfuGOZNhcXmn
yD/C1ZDUXjrXxvKnjhSu+1TC8J+RaVaz24rjQ31liUl6yPMt9jjiOoNIV16RoEJz
2vRwfQ3KsWxWigQirlyVY2mReqmlXoM/S7u6+JcKyAs2mWPnlpGnTF35tKkBQvtK
QzMHYfq7CZjwwo1HBFdfLimYuBPo5ui8Roc9RulgtBrlmkcikbxCuQ8A2F/NBQvk
3vcF+qao7pHdyTq9LgbQdT2Jc7xBOt6ow3Ub3F6ofRn/c/H8tFkGiVDrR/eNxyFj
MJ4CewP7N2ZMP6myE9Un+p0LWrqKgEas0Th5zUmU/af/4kfIuladTqOr8/HFP1Ew
WlxPVVBrmmfszITLCcphYKW2yCN7Awsl0TcBxZnQGdhyCM6xzXQY1Z/HqAmkbwcQ
BClByBXhmoHDgmb5wYeHS9zoyd2X3KBifi4r1Bclq6ANtViK7Gp6vJ5co8kmr3qv
lFc6mbBfDvrS0Dok/kaV2shvWZoVLJ85YTnG0j4LK3IITAt2N6Wd1DSpFH9CvnHJ
Neu6VqbWYUkk7AsYAFbszKJ9Yz3I6TWdet5QkCr1mtleTZ5VzMM0qzJSx/7DBFUf
DvXxYteUX3Ilt2srz1ctI5beOlait3JL/KsATgMWhV1Uj2H0DuxZClPtwFfhcrFH
1AI1cdBGcSNyo5l0uKZtgjmhwq0Fzql63IXCBQsKXFaDvrfA511EX9ayXAwHQ9Cw
dFlWhAS/+nlMbhDepOsC2aVvmA/zTfrS8hj/Zh9PkiD1nTxy1VZx6kz/AlliVZtc
FuEv2kaFcmAsCfD55nqJ5mCIMWV3Nf6FU5QgO3HmSfRelJ9WtGbwaSRJz0YETLLy
bV6r/rXtp0xdB/fFrs/MiyC527Dt/wJAhHUFmDX77lZQN1sRROgmlt/Z+EV2xYU/
StKvS5eeGdIY9vpfmbLvq5De/kTOaXGXDoD12sV50wvNqm9IAWTUiBSvfpbnkZfb
UiJhaQC/zRztEcv84YUV/etDHDdM4hYnoQLCqYFCVDcqFo2zrT5Tno64JtFf8mUA
tgOe6chFyMWkJKBGZGFWLl05W2LeWEd2N6GZesjadoy7AAdx8iXsedEkNyruM28o
SDDG0TzSl31UqI4NNZ5USySyJM4Qwpw+GMqZOs/xg2aSuA6vpQnBFt6ChHQFGQkU
KmUNQDkpP2EEzpSwVZlghu2k5Bl+M+GO38DbbyhPapTmipwzzQZs+ZxYYxmgfwdq
+WKNfr2mY/vCMrR/WwRjFD+N2IjtOBSkRwPJy0GvVLvsi7wdcVMDRzej04LJOBDr
g/6hhAgJ3Ea09WVmRoyxOB5EaENOdviSVNIuTsdcpZHPGYgJwx/DSfAyjW/Bwlel
PhCCzKFh8paRHewGPjn9CyjkNZBFgwlADXW2h0hBKiayTVUCc4sQeZHrDeNaCNQW
o7PGMgRApk9fRa6YMyYFGqJ0ok67TXvhUAd6/PgaP4H0kTBa7Tl1//P1ihJELVFr
LsC+4a8pKSSr8TlkxNfwK/+zifCqiIiLX0YnGzUh7QXAH4K4jgunHFjUnLHtCHkJ
hAuhOrPKOECuFOToECKkR1mxewo57JlUrKFYu05G1mpehz7qwhWWAZJBo2HA2j7Q
YNTao4muiO7bBJo68YsEqNoui69GT7mw3b+8RhCHeBSZ/OPl1prHU+/bMq9UY+y4
5mMc4rO2SH+9oN76THJPVo/bjurwHOC95cw6XA1Vf80qgbb0oi/vrdGbANgTD7R4
BvzHhdnIV45Hl81vf8gXZlmtt1cVm+xYj1FLNoOAWYgDEgyTbYScfI1tBP6lNgzM
ZISlYKcFJItM5E3/DCvXE/4/Ng9WX0kG51CpyCNxyjT7F6InO2cInTVBnwjdupmp
Vj07tte45S2onIur7FH1Esuyh2Nz/4dviAHJclYetj4vVu6pLyOR+d19PlPvzU5s
4+Hi+n0bSMAOxCcomPWXajQffiGNR194TATvqeC6tfYI+au9jMILttXh+nKFIGf4
kL/gJuA6uGa2cFfndInvAEavFJU1SgokWuHzGd5ldB1fKLyEEE76m5Zccc6avLLz
hv2EAN/+fCbPCoW8UsusBzSkBd1HVEL39Xj5xEv6C9QQbuNtZcn0EXurKRBBizX4
F+ifeexZTtJ8oZif5L2aQZazP/e4E+CysAjfLfqXbjvNcS/Zw1QDumd6eUING/Qq
VoP7YT3t7vIczydgBBMiSE5H0a+e5dZ7WC5bLxcaYIBEEQK5Xs3DFq+159mANYtT
MfPmO1717b0YGnX6pgr7aOUBj9OIUVilkmMoTsFB9NPUlYh7ACzblovQLIU7kxiW
LcnOQkyHckrkYpB+y1FH/s6Szy8mH7+PltmuW2QIbASTOyUUo41C+cytttCeHIRE
maQX/lfr++fCKd8ATDz08fMvBf2xVPQuFGzj3OQtVhcmhcphH1/PCO20RLaKfwVA
Ruo2S4if8GVxaq6krFWkShkc0Uaei1R5zN1bbS1XGIYUDXlm/tTd6tcOKD2+ktPe
5NT+M4laeSkzVmUQHsfvFbKYwe5Jsghr0RGfTTtYH2xsqf+0NP3LP1j1vBMdjkGg
y7wGq0jkk3luFlMwukp1MsXvpSLIcMvhajbhmFjDNr7I5h5NiZ3Hp/Kgc6S/vmwi
sbDt1XwJ5oAkSjnweN/mlIa4pLAofMsatHR3fmnT34iXHrRQVG8S51pYQIiJOJ2r
FQEGtR98/pXXl+OjLrXDqPbj/F/GMk/24IPaePSWYgQIe+o49JygLccxgWqs2Ixe
MYdoFh37dl8lD4T3H3R4b3Z0Y97GexKCgHOmBUM13ipFwRCV6XN1wjG5bIB8ruqx
PB8AbTFgwEXr94NTJqP28wOFGfh7VzxinCll5pufxFqKDa+UmMxmcRRFv87iWGNY
PGgWHa0NAGnUljupVz7w/BvPVIQPKk3hptJ6uVfdhEnp06wCWGBxecstrJ4mjAV3
VsPnfppOZ0c5tubAd/kz9X8hCCwMtYxtUYRelyzUlhPaEW2WqJhrV0US0Kn5uE50
mSOtnXi0JSpYxMukofmOzvaSoYQnsCFcAW/T7Pu7Rrglrl4TPE6ePWR91Yriwo9S
5jCkqT/7sorV8Xc22hfwZ/ziq1cqFM/Zvo1ADsxP+OK3ffcZXz+R+i+IjHVPXIGV
BYuYKi5mMgOJK1HTjmXYeLQ6SqdYWb8HNrwo9twyw8yd/GOeze9gB8O8IE0EnwJH
OnWOpRIiRKAYmJAaY6ZSiMIgiRmsD0xQR8hFiwrhpP1ev7DbfPbSutarTIqVoPqL
+fXVqsyYBryYXdkQXdr0E2UONmSQTr9mNzVTHZk1s7emuyW4wYfabjdEoDNx10T2
gJKC/81T2XaNScqF0MDzfaTzZ9DApLLf1HPvVsI6NpBKqyHbpXNJrLgAVT0wBlbg
Ky5tNrjhAQFxPMzpeXu3Gjn1JpfK60sXPE3/w0GckUaFkdExcff7WNl5JjR+rF96
o9m5TBcCnoh/a6Qam54fl8AmU4D2vrU917UbYiwBQSjhIFRmW+Pr4qkwCwzs3Qj0
fCjGUx+OYL+EWGOfsRAkGsAWtKzDkFI0qFTYYL8KfLwqHpUX9CeUhSxus7qNOx6L
jM9vDonVpWaMOPhDfHYXwrAiog7oQmDRDn4RMBYTmW8U3pOveE4lW7eHxpsax4hd
KamJlz2G7jcna/WNdhHRlTjlGNQN8vATIGLkomgoPSLP3lR6e+P7pjd2rIf5p4HH
evsxSJfjGLGzw9FW0V4FY9x8vh487qjHYgCJfh53c7lvX31gdNaol8DCESLd4+Ds
XhYfzZemrV/RC3hQMZ7B5wogP9RDoIG7qxtmbTjvQRfPo1bt+mZKmG9aNInnyJyF
oz3uzfT03Bz2VSPiknpd3GYTGNUOmWqKcyMVsarAQWIiPvKSjypcf/WlLvdK5dv6
mjZFUjS+sX3UYDhnv4K7DKpnRfLfwXtSKjpl7SXhWnnSROn+dwdLWdmPkpxuB94R
q4MoCzOh8hE2eQnjeKzd4FjoHAwPPItXMQOmtwV9a0SidiWLLfe9yiBBRvMlhPv1
Zs3fpA5HN6/X8myQyc/3RMLiMrO53LP/H2lVQqNzAU5eHGsUumynIvX3zRx+5RL6
JSZV5LhVRUoa6pedNMgP1eF4eNZNADAjGcYOV8KONzU5v9+0nkuY/90HGYqyA2F9
nrCGumcbXOE1BW92ObLZP5AA0O9KKsJGaIRADo9Xb2i8IAgHCmCkpgqErzpXzAGv
5veysh/+i3+QYsj8z7UthqXBQ66VEyvYwgHQ4eCvWorpJCM5oDA7kvbgM/cC74yw
i6vAyED9OTvClow6jCVqda0NBjHsmJFvVDmuDICtSEli+Lqe0DRuxjBZAPpXJTSH
PEuPaSwJe7gkJFuYWD3I8uElYLgpm5U9mcl4VPsPS0u3vHV7EMIopfncDqOkoQnZ
xRCK7MnOIV9Wt4rQRBX0lCrbdgnuET/rzsaKxGWg2PX19JloQWe4gfJiM6fof2/9
UfZG1MxcPiMn1EDKyoNmshmfke+M+/5+XlJ9GcJ2rIQgxALZwbp5HmvL1/qP3+44
FG3V8rVp2Fkyh2q2I3JsoKTYkwOdUYRqkiAdM0fWsOASInY81q1+4x6JxHfJzOYB
TsF+4xi384dWFdqnHN68Dgpyi39Iun00I1FKFEd/ylcq5gAtJ8a2T7OSh8fDNKK8
s909naFAGo0hU1xLH0H/GiN9j7ARLuWKjStAEc53ek0aPBBRsgZhiSS5oCAi+/sr
vsy4LWlSyrqtWUcJmd4RRFevGEpZC908HCpODPRfcvzsY72pSynJLpcvZviuUQSm
+NDHWNrP7SQVvf+XMJ0ibrKbUkEvhCC1WUjX9xjKWviWj7w3LjgxDIh10LFh0PTM
OJQH6TjkR73hwJrxP12L0WurhRJ6yzsanT6shRyUxRI5diqEuptMECpijk2gPIFe
yG4CKj8fJ8YSNixabyvXpfTJ7lDFn8vX7WZEpsM1zo79equWPUT+imSGT5jEN6Zy
+HfwXKwAzJH3Zppo/PIYqQ+0yQAiF0mCcVEc/JEYujqZP5qOA+kRGi+z18baJMl6
n88G8rvsXcP1OhIJWAN+F+A921SWinmFUhEyyOSixsA9wpbWSnlz+sxkh+qaAn6P
2bDT2+OGl58dvvNx1Sm0SaDncJg/uD4NG2sNp8zPXjdyf0D+C3Qjn5UpE95Q113l
g2s8m0xh7XdoEIp0y084H+VMxR80Iu5PVLOGxtb7TVKvP4gha2GlQlBwmTNhs/Ke
Uuf16vvCtg5fkioEcAl3UZc43qFvflw/YJs9j8bnENg//K08G6Eu1t/2ZU+TAAN+
183UF8leBHmR0G3a8UK4y8jXJQEQOeNilqZ9efcRkIBXGGN51X0EV43PcjQHG5yI
q/AISnPJwtnP6SpeRL6USnMU0Vk+6Hr1cFslcRMHEwsSXrRykZkksVqBZapwjXsc
ZitCnmkRTMLLYGddT+0GiPV23nxiIaY4bxoZoR+5SXrhFYi9NOj/aVsyU9X7Ox1G
44VOKmyALTiRFJgttLAjKP8wRoBtZzE8iUsq6fBeDpMfvX6L2NNXv/aTKWbGWTmD
zQOVLCFO4WJPsDdBgk2MBDVp+5AIYsqhRFMldTWMWVkCY0NlHxeX7oevH/xg2ptx
myUAa5iaY1BaK5SJUPp3cyAVely50uFObahCKeae6FOBtPZOJWQJxu5runzpwNKH
PjVBnzJhn3KVEI0w/0niYpOaDMXjZsy4RF4up6qAi06W7ClpNvTcQyKzT61ibIcM
9gL3bTrFqYPQSpnSl6CQL2LIEbe4w7CbrwJ9ojhWzJQ3akrAz4HGK5PQ3uEsci+R
oRh1KTqGEbqHKuWYPfuvtbhu+bOKFU/6WDxT9TradWtdS5qM4rMB34r8iACew+lH
ohnBhQIZIoiKhXv/xsK1aHbSABnyqBa4p8QbmjgbYiHXwGwzkw0yAJlxlsJcp/Ln
rJSY+eOsQuRi+z/bcrMtNu0PKscKnbm7CO8gYW1LpNUh6hPCMPEOqMsRR/EsSajR
T6BThYnqwwqpuVWOaTB6VT5cZa4XMX24kVEhe/UWqduaFVXssk/Z95xy4g+aM6j0
6fdwA0xmI6jf9sUBOyPAkNn3htCuecE5GOHSmKba3bvpF4EOSqe8EeOcQ+VMo5Fh
O9uB+0yGJ0AbiQmahl47VGUI1645QliQCuB9s0Fp6AhNbmMHcUE9k9sxson+ZQY1
xitzKUCxXHbukNg7Npu71t5MqWk9aj6NIOm+QIFlkVzJNi8xeQMYYpsxuLZHih1m
4J2ojTSZnHZtp5tqPhAJVQpGQXuMEwiHKeXgDToM5X/QoANz891PNJ7kUxiWMBWM
mnSjd5iBmJvWxTAJ4Q25R6Pb4y5rAqYZvQIHsm+Vu8va0hoErSlJVdJ3jwFyH0/M
j6Os38lR2wamE8Io0PiibrcVToK0ouWCsoP5zfrSYNEoHzU3qwCg5P1e2g48sIAV
OgwHlXtk6bPc8/TaCpDWh47fcUuybCz2zQW5NlSwp5olBiBgnrzY3vzu3rNbXgGG
DIjKcE04AqITcWBwiFVD2gH2WRU579jiVR4MSc5vIi7pJwi0aqBzWmPSvXXYfGcq
iuMfvOBN0VFQAGqqdIP5YHlnl00pyLkovQ/le/dDvQ/VMxbOoOgae6lL+g+6RJyg
TFhWi2CNV0QXqgrd3E8HSpB+5P44FBihFPrIfsmvXAESAM4h6AZJyWxMcSufknjq
cANqV4niK1SUhZJW+jvQQV2ojdFFEmEdS7b/En2YEctzz3+lmMSp8hik9OnKYKQi
Fb82ccLFSfV6RmgWzkZ1u0VvlfG4+zIW3nNT0e8Q9XgZVdbUf6uiDa4G0l6LZV46
F0YSCdqcxBDmKw60pqE0LS2qFAaoxGsHgJXWt06HzPzaPkUEt+vSQ2Jq8UYPWQp5
5E/dV1M//0v/54tb9o+hMi4Pe7pmp4PULFDP1GW9AWnp0e+HyPLBHOm5H7QCxI5K
/vduoIoK9mEiC6lL7Lrz+daexi2QzfIdi0r+krclfY6XfVnwh+b7/Am+rXOeK8gP
Q809OfCG/JiA5mcWwpWb/VdtSkYLzJoI1nSSF1MGrqR5rpkMFtaptEdLVta+F6Nv
A/0tHjB6MAAabh3UVVEG+UnpUULrtSgcX7bVIAa9cLbiWZIcd2iWI1pY/3nzNrBW
oCkslITuQfo6ifyqGBL6HGClHDajGLRCX0R1xpJdc/BuR8Yl4f4b1uzTOqInTRNw
nUnAMWacL5i7pAEBLBHEb43nxIkPh51JvIpeyVzdaI5OEYxm1S+2oHY5454ysc2z
kmVbIbtqnPPGJUTP064PELAC008mYrrMdLh613ItoMKBzvk2lNunRC76H7/aWGKV
/jw8b4Ohcj5Abl1KrJDsofCXLCghzKuq6fF46ANpOH10BvYvmNeN5qkwquxX/cAB
3rFdWGheBxo0zcg2W3uPofELskuzST/oRM8kmDAr/stfgVd9M6AmJZ8akNFU6wUa
OQiNn6PVoImBI9TE0SVLioX+xjXJdWrdSsoAZqSC8vUh20HFYefKbPa4ZgNATsmB
P3xA1jjjk3pX06Buzc9gE7if+h00hOBmfytP6WdB+Km3CganO0QX8eMaE57kXCM2
xl2JtnZI+LVOXM6lLuvpHiBVN8Bfz60OdKUKCLqhof1j8vy6hhY1SlO/YHzpLhFH
W8qNn6LhI/modEC6pUUpNtni7uKR0Yq8RApsoxALZczDKJv2WvCbKCR04q0yEerS
J9skelILnGzv9fmvJ0zqHVt0+tZBggstzeo6/03Gx1Y8BAA66ufAFvGVmk4vPc+W
phX4igLyjTxZ/AI8aZWeejZ3itbyHZS7/ZqaWEvVnoMDLH+JrQ7Rgj6awbny6nuX
Rzz9UFxTyOZIESMat4KwHFDbmojH3SueHvU9Ucf8eU46XPGzeeGzn3qshm+O4DzV
U5xVMKfRpFI1I+BJEaVF08vcBmp6iql2NEWW/27auEPGI7txc6M5Waa04Mjt/UKJ
31SxhwWaZKS+W7iztzKMiBDuMYosLwLFcXX6kL62u0PKLgVfNa+Dr4gDuE/gzyEN
3Q+2uED8/hmsIj6gu9m9hpnX7H/KtNH4dr9d3UDZO2+4fOby/WGqTJUdx9KLnv9n
DknOdJEOOYNPadyETPmRvUAHqVoKey5pqvgf2TxwFf+UKU3nnAEqaYKAT4w1iFhb
GyocNSb7NhXPU7XUPbZb4irGwzpCen+KYnxaNaTgggzR5pdD4Feg14bh74Uuz/5q
g9sWebsSat8+fhoMntpXL4uAZjxWUsIckPDDVCpKueggKNGBCqCtirjM0Ba6dEFj
mfplKn/9JK4G4ZxG5eCcNp66RBaZeZQO1XXvnVnzlbZxTHfy1eU0CVtXO8bG1Qol
ZdXCQgETCX+p9TDsIbAE8MKFVUKo/P2BrdeugeSkrFRYREPji2YbBr5X7YcUQoYU
+KXymhbZ/mQWVUhz7IXAz88/gjFWSw0Jkq99m9UbwGeCsGB3Vsk3+CD5En22ayYE
uFxcW7eHZAQr2OgxpQT7Mfy8zL+QuMxWgvtdeg2m1cU3pMbOmiwf6YXe6EHBYq2x
bYxQEsjI2jjsSMFXAG/393pCPtJ7s1sb40BrtlDfuasttGITT3Amb5EBP8MXxjWH
wO3Bus/1tXBNsK2x0XPUBUS02bVanfnejKC+k4BPt2fawCltrChdTo2MkFYZm7/b
fkHiB3ByIzr9/qaozdG66rnHntb/q6i5/136wFP0hFSYovy4TKE8Le2383+ovNLK
+2vqiyBck/Bbf4tJCPPr9QDYcjMViTpq3oCRcCCds2mqJTp6omYtlAh6c65Hmbcx
ibijZNRhe48CE5faS4ycIrhEDi+aTgr0OJg9WQhUi5BIYWHviueu48eFjRSQipxu
OKNdA5j/I0tgWU+/zBYeUdMJpYIiX7AMwuEivjD94RFe+lgXMA0G/O6UEM16pDUX
kz8/DVz7hOUTLGSU0WKNjxSLhEImDwXeaVScgGKWcoXbtM40Pky6fuzCwurLerHL
Hc9tEixz2kIBMwK9tFM/F0elmv9wcoOA5BxZ7iQI3I5+4HcCB7ZeHxHZ6SmVki5U
QI1W4zCc61qWKDm1Ygd+VOm9X7QEIR60PTV/x773eKDhamxEqsviUTcaiUHbKV4u
wwIYa+afbNHOPnLPujRoW2mRFfGVHKdnHoSTEamDHCtGna/wQNMFcY+X89scCdBQ
lKagZ7CENyzu53AqNgYUuxTkRVjApcVolgySekt34vJin0BtVnqIqAMZie7Q7hmu
oOSasxhdutLVNm1ZIVsuF8n1lUKkbul1zTWcl8yZMF7gfeOUJxg2/JKOMtDHIJ8+
SsDsBvgP44UvLQEFLuOGXX0pfAX9YON8v1Fs1lF8KG7H/u9HRkL9aE/zu6FhZiW3
7WnR+HhS6QtRsh0eKYq8TtzlUKliBZpNys/XnT+FtQnEpyKAyS/B7tos67Kd3q3Y
ZFqHdnbwjHk0wb+XlE3KXdQ5lFPsw2SFNOA2h3jHj13XIQ/N3gGPSu1FxPH4mIRa
6Z5WS26uiLo5NTEHZoHQPtCPtvxrmKgDE08z2QaXDa23KgoDAQ5F1VVbUmIo2B7C
dCSw6cJ3l6KmxRWqLGdNAPK2/YCO8DI/pZ7e682QQ7wcz/EWPxIg/o2zuOYLWfuN
vC0U4lp274btoYQrsn7152BkUL6BRCVcOKYN7IGOosVx0/xDfkMr4qM/khWm1wmB
9zUOflg0ZyM9d8qJZiFOviJzF/mowf7oGtWWfQA3HrKY9KWMOCDKDiL4QIL0gW0E
tid1GFHA1pk6iYe4ln05FvZdVYLKcXetIVrUa1NmS4/Dsj2RRPGddSm/aMdCOfvQ
dM0rVdW0RZ3j9qf084dSirduDT1O7WStTBNCzjSkBwHjWQcvtmlcglu5LxytoU2m
amT072lEiN6FksHBvJ+GlKEataYMKkJBPeHcYBZv/MQiCZIAbvi1RJs7hcQHh+fP
V5Zu+9PK0ynN7GkvZ8wTyjXzszh6PF0Q2a6d6wuKmWoWYI+JHUJs2z6X5xRJ7/wL
P8qZUx4oAJjL6agJHCp1EA2yINsj5JLsW+22uKBvfqeYmOcrMzU9F2Ih5sqyDJBG
VFTktjJF8r7u6Z7Bo0jVAsTEUqODCeF+cIeQd6+bQ6W0o/ZnbN7DbFbHeI5aWIbU
SW1czyjhhnaIixng6JP2ZZLVsZKqBIusaNC3AT6ox0e/93RtkvcczCcq0WBmhlQI
j0UbqrD5/oLC3pA5IJCZyxQC8SSBFqwgV9sLwoeyCdRuzujruvpOZuSeo0mFEiuw
DrCZVCz2PFYQB3S2KiCYR0HpXEMw2pgrR43/j0ZMLY4+eYRY8zj/bBg8RoiL55lT
9U77f1B+XfHzXss1Amr5Q1RtzCr1ZWlAGZB41gq8SaydO+pQbbz6mbPk39cZLTgt
SPsng5uavqA/J7kpmL7yeyLgxRacznz+xuMyniNJwQo8AVJmreh8qasufE5Rt2yE
uGO1ny5rF02cq5wlRIiNYPrl25Ozsc8dBRJY0oTPWGF/n3zG6HoooMKK68PbU/wp
sH9YZZUvh4kzvYqJcUv/kLfUSXINypYbbpV4cmpaGTL4ARAspO3L8JhSLzlXPvQm
SY+hUwCdE0cNO82bfhhjpsH+pUiXMsDLwKH57mAgbVtOZv6A9YykIUupeDlZ5OFL
8U7PwNF7z/MMxwS05lQ2UUV11sKNW/ouT35X0VPGFio9XW7Oh8dG9S10pctl2Nxn
nQggu/kNvrUAFB1lRiFtX19P1FdKvmg5Eju1Kwbc3ucFovlGLJqMGfeCS92cfdR1
dQ5U8USzUYviUL8qMg0oX/ZZf0SIJhD7jX4TmOc1OGla+yEQHgeGvxlbgm6qDIVV
h1HkaxqEj00+Hkmv9yQokKFccVAFpduQQB1FH9xULX8vgqPW84zZ5WzHg/+++hPd
f1LxtRtttn7fkhsg+p72r08VSRKsHrNTkLQDiVXFy/nmfUv9CVGHOQBVaCYUa63s
BoIyA6qfgK26qesa//S0cdxPZiXiW11x88nZZ+3n0la/zAoEAYwI4GjLsYC+MNc4
Cb92CwEB2nHpH8/uHxhkIaBnQ5msr6oJrKc4MPu1Ko7SPT50qzehe4JKmp34Reo6
42d+G86AzgUsM2AfjZCO1V8fYMH4x7KVoqebHLXmB6R+pIXaR3j+g5KZdCB3eds9
DBdp3ANZFArXTp54X9cRZM5OJAYQnjip61JO4woympmK1Tndy6dB0h7DUubebryf
DDrcbLmpSBQbEfO82oVbnWhAMvGr02T4qdCrXaaHivIejS/nq1I7uZlpDqzLmLpi
nB207SUUh45EN0CkN2CLxxQqQyhrPVATVztMIRmSyCbZJQLWU9r0eAKZ27VrJKeZ
ettxTEgxnJrh0goLBd8epieflbjUDY836ZYLinvUF2Uk25QnjSDerlznT4Z8w9Vw
L2hWHRhIRZvllMKSPMW8+lk/mSdV8X5F0jhFFTGRu/DwqpmBQ3hvD9UvnOQL7mdj
WXkuYJBHL6Acp/sxC7v6Ak0Rx6RV7UhJA1gZDpXV+DIXohhLg6CEbCfCSg5MEisY
9V0945QoeK86nkvTln1ZWlBExwqY4G49NBwiABEKd4SASkOGWKwOQmWByTxBdMo6
N2+ROOl7xwyJTIZ8vXLwfj3Xzw3UhLqa1csR/8QVW0cbpV4CZaNRsw7IIklhlBv5
1kDTUGq0oFzVD62apc26hl5XprFCYs993WNqAqmC7NHYKtoLch90HcVnw/NO/dZd
EB6DMMT4aJDZ1J5ThTtxOgy6DHqKzNtw65TrbgTYDR2TCx8o/uRZENlA82Wvs6Hv
XzIYoiLWnUnSwPO8Vq+YeknhOhDPnoh/Z7fM97e2XwN/7SdkpcVTgzjjrTsEwv2H
kmzdHL/dQCmi6/2EyhAcVVCVLH7VZe4Ydg46g2TxLsvE2IVIRdL/05I8fc3D2cBs
rhAnfAC9egHOB+J2aJjcM4VZ0tvUeh2Zf47Qh0XTh6OP50Mr8Issp3ErrlTvhFfJ
KY9tHfwZLJjhWJXo8IqOHRchXRYavwZ3VEIGI5xJ+sykhZv7WwcCKpA5RshrZz0a
P7yQ638Sx0+gxhYeVkB7UB3zNij9G0No9n3wPXKYX9yN6w16/vZ2aKSzw0XRTmf/
d+U7+c8WuNPN7zAZghVzlUEQ7eRk2QlD0PBA2hGifd/2l9FahGMzspGtMdmv4TXq
CFuLg63be/XLouK0hh8SsELk6n6Q76fsQlUWdgJX1AChDHp5bsy6Gf45QR5eurBv
lHYjxWlFJ7SQVsrVi9eoON2x28aA3/vjesxlRFwO/BTiuyf6RwP45wbNyGUmAJSK
ewK3ycNGfM0adO2KIiZH+78ei/zdda0AFR7NYXDOJZh4ef1cltz8uOEgSYiwqkW1
vDYYBThuwqCCRm3ORUUv5ycIKOBMZiBpl37jwgI4VlfY744vFIMpVgFKLV7YBVNE
PXA4SH4Xrwz2eSCgE6gvaXKEMHKqgR1wnbyJ4CR42Qa8mBD3WvkdbSK0rSiftDzp
wZUhmlYuvehhjrn40/3/PM6IC8p4V4LNCmR1ORekUrCOB8q3uluPW/GiQozv2Um0
06YoDdbvvbjqhouSve0CF7icddqgRlY9ZI4llXgYZ/fBRFutYeOVjOOWEp9WFKOu
aMSHbO2JHMMoByzcfTDpBpuTJqIrQZTJeWRkMtblwRKxRDegTreR9qgHMSkuKKGK
Xuovbiz2Qanr7R/lHIMYOlrKV0h7Bcd1eCXElKU676ovGYjZ97OitMGEl+Q+baCH
IGOT8fhjWR0rPisg1xiF6/g5FOvoFP//LUFJ6yrSEKRPlBzZyw1gga5LJuUDMs71
et56Zf0riGvlNZYIf7tJygr5M1ehIjoEoO/wYu8JOFT+YNujfCnulY1+ojeFkUA+
eoLEMhjxae0YDVRe/Ai/aDEWV4BYiwFKzu6JVODoH6rPGCNNhWFHXYUhSXcvtpSr
o8QU+n9pd0jCcEoGF2xoaaxlLq9TwlckQe+Lvhnf2/Fn+GlMAS6tDq1OOI0ffWX/
NuXVVHj2w6jQd+muoS+217l3H8+hAYPsIYQvzbYp3L6TWN2TUG5F1z63jR+sLJK3
IWXhZxc8Ypiz09nMy3V5qEd2Vpitp5Hqub8w9kfG3vSyWoj58mRCLdpuiVs5+YOk
t5+OuyZWDWNTJCP3oxlEYfVmqb2uDSoUTxgSYntP2UowTjrqbIumLAzzgEExxN9h
TaHnjqF05ZqbQFt2Fmwd3rQ3cUX3+KfXsZU4/K+eQDs+rfYYeNk94Cwg7sCHUlR7
EVBN2mYd+8NtNl/iLx80/li/2PYT8FW709hdX75DDDlIx5O65G1jVEPloCRrAs8L
aqbtV06mGdjJmtktiSuiXr3fCk5h3xoI8ejoO0ZHXooig2D9w/Se8QaxRrD0hM5A
DulNG/BDfvN621lcECrwooSbMlZJ1GsGDnNTwuDE/tBeAB2Pw9TmtYtq93pDWMvj
DDHgmvx/yxeZky/KbErJMpwSRJuqhyc3qYL2GgRpHZqSgKUAgn/hJ955qLMVvfz+
DRiMBirVnoLOz0UpHNrDIscc2pdAkAghDXyjzndu+Lt4fVFppvyzNw+uQ0tMkfXM
tAfbz9eTsWyABmo3r/H9nCi6lKJV2xwV5fU3ElAUek7cdsWDIuAiQUKV4yf8ZeFf
na849MVyVzhjew8JIQSz6VT+z8v+pJ6+wZ/a0eWS4kYOyQeDWRAw7hBo2Fixl5mB
BtMD+Go3ERlaEb62ynR2/HRRVueAOvv/Sue16iZBvQh+xBIB/rpFqZK1IleIpgb7
8r7Xs5VF4E+w1j1LQYHl4vA2R6P8+ha4QaAoJCUggBkoPs3may36qwBAEsfK5+O+
HvqosBtQ0iLOslBx4FOkN6zbbPadGQjwfVfwAKPQlEvZkLdxnWBMfRwqKcxKfMTC
0BgkJvHRXTmo2vxVdBJjBIHAOpCnKWydopRZO0tNNQism2QKCJbDvqZVfKgxJSbq
ehv1i65NLdhUuaFzv/6Vr/EgUP1yrCEOyo7EROWS50FeAke/qfeBqCjXp6pe3Deu
OucTtRoVT0m6pv6tnDhuRVEZXjgmLkBud+qOFOXGYNBqYu0WIVOQlhfUyXVQpHZc
q1FSEW0rdEg4RvTbRWjo80Kybqat/bi5pYw/6tn+I0BFhXGuWRMwddKn1ybm5i3l
S5OT2Pvby35rTHtz9DIpMlq9UkUFnIfdmc8sC5jDVoKPIx4fQERRFyPPgUtR6d13
KQWINLjqCuM7JiFvFBsEUQX/+qilXILIthm8BIqJ2AQ+7vNjki/437uDyeHj0pjG
49q1ddMs9XoJmes2Y912LaWKXwUi8fEaNQPeouBfQ6aCTtPml23noJyPzQlCZIdq
2NSIfusVGnytNLZCTScSWBaL+1xydgCOj3fx+yb3a+44hR/dgwH+ZqkbuhfFFWhy
XDtjSzNAuD+6JBqTM3tTvHafNMy43BYtAo4Bf0aGvcBkOguSv6Z78CK0hBqPh/ht
lQCc3sVAlt7t4NPT1He2EumItCQo+ncNnaqxA20UvWbpqEKZamyJeJvDBrjQ5QM+
dTMGFs00GF0yXuebYl8Q2H+/crBRS67DmUnDxlG43hUA06eBt0pBUtVcVrzzV4R2
36vkY8OlFkYH6sF1exBEU+nQeVIy16A5WvP4HdzUGx44FV+E7NIEn5NQFeHp9K2b
uIwyn8qI3W5oDoZG+YMj9QMgm2SpTFtObtD7czTdmL3SfY/Un9w/r6bFh1dca+0J
/flyyE8Eyh7+A8SRR0yeV7q1gfyNJCQOO6KDmw6KzIT+sb8jQ+6qhFN0Azc2d4rW
kZ+RwgekFjXnIoIa9AlN5G82xnJlkSgBLtEHSlC9RdnRGpMBO6oQdhfH2OiV+7vi
4yJjEusaW4Y/NDmpkDh9D0ftCUN7I+ijHTaWoBoKDh3zsWR0+QEFUnRTiIr3SMiN
0IjA14SlHMRKQjYXLbMAJPhaprvyzwJ6B8cdkIPno35IZbZCM5omNQBcUdW8aBTH
njXDVTJwa726dzg9WcYEtAVwLMvw89EeweBLAYVFa4NSHzt/5fva6Qo2Apov5EIK
q4U0CHEc0sE6YdWqKniwfj77qkX7hdy4+LQeai6Q2M+MXmay7vb1oq1dzGswd6lj
neq/jFWBxWWrmF9Q1wldZZ0qSdt+7KzFCXZTBaNiaIrsLPqZn9cfLUHyIEoLIdbC
07oGaihthShLGGruByMUK6/pcK/I0UjnSCmhQh92PdyteELeyTLKXgBPUD2AbxQh
DxIEkP7+UX260MYXoLpfgfBiGUJtZ5ExOnsjog10j9hGSwiJt7y3wuAHiApMYSnc
Up0JGbJXennhXopBw5x+58ppzWzlX7und2FjYq31Rz9Td/jVrjU+yNmVU3zFB38t
4r4D8zy8Uit+MJ2uM7tE3b0yCQYt8PpcPjcyULtlDl70WHNtR7Jdwx94fxuVEm6s
4xzOtysr6qj13IcvVlwMW0OJqezGXU0gFFyeP3KeIVoUcnFZRG+VgBkNQPM87PwK
CIaEZ8lYVD7SPuVm2Zzqy2iFyQjfDn/t2Vcd5s+F4t0cDSjEdaOHpZZh0EtqZlnJ
Tq97ExGpswsJ2SFUtIGYO+XwrQFNOmsMRQTURYgOLZTUVEGMNRQXfQiERsYki9Ku
RvVvZ+l5A/BZfn4M7x7p7Hs70O1dbJtTeGvEmu74+tOPNdxbAglZCBuMDyNTgq/c
SOLibwUvC76qzE8iZGyIPFHGm9f3RLycsNAuBkFZNFNDfAeA9d28r4VRhkICzTJ+
45Qhihx/urSxWO15mJy+763rCSu6CUg0InwFa99lIyRLl+87JkfoViCglHftrpbq
WP+yPdct8SH9EyfLvBCtBdcAeZhRkpCexfDmKnFKxOnEGDgBAKJIkyJWepH54bI6
4vkUP8zFBA9hBrySfPgx8wfRdLh7WI0nOgTQ+JZtUJBos8zUp3865QNdZZypQ7l7
F749qo27pA32bIAzb+JshSROOlK2LpsdrpIzVb3r6FXS3CY7LkvMtU8nUVsLrTHu
Qhh80MoMoZIWo+jMhHDyp/uDhDXt0t7+M7/4SDDEwlWhyOe/6ZzL+zPnQ8d2+eJR
CCsSmJK5zaisdiTmrPGcFaAz1DTJs7Mzou1koht0VIn9TO151P0v7BfEkcyGX9QK
JqrbEZ5cdHajs3z8BdckG9br7Af99hCO8GeqlN5BlSh4z/rdJRP4MYSY+/QsrQ8x
UFjcuGcO34roV+l57PFbNuVUd7FMdtKmj7AcxsYiqezOQh+UeeZhylE19hNX0nA2
9CwlnJxUQGPa4hYkSze8B0yUlaTmp1U0o+W8Wwv/zTijNQnweFOdLWTYMzbEA7Kb
tI9QLLEZuTxarC4vNNV9h6/xZjh86abSzlZYKgWcZXek7Z8pWhHuPeiqySb0W/Gz
Xgn+hIXkVHqYaOdiUBLs/SjTNHaMvz/wSeSSd6H+cDfH23wyVqaKkqaRukNxJOTK
jzmuCXy6WGx8lcFFSdFCullldMiKB0ILsQ4tYuNaDCsRgNmeG6ia/crC21lk/e1S
h6kWo8YaZxrONhPNjoSZeiq3I2ZnJb3miVJafGXvjv/Q4fTOH0dXwtEwzzjjwCvg
ai0kduNlnVlK95e419TnVSYQh+YCnNHUr6ezsI2TcVDH6pHMLM7PeR+zXMuXST8S
ZDFmL/iddY1CuualRKd0kIqSG9IzNy5WAPEkNjJeYi9g3L/t1zy60xVeYtI4SUxU
MXyS8JNZf0e4rl9N+y+Q9l95b9UhavXaYtsmFLcMMrOkZ3i7YKrYl9xmh0YOudyU
dFRExZNjwDKNy+TrjtWNsP4ehQ++6sqQnUP55DREdqtGpcijdy9y0xsQRw4VwBf9
etzXcesrsE2lPsLGcf+3VbudQ9hE+hMNjK9EUDez0TZKfZtJ7TtOUEZtCejQWTKK
4GsBiLa2aifKPQsArwWjUEq+pPrSeCQ0uV5cULdjm6Zad35Qk6Pc73Of9GmdIs3j
5eXVOAtsCpxJTJ6hHmd077XYtUBjQP7RWIG+7JMwWL6YQjPw6g2SMj8IeURWRCAh
wifDKx0KJXhzJPCBm03l2LRscIPvY0xPY/L148h4LBPefwk/6QhmkPpRa8hEwLRa
oIjeQ+MUH1hJyoNMjFWHKfdLHpLLWgRD0rRr5yKYQqNx3HgQSdotgIMLx2lkc3Rp
qYdZ3Krh1339qkZ4LiOIvAjnn19Ii0H38jN8fDQ0i3cffYHAgivfW26SxNlQ7R5u
5GSiPs6FbiY4VHLRdC/25rTqt9d3Gn5I08xQaXrir+6zCQ2PB3MrsqKHK+ujb2qN
pO0UNyucmlmvx3c5XCam0lAo9Ys1zSDErT7PnV5MAB4laptREPfTb1aYWQV5X0+2
UAa2nltn/s7l4jvMaupBbKRXOoDIocGfve2doNgsQv44Xs2QPVA87T0Dk6gJd60L
tIJ7HZZai/gbquv7JDvRjsuunksW81CuVRVNFqK9IgDwFV4t8mDBKMI2rhzlAGNb
SnYFybhdt8dd3T2Z5r4C2joFtIRTqdkAO2SElOZkUSeB4uIe5TkBsia5rvWiAvCu
51bdZnrsRpQU6lUH9UaRu/Dwql453rorntHVziwH6qpbTiXVPwvBbUBzrb/wYffe
uKmAn41kwbX70vEjIkEJjs1k1+3Aisg6oOcXRnH0l/sVn0/l/7LS55A/79+BLauB
Q0gALW+re/Tpr/myI4ROWBsZ8rZ8LJJ6/txXFZZIDMRHp5K3t2yYjofKd1APVRdU
58jpfyCY9hb2v3fQw5XWU/H5aNztxBkoU3zWaqV797g9lR6Y6Di8+Wl5YU7KP8Vh
iGTKx5fCiRxNDRlSk8nyOha28UuJds/JzFn7a4hSVlCp77iHSPrECS90Gk8W1rgm
xi2tq1hdEp1ZR8RtXyV8I19Asmm7I2bqAQD/OAh7BV/nUeSDLC4ApTR1jofykEPq
Ak+hMYEcdASYGio1DxHP6DG8kZwype6GhChBGOSFDm7nwFGiyy+XBQ+JjCHuEkKu
SAd2ba68j7oSOqbowy71Hkk9iciDjPgCacdB7aW5aioVP6FamAPoteAMC/mGm0d6
tp0yLPSvBcdYSgpGdz6Sx9fSrx0Zk6/OvzgJKvMX3NGFnQJlXMmmZCTj+hQPMd/t
uy/mLUjd5RqW9R2okUtirZLGF6H3xutT9oMuYLheBm79yMES0UqgRjJo5LQMlaV+
lbrdlKYmVitUHoTJJZnH2OGks78fbCFtVvDl21Nv8ZrMDjUjkaRE2K1Ll1DSN6Xx
u8P/lz1F6ehKdNDziyEehoE12xMw1tTJqtKh0IB37DqGC26+Um/NibXvGXzvfeOl
ZyZTLmjJut521VUrBWHwN7w1wbxxN+vG5O2uzXXiEKdr7TSG/1Vny0MUt+/TxuLS
4Ax7Vo8ssdhVqF2+jw3MW+QfH1VH1zedHb+9vuJLN/gVW6ChBteciWTH1WyfBjZC
pCcxlEwi8X3FqAhgA80d0UQ0LtpQmnEashweNjOYohqsKZWs+sjeZbH113JFfrtJ
ZW5QgIBPrF3H0rQbpJHtQgjO+W14pasUaGWs3flHkLChBWAHm/5WrffqAz3r8+4y
B4LxyiALFz6LP7XdSieRS9Q3c7nTzrYMAIxxVw13xZSAE1btoAi/q91tVxI2qD4W
0E6iUhVd8yTmlHR7gdUAW8z6qaVSkEIanbj9fSxIjFu9+pAszET/mkSUEltz5xSj
BLZSt1HXLggsg+2RtMZYRb2zXBgnkcGIn3EJAY4lZLdDBVtRKzeGKXP77M57RZ1f
PHQ0HFQsH1J3U/KDsMnsFDqKJd0f3T4U+3XiGSVuvSc5w5dJeAGwg6CZ41uBts1H
kzIRukG8/boFv6qwwcMPKWeIs1iR6IlNGFPAYB2/DKIIMDfVT+yBCMI5qA5RGOxX
fVdlDPfWE057ttQmJWFIAR5PpuMORw1Yo0rqpjOQ7oyEUEnDuUCm5FjVEA027/wS
EAcziFBjOTwFZxAkNjrEjjUpgN6mbPZsHntyCcXmiwn+wGDTU91oLX795wDAp91q
X7KVYxgumL6qnCcbATEkrrI74NpZYDpWeALnILwuE7nrKHG1JIJ+hA+pQX9OUQft
EnsaN9HxVDLAxmkSyuPzTdsIaPt94Vo/esQWwMWksE5+XvDxGZEoLBum21sGBhrQ
kZHQFwYPreHkpu3/Pqc6gp00Sr+ug6zUTo+CYaRdP7VfSB9d34NGsRYxK72riLAW
iwKRsRILh1WmFYt4sey6WmXWzNQy5L9VzSMHwTICR8M09aSRgp2PNmZWMy1t6lWq
DqNx6n1v8xWCtpAntiv4v8SYkjbzeQIXEXw3XqIWaTc/euz+h/ikp/BN7kwMLlZ7
buTky18za5msHxlSii69tuMWsjbSPCYdlZNbvQXNvpKjKqMoFsw822UnIJcK89uG
QM/JL2VttIzR8cDQSJHoh+f+vK7OjEbZm6MJwd4hsPWbvtYDodyE84bBGAYJigRx
1mxF0+E6pvYNxkZblcvZI3RgYP1QKAYczyw1vGxpczvPGfjT1hNuuDlJTjLFTF9K
vDTdz0+zxsIGt0nCqkVfvvElJ9Nv145TCibza1r3WVNme3kkhu4RQUO/Jl24KWqa
ssQh0/JQNXbhVxz3d203f1wYzQtJ7ClIqQrqbmTenDkqtmWBFMQ8UrY+9qrR6ta3
Rx6ZUnSvc7fhwWLfukNW4tFWBbihE+VbHWQ+JW0W0n64VJW9FttxqajJHRL6TFfo
/lao02NDgL7L/zvdScF5wm9mLvyHdAStdBep1IJSNcP8foYVmRSqaO1mOm98/swD
is3wjwHdQCM7YtV5T8L/5L29Q3j4hCEzQBrQKNxP4W7RrA/DLkB3USKMwBALm25O
wVNsX3Kwa5HZzjB0uf4rAsA7l44WqdZCnQxYM4Xbdjo/9h46Dkjd7/k5fnkOCEbd
8FCMxjTy20aAiGt7fdS46+i0fupvOsX1wS2hNud+2kIEjecf5da/7cAKG/V8En2s
s/PpGZY7aGJPkASoU6qC4mjqU5/mT7SbhXPnBJNsudVdBeO9soF3gAT4w8hpLV9E
+JnI0kc30UKjixffkxftnHXo0myQD3RPrkyZh2m8kH6jMpW1KMHJ2d7MCLAgga9S
Rd1Wx8NRvHic/anfCnKEIUBQ7gu6oZaZzYHVsamg2OtRpOdOb1Rv+qoAZFLAqZff
RMbe7pOWVvoZMErRbGH/lKfWRxHCayefx81Vn5SDggQfxMYJjz4fKKSjJ26D1yh4
2LTkznyCwkUrspNNJCvI1Ua6NkJYRthPwhwpsy0b0KlqPe6JbrM4yzKcGdXhYmB4
t8RVqekbfPrWFkJYhlhDByJ1pj+QUsTConar04NdwsSfns4ldqXRdzNnpZEnvTUc
F3C/gecY4AD85DUIvZRlLwLXyrVCCqzZg7cWSDfd/a5DNfkShYQ6aCAfm4a0iUDV
4/6vXcujsVtuOHr+hJJu/YMYye88E8tTOsKwPO+HQS1wDnze4KWAT+LFwdfquRVt
hDjViihlCN8jw5qM+RXB1ZucaasVXuY4Sc4oyyDeRtz1Rt9+D/6qn/VyqgRAlQzx
ZstlL4yDZolRWEELPvtkaM0F3DKW2lJ0A30x0ASnInyd4IFZcAOEHxbAWbSgD1N9
nCSn2OmZiXFLAaaXcVSweAPvmWWTut8+UbHgnvtmfNGe8ZfVdwTDAdO6MZr0IJDQ
NT2gR3G/IJIgvhxyHkQi7uV5ahgr9W+ynesQLVhxbrbQmgKzFJkAwd//gTRdmZf5
BVMTH5DsFfbf/FjI4wdwhlodUQbbcVmnQdRxnWykX80f+J/jN1VQpesrdivxErfS
O5e1rWPxfQ5ydTLKIIS/xUa0ULCf2RRCsReSY/87qxAzYBUcVMykT0IoKZp8YY09
VKVHPhSmjILoomxVPVWF136XxWvSmUvBhy/J2Vh956qpkH25vqJvXqZDYT1Id4+N
gC0ygMR4FR8RYrl/fDNIKlUk3ynPsnL5h7X/AGV4gO+8okl70Wj9MUcbaxQygWVg
SzZKUD4xG/b1r5XB0iKTYgIzo0gZ4XVhd6jl5wtq+CUlV+gxh4RfhPmYVZRORKnx
fw2Rnm0dmKDMPbUZMpDpQJF567ZBTLlhhJX4fL6uMhnT5HY/nPMGFThd5IKFVj86
53JYr+29pMQH82SjF37X9JAf7He2XxVCyKNAQR42ARulzc8hy63N1neVIkFBFXZp
aCIEihpLm45/vsxP6u5o0UjHL0K81zmOZ306zqODY52i6t4vraZBYtC/9W+UhoZc
pvAwUxX7T7xkXLQcruYZyGuvc636c7zuGNgguIzCxMgZFBQAWnSAPkRa2nsL8Pmm
1uW2t0MO7LMFPncai6QbkUuhuM6lD33uKCMUc2mOekYTR5zVXP15z1KT5DyXtSqN
0iUO4QldKWQqMFH6KxbbYR3oyJX5cXp9NaP7P8eNSMtgWwxh+JLb90/ilOC5eAUw
udXAmnKnWWY+0bNMQmVeQpE6vLQH1LXVXVKu2EbSQNkrBBzPUJjLq6dfACdLZ422
nfL8wxMbqKAeeI6OQ9DC8uO6iuZdaMJEMf/w/98qwoly1bJ6FjBEd9dgH7ViXhYZ
Y8jR478r94on8Ne418p9Xz71mx+wJb9zLPneWDHvK1GqE5HD95bpGcrCD2nl36Re
zvDnq+A7bhCgQXgg9tTqNNT7GpN8UH4Cj8jkx/lAiFO9Llp3pS/7xLdfJqP7DAEp
yW4QLzkG5uHFOxM9lcOeKd1axLYX7UDYIbzy3DO+P9v7hBrSeP3kObpNKvN3SwS4
b269Hpury74LtUYq7ffLshH/t13GXNdTm+3lyUghwSN/Px4BBxjZ9cQPjz19+IwX
DCK3DfwcASIlsv8wM+aJP/ZaMOG35PmyBpnouq0np6vNrrAx38nlWKqVNxrAc6GL
Yfszb0oJjfJ+58fGLU1PCYyB33ppRI7WMOesm4nuADKApdMtIopydSmBP6wKXUs+
myO7GN6lIr4QffuywHzi4+Hm5sz3YgCztvfwIuXDyRTl6WfbGJGOdoo0t2ZmMATH
rQN8TpC5L3VmN4roQYS95eHxOmJ7VozrOL9PvthbGDJGFsWqBLDq3W8vm0eitaVd
RBTgLeO7jy9A4PprMA0hlYVXd7+p/Y31Cp/kk0nIUnntQ1+UpgAgSnjhZObDvZRm
PfICVRulcQIG+XZxBGJGDa8S1kROkGc49Rfyj+t/tYz8KWgpRBcZOYJLjaHGzTHi
ompPC7BDfhoRr+spglnpEM7WqTG5iijNe4tlsKZJDyzuOwW9AO04gSf+DwzIGNDt
SZSoOeAKTKUwMcC2mv7m8EcGCUcVDuVAGzZWfULzEOvUdL/uRyq1Cp/6R4WxsKb4
AMvxl8OL0Cozj0ws1l1mDC5ruFF/09N/S5EaHyd5aRS4WlkgiSnHswMaodMRgoAe
q2pYHn1ZsDY+xDSeF+OXyH/DqpfoYBVD7tvv/XNphT9LQRhuEnPhne4ZELFYODOd
zhnVqRMSyX5mQqJEjB9ocyN2zitcFrf4jIuqCRAYXetJm9kUteG5KfPaDKpcZYBq
pUgxIWiYiWUbvtwKv+6GGaALdaEsxMoWuBU9lQLI3/1oh1vmloA/aAaBDzSDyJ18
50uCVyEeURCS8F7Qv6cUoVOThE/2tQGkIhXFNZDuIlgjtCSk+wOrYrE8A6thOTBb
1mmLb6KFnmPzuZuT1v/eWCeY/mHf30U2qTizNcQhJL2Y1sjwdzEe6wkmWvGlOEco
ygIoqJ1Tah7X9S4C3ak4acIi7l+QYn9/kjk7N0QPDo0fDUL94zFqSvXvd7x7/7ap
UiB+OsbuVyER9aMjxk9lPIzRvzySyENowYYwyy7mpz33Z5/+04gDpw1h+fdQJPHU
B0ImWm/bLHcuEPTxml7zPA5HeCVPaVjNOKNxpxsIWmnfQfbJUDWPdGRUIkSkUucI
CoCcOhspCjjPhqsOe0EeMA1uVgSmeRcu/Hyl/TZ0jG6C9Yx2NNX4bn7yS+oNZx6v
vrrhVthRY156gbSp+pjH50RODLzEL4i4WE0Zss+carnQxzbXUNf/S7qtjlq7YDQr
zcNyxRItTQdPdJx70lIe0BzPnI+6RZZqQTxFsX4a9lmWOtxEgITCKexWcsYYVcsi
6R8griXv17Rwi2IEY3Qo6XmTKtrvONH+OHmIaCDJyMCsBWf3Lm8Dn4SiuntPNLSV
4ITpzsrE22qNn+3U/SE4xw3aDMGRxzDLYs1jGf/zWtMJWcz07KrYD5w0aPA2vVTY
xpKrWDXn7gUkB9AHvY7QbFMhDfhsqwAB6u+jJi8ekQoFTgA20J10FrT3jkJV6tEd
o6RY6j3D4iA6Z5gwZhuX7LxHwuUsqdEPoJw5uEaorkJT3EA7GjN/qWoP8DiptPgP
Ifd+1nXevsh01wjH7XpVAlOdmvMXhtywThVo9NRwRxeN6kBR/m/v5Y712fZnCxoM
cL76s2ON0lnxs10CEiyamlqzTTtLxKa9JVfJGQzmE9DIBrs4aaue3Sd+1wasMBMb
v0qwRTGyNHFQMsKqa1swmP7wMhatmBPjeZDovjOPpA+JOp5V7AM4/PiXpxE6hDK5
hPS50s5bEY5lclhcVULCjVdi3oA/toOlW/RAZcX+0hWPcAXL0qtm5EPguw50oyDc
a/pAi29qHVSlNpg3YKgiQG6YZfMBENRPsrMKmLg7brgH603mfpVDpW4+DsDxWM5h
N9Z64ZQ5eD49X240sWKeW9AR3gMMljvfzan9WauJFi3RZvLV95sdtA90L6OuuZ3f
gWR5k4p4uuYc3bMpoDevQ/phpGTCwYIp5bYv6AacUsq0/M0WWAcbIWNb4tX28WzF
+Wk6GLXYadUxKRFfjtriXZwrILjYemyahCn5/Pc1UeriSvaWSXBVhVehwielIjIm
uQ4huj8uteU6i7Sq3LDyiOuryb1LGm+3zKNSYIduRiFrT23VOgM9Bn+buHv/3bh2
fnE0CQDfbbsL5/VxmE0raOVsnmpaeofQzle6Cgde5cRLclH/43iihjanZkL7wsv2
c9y8/45CwJTL+IiPbARS7whDy3IGLZHQGIce6evxWN56yW6yMxu8bgFkJ8KlqDvy
oHruxQd/wz0317N3IzDjvDLA7Iluye+HB7AH0HPmc/fPRjkRIOQdmVYL3Do+Xdvh
aNThua92yw/3ws0ifAQTE4mL/GNJe02gL2qRj0kB8RBanDTsLRe8zKA8aGDrUr7I
HEeWLJdk7BAlzNr+vEmB33SjEr7zV2HQpn84lcUEfIwkhDzdrVeYHhNV+HQ3ugv6
IP2zQMV2fTmkSspDCfpb+cP1wiReSaftGu2sDR0Tc23QR6F0fWp6QwmFFp6eNkY9
4x+ovGvbL1mbym2sSV7ifZ99n0DT/Vip2gFlP+xjsdSEzqoXPmtoAig8jTc27fCo
qCwBrMqUdfXaRCqS352ejFBWBDM8NkY5zt/AMElaY9kr+dyggswE7ZrPNDRxZYhZ
LHhxCScUFboipX2KUj4wdZB4p+x/9yH9C0bnOxolDHMDDlVBEp12pwp+Dfhe3i2R
ZwVvHeLg2WGv4GnzddWI7X4ZQRYUeX0lrdh4KF/BiZtwLsvxn82Zufjg5uQUxBHd
MvuBORFnTMmyyPzUGylWKAm2vGIw8wx1NysOaONDaw53/DR6vzWshfQnlQ7h0DzM
NtciDfnA098E81EDrtOid46GZcaUFwR+LEZYl6DXhN6AI9LGmidk3YFvpen+koPf
t700lCzGhQ9HXGuiZMBF5+x6Ju0mNc9QOjSpbwsyMyCz+BT3CKiuGqwMLR6gOfKA
t2l4G4oadELgEtFhN9aCNgXcuL0qc0RDRdOXmw+IKAhcMBstJDHi3e3dIV6/3r1n
YrgvZ+MeoBWdpY/bUSGugaQoN/NKEOfM2KION7c4rMaSsFEcUWXxPDcATMz8+67x
/7xen0UJaJgw6cIJVUhggnqfaVWGYCOOF2YTwh5z/rXrQbjaZi55cfWwLsW/zXfK
DGXDw0alJt18jjNsPMHhXRZxv8fbV9FMFiPQ5udBc56UkT/GAQciu/YUq0b+cQOz
jqVzU7gNALe8B47FhtcazSFClucQHFN27Nvf5cCoey57ksUUGbcamhSYZmw4g1/b
CvioI17I4wOpDAWc3WWifT82N1eooj2KUZg/tPXCs2tvY88BvzfRDkr0RisCKcgd
Vvlv3rthfnmG4LhHg8CGWh4Kvov7AiLPER4x13uzkiixs59CyvTZ2yt9jILXZ2PC
vI48kVO2JBwOonKDzIG0HGXmIr2hO6Rk2EzY3y3ffrq93IX811wnRZSYYJcKVDCz
rjDTwh03atjfqEvOQGkunOnWEViFo3HKnzn4ZVBpFO8k6DEifwigY8WVGBSfh+hd
O5JDbWRK2eAXvyFKwB43C/NFC66frZBfQOS2N7WHTgKhvY3zChKtvy9w15FxTZJt
mjQv99RNnw8HOaarU7WhCD05t5hxL3tUDp76kceeFfmkCr9SMo+w9hLqsqC4pny1
fs1oC4hOVHFKrmecI035kuOZQhuxiwmzru/6GGroamAkDvO1lXxrBBghmR898sdN
b+6OGfGNXmM2+/es7+eUE4w6wcOZjeV3rne4bEOjueaVDr8iseF4J/F+np2628fI
uwgen8nR/7dUFkzuR87JPdsySTZzC9umCUOYxJBtEwM4c4Y/hYp0MjvuYopslbqf
+MDE8pieUkVsjPgL4QxEmTNdF2vpIHXGM0wl2WWst4Slcq6zvwoUxYVnTSSTd3zw
2dYKyDb9kbZD9t17ZcNPsaFkbxdl4RIC5HWVxI6TAGu1cPkBWOT/Fexd4hdghs1W
df9vIE3NYqU0j0IxX0pPOocGr/kPRYq3Q3i58axjtXClFRZEeliLCIjozYVoCS53
el3cvnOqX2gNO2r+yki1VNb8JrYy8d+I4czwKKOBUppvfBGH4DGtTUaRqQXT+Dtu
piw9sKGWzuxUFXQlHgQtujRZjnUUimmXPphwNhBRWPfMchCEZFzDLwD3g/9ipWMF
mgmdPKPaUP5YI+a/sDjDKJeguUu9yXVaGCfdn0zlXi9rCAN1wHrQW1Z67E7YVbXL
I3/gJ6WUXD/wzLb7ycTHC2UiDQBm0vaDSU4e43CWWxDNnR7id1cEpdD78AOa8fUC
jJV2Jcn0gOEs5+YSsm1wzjL1U81YUOcw+azWt3jj50IX7nTsLNp5I271sprHxpSO
A1O8IwoqRFnH+s61GeHcliq4jfXRoABfqadaLQwMoRSzcp2QtDzQjpZuEjDkXvQf
VPXNv+UxpBZ/Od3p/eZgPXQ5eFzJrLUWuNy7qd/OP8rnCkAUkvqiREDeFmqB6x8h
DKPVAfVUtamxlk91wP56rPGDVI9JiGeMp9tqqwqPO88x4R/JsjSAiwg2YcRhQcae
8RXx31x7laKY3sJpwWr8D42LgtHv7jvaXwfukQrdYms+cg4C71F8UE6+B7DaEqzv
jY25nZQ2m04LD9RlVlUrUpXGNxkJIgkOi6/3IChpbaQyOdx1hH+naHQ1kTKZDYHo
Ho7qAAO5lpJtqCQ1bwu5+OGUWeD25jfiyiAxDbN8EJVC6jvY1aGoUL6IMFdBmO//
swLG7cEfKSuiFaouuTwvY26ws/rbRaud4+Eup53xiKMDOSN0ISOYMpgXi7GEFbl/
iZuBRTSrLAFk1c0NVNIFqfXsQ4qjCwV7MDvkRGAQCCGsi+0YxU0Oe9WkEtzwQi1J
katLfJjgtiLZtAByqHVL6VhH5eNDCu9oN2WhC/D18haXWLlQJhPQmZyohMUAuAJd
iKej17yqgiDhnfSalnlffeFwOQGW/VEKNwf0ouhb/aZda8mPhhfBFL/fu1JlRNy1
h7oc0njt6paV4tkPldKXrZa/7BGDeU0nCqk5lt0hr4rMUnuO0WWbrwxa9zh8C7HC
1lrwTl3ot6yRRkY/ss4d+wXUGEdtM3oT7K1RGED3bkcaJwNjDTWWVMdNo8fy6Ji+
GMRdl2sa4BkR2ccJLbtLevqqkIhTf7QcKlSQS0GCSxjq8DFTWx4tScyPiB3Sz19p
EyLg2BEoVSB9zLUGPLW2aUJx+VEXtglgF36PheQLMy+hUswKKqx1bf69bPMeDTkA
tvMADFDCD2SeoLx5JBEnu40J/4gU3Y5o6nm/JabV+JKX1b1tO3Y3q51VWUwzcS4c
4n9JzWYMEYhMZM+C1AfQ4sal+GDLL/kNHtMBtqTzjkf/qD1+exAkWITEQY8xr1Ov
b4gpAAdcLI2m2FhWfHsVDbIepkoIRC3CmQZAff2a48+9UXw4Nsvnkxh888C2neoa
bfi18oERfxkiApZvSqKSqK1tLRkRNOPef6gasr/MNAk8Bq/SYedCso7e2XVJdk3t
Uw7DmRM9ehVona8kNm7yNJwbqs4SbD1GN0A1Qn2kxJ1RTB1usGSuAWopRU7dyMW9
xDwTPD7aDU4/9SNSWe5maRS2a2ejaWvIwrnWxKi+LsXiew1ewzf8SMC8Y4rJIaS8
1iVarHmPk0vUd3bSPmMJRmthcCmYRc2m8PKL5KhEWHSJgLehg6Q9Ks0iTkMsOy43
qc/tFd+q0usMVuA/sgZqfcby9B0kKHJ7QmGmQcNj+HzyXy2G2e8QfSXcWnQrPB+0
QQWE5GTWa9EWKGZIWLLrW0QNxnzG6rFWHG5a39AV7IV5pgjwfW4KndYKDKVFRIy9
CMP80xSmBHYS7N5XXdGfdxPwa796jXBKCoSEBqOJZnmdl+96vbzAOJ1h1Tu8KRsm
uuxEWmrBJujOmNQxjzt+U3LM+E6LmNPIXsuYJDPeP8BJ2o/qJbUOnuaQT/ovESYj
ycPu+/QdZH9Q382XEYFnwyxn0CYIB8tp3cavslCVZi6Dwvj1xQWg/qGkLWtqla0g
99LSO3hbjxO7CDus/AWHSMrqlIZxUe8co5RWnYbm4uPhT16AQwIlJSBTeBPD7Jiu
msOABFkahydC7s1iYDfqWFrOhdMxrHfXzORWPWXutUAMGHbykNeAnkZ3iONzMx3H
iObgeTAEC8EHhUCOVHwdO7DAbDcFpmHGEWB/6DzgQKfoZVxJVeRu9qRVCd4GMYyu
xR1mvY0NJUwNjaX8KH7hgsMe0R231K0xQJd3hTb/8Z/bj3jcO1kTjomvk1bv4jjg
ggvAmZwOtkiXEnuDo786Nycz9mt2yeyBix3od5+qjYLIoXzyzdnBI2SXmmJUvw24
3owvxqSgoofXXDbG4KlXfIAqilgY0lgewi1mOLaV3a/q58AMzKL8qhYDGVZIr/04
sZQc8QAtJp0jRefsQBENGVZ4bkeeAG06crElfO9LBa1d1/MRZf3UsuNmcLyNhDBn
Vm/iwUZ0i6yWhBW4pdwLUBPK1zXwW29nB0RLBRvQKfC+1xhlJWRM3U+SNq2ywoww
VVjIV6ve6lb/PwY8b3KODLDa04a/aXU8Z+OPR+ytrJ2ds0+Rb70d1b0nNEBkfZQ8
nQ8Pur6Bfu4KKYc2ZZ9RkYc6f9+TYZtaYhU5nBmzie73tPxa1cSDYbo61ampM/84
PHESRRM+7ezU0yy3acEujOW1DEWb+YDu9d64HrqpMcnY3UNHLrXBYPori8W51+2l
LbsojMZen3YHvIrCp+rdM4j4uQRPxjVpK388MAAsa/u8jOSct+iRWt8s+ZgnvCwK
1iQAWE6e/C8RVZKtX72TGf7K+17XIN5f19oZQt6T9gYfBG+m0lHoQm0HbxtJDYSx
hFO0o+rPl/1MV1JX9uRfcZ+70SQsieEX2cMe/dpk0p5wIWL1JrboVTALl0KErgGW
omFom5xIzw2UW050xK4VOI74qiPolA/HIoiH/ftxIMk70+IKb8Yy3Mg6u3x1Vtqc
gBOx5SfY2XHupVR98Lvr5IXb8Xedk8ojp5ggloqnDh+j/T7AYeJbUH0rBD4wYdXk
U3VXnb57ZRukDnPtNVGmPhnyuc+qmD0pzUP4vwsfOcaZ+tAnY7fPaXpD8lcWS7vd
6g7etbLdWACgX1CCWFScvM4fITpxkPt3//yEA2uHsqp4r+9YK3ZU1ntEHgVKCZnt
T9756ymTjzIgNs9D6p/+wK9BSpUO2OOn2MRK2MLe/+dwxXFu2+c8Igk+T56i1XPz
kjLdv5izFZO0ulta28YxdSKjkdST9mXSB/UMiTSGMfXGrx0dD+XmSAp1slmyWSMf
yPcRWbqFNpEQBKw0cvLXiWnnciAN16hE3t+mNb43/pIZKotIxDAGKcaywFyc5JwY
yhzX/gOMByz4/IbXkBQWY2Zybg9Hg/Tgzgw1Ilcpk0a1KMRogo8PFcGAC1B3lQnf
HMxEOD0p5YnRtWFTLgw7I4uxMCEkAyxOiER8S141OjiliTcToJCSC9e28iBPqGqI
ST+me2NevOkGGDeKYP2OGrYhf0xJ3/9OqBosL4Jdsg7bU0eQhsXcLB8FLFhOgtCm
BU/LnDC2wiOwba++pRPVhvNfFrwu4FmkNMYQ0cScOI6n/U6napDX000aF7EEzQWU
LcvQ+HDFBNMXDzyeC1kos6SzyX8kaZBQAuV8895Lxggi26iPkBoIrirTxx2q0vao
iIYmdIunHtG+n7jvLZH5VpmzrTchnH65Nk+B8PGRjROC6cdFQ8FB7xEfs70yyOpi
ptwj21L4+FtbOeo1zV1pO9FWaG2K+5b6MyL/ii6usv0E43pgy6CS3YxUgcn6T5m+
j4/kCjk8kv+ZVAQAfVSMJ+0TRyxJmG5gRm1BiZqSGnAH52cEGaBVsWfHPvyb4yrX
VOaprWgbFDGQNRUuWcKbstEsQEoyChXIjhzjJ/fQknnXjc+/45L3qCc/ZDJkdw/C
5RHHOVzYqBk+05IDc7lmnB60TaZ/5IC3MrXUjLj0/Lo7UELp6cHfmEqIVrirIRcD
8Zyt36EisLVNfUn7AlpBVYxh/vVlaOOfxj8u8i9D5s/Zw1K4n5959O9MsbbMYpMa
4jqnbrbhFqrtX9olY3ZhQy56gy2v6/MmYeje3Bss/E97Xvqj3MadRxskMHd8IcTi
x1jSey1agx47zyc8DwIH+S0eiUqp1qakx5xuobQQ/VCkBDLR6HYPq3OcmXppiDux
X9MDKwLIxVZoH638w6vKNJIC4WWSJ54NlA8DxUYnFfqqMlYJ3sODnYRgtwAJJhCQ
MNd+WgAXnFmpNf9vNnydUOFp90JP9SR4Q7sCDD3thKJciyyhqcLS/G377VBuFB/L
71PLNt3xc3PxWsmMaQaELgLcTGh/TatnIvh4fErLGZ+8KE9Ml0NQ1fo5IqMLd43i
mWP5wwGbsrfg6STwPzsvhKFL1ZU0LWcRCke/6o6JGIbWhWosdbAb3Lx/ZxnlaLqm
9RM853an7fSCBt3gxEQ4lYwogfYQQDjUrcUiISO1S8ONoJI/lpTbURyreZeKSboW
vA9WBkAf3LVtSe2motQfyJCWN/H1mJd2HAKYME+kMmWiU81Lv8A2iYKFdwrqp6IE
Co7AFPMIbNh8izWULH1JZzYjfXVQFkEpPUquZVMDyk7OsPo+ex9F7TrdEP4C2Lp9
gWCeqFtu/dXZkL34Ud9/0QobuSo8tFFO0DE7ImuwdCbTc4mORAVZgQ6U353Qlctj
XkiyH+A0rKWyerfTLzFAB3BD7yaxVmjKexOpU5p66ny5PoXJUHk8EaVJ4+VRTKZT
81jlyKgbOYpeHN5zB1vj894KK8tOz55fKrHVT8H5xUu4AsyQsIZpAn4mOrp7MK7I
9FtwRk9585eH2w3BHT4eRlJt1N3dZYU2if4M87Tew4TXKdcrgqjkuDgqsxUEVccP
/FbCMeITa19qz35vlE4UaaVKJZelzkCnLrJuBq+aSkNVVBumJdiWC9wKo0cqvj7p
bi84xhlkyVK2dzR3/H+llz1g6nd8qk7kyTxySjuB3k0h6u+FnDcuAYUrbx1gUDxY
P4GSc1pjPgFmfLRmuNpBcVU3QJAdj3D8p3tudPe2rvY1H2vzzsliNE2KHINRebCH
9rP0ITRs/GIh4/UQ1ePlHPVNg39E2dtGDblMbCXmcTvB+g1O/9pk3ZrWwaLjxI+U
DG2nMZccKTR2OPXKRENj2ix3ulP5f+xue9MAgOweORcPQI30rfzyw1/DHQt1JAD5
MVP5F5NhbjrE2SR0vL4ko7oit5WLeXqg3qfQxM7wRfNWUoAINlYqcij9l2SrMvR3
ogIbUrdkWTn02TbC2TENK/vRbiivPFCKoVz6odol8jM3h+dZhI4f5Cc4FZogU3P2
khFvjqYNHKLqFpml4jxvCvWAMSv36rjatx0/4PtDQZ4dZPh/6h+9B8zoYHVpXTqO
kP4gK8o3DDOoLl6gUYPJe0NLBJM8IjK2p5krqTg/89d9l+uRNZ5Z9TKuId1DFhTK
N33uPKQduHtG/vG1W4nxGX2zjSsGOWYZBTspD9XeOyw4xzbVt+4jyjClDzhujp29
4OJLicYS5gRCipvZ2Aq5hnAxAZo5DoeRCnogOTHXuCyQRF2SPQLHnh/jli/h2CYy
KRpTN6Xs2NBv4n5JAsobUOC1funSHmMXZFWjvVtWIP4wCKRjgdGUQWNNDs/NbDUv
lb4w4Fh4GA5LnlD4hj+cpMwE/A2C5DVJirOrbZi65X3bTFVJYVu6N44wTFDrk597
UYhrZDYnlBTTFGitsX7GBrR7JFKUtBj08p3k08TSt8pGUwhUHDz3T2j0UEDBY6o8
rzEG7ZN6OIX1riUu9Dwco4hEKoZHS/tqoj+Xgsl/arDQediUEVEdtf1t/AgCplcB
yw+2NP6zg5GC+9ZrBOLXMU5cxJA3KdL9gx5v/3umyxpV/eaYoZYLkrebO6gVtGze
zHsd8/UTHeHdRy0K30BpLZDadVcj2pF6qvt1cQI+YylWxpRuIE6PcbKLMqbTm2xg
7o6aLtY7uh7sEE7jyKU9wquDoASJtiA6A+kmvMwYmKidqXbsTbJXjK+55qXTsSk9
NWYMcPZ/K5JDT0hOTvVJ2Yv/hRvcrVEQw/6lehH9V9jOY/6HVvCsW7DiDJHqBN3o
2sccp7E2ZSjuD/BO9xUbeLiC1729x8TqHF+eJa0pR/fy/dtAFH/x6ONOIHxv6l6e
fzfkT/1qdOCTqjHqt/uBbfbI1jUXwFpyrEkcg2KYYzlAS/5s7N7uprXQp4u2QI8S
mL6BK5fxAcHQhdku+SoVRFt9PHLrszMp5KgSZNhtN9hxCJ/4sdKItaW3MZB6fviN
oVGbR6F4BJYdVDPX46Ac5F6yPBwBtbsYTFoYoR5NemEQ5KNbR/Th/Qm76epPBO8R
E3D0KmyjvOBO48NVTHu8WvqMfvIyUL7bTMRbZ73jiYXWiU87YVCbhg25D+yDbFl4
BZVKllfoAOtmv/gKcAqkJ32Ayr2P6CNCSXiJ3oIgFo11hf/VEiR1TviMnMNSqmL/
QF1C+K3GJguTz7+0MEojb+mJAVDqCj3B+oLqio0PQCU1xES1KyqbIMPOnPPWU2Je
JqzhvCsUeMjj6N0nT0zsYlQGmBu15STaobW03nkhRCby7N1vD94aLQdItUZokQdp
O0vfe6gn3JroulzDdfeCFMEhvGo0T8IUp239z37/3idnWeRrZr3gxU9JD2DI1bWD
TAWkxCWaUm00soUF3nDsSDoTAqsji6tvhHIvgn4inCLytCmlNDMjxXBs0Kvoy7TA
AfF2hXYpTPh4d27yj3VmBmimD+EO0WqUfYPFzST/deA3iu6cOELL7pw/dSh9Ki1u
GpNgTFWwfbDDjiDBgc1Ku4lfhDDYNT3ZjgiTT2lcKdXXzsX9WkO7I/3zEHn5Erj8
OabJa+A7Utx50I5+K7XAZpbq5pRSuD4xe0xIyzP6h4HbHp2gGnWwFw1j1WoJtk0L
8SEYgXOtgpfivsKxk2EggX2IyZCRwrobspFPXL/0hDTal4jiQateKObtvsuwaGw4
HlpAkyMvWRwu5+9QETJ5euwO6v+TkW9D6cF+HRzXVmi62EDqEvYYff5fyYHF4Foa
e/Wev1wo0wzb+GVkHMs/ng3r2Gl3UEmOrMjFgarJOHzLwInG42O04qyvC0oN2aMD
coK1ELF2VTsFbGlQXSgKSNuHz4c+0IyjvPzATu+qKklY9LZeO0jhSGrA3nUcG0ar
QkTWKob26ZEXL30Qgj7dAXe4N+nK/roa291LdAvS0UKsuqsdh7PvfYg4UJE+9p3M
e4Wvj3IL+QJSz/lyhYd7AbQjazzrobPpuFe1fYI8K6EcF+d9WtzcSshVfMBKPSwl
eLJC7fTaTL4qf0X0v92CVbsMgNmYtDZCszT0+8rKkwDerKBY+gcx5eAZyWDSIf6O
qwYWQRocl1LJf+gtKlBOSbayD+iLKnizvKFuHs9GTEuq0fVFdsi+x22PpfrPE9jj
h2E6LRC9vuCRkoAVZrVK2/4ECMOWkwdBQ1NcU5vALvRf6bNSbfoBykiIr1A4DRYI
BXiDmK5McMA2Yj1WiCUc4d9icOEKq8KiG/UuDIo9UXz9TwjtpTGkJbTGT7tBcr8F
c3WIHqTOhvGmcxxgjYe5zthC7cAftSvJITnbD+U6rqTRilRdWlPc8FZdaTNsg3Xy
kjcySn5vUdVvZE1rD/7GSGNdCiMiChYONKhwukHDzoKK9lZzD44qA2ftQ4LYeUH1
PvVmpGlOU4wKbGPDIiqmKDYgjKFyeG9kkcLBEjXY7v91bm6Za5ksVOOeTOwTVU1H
ugx+NRUiJvde1LlHXYVnwxsmyBd3GkrzdQlsahhKInOehCuu4zMGd2kDY3+moj0Y
+mysAvXNR9yRataoB/giTyVg29Z9NydIaa4o5HV26cTgXrkk84mFVxfrKIL7xaIg
K+8tFaEuyiYJjtFJZk4p6R4GbHxY8bln/Vo8dpA+01+QiHrjXReUw+9C4e0O3p2L
59vaq3B18mQ4uWD+EOvsly0EMY9DowyHe2h7WNCINQyxoNOErSaE8Bzla5ADof75
4eoANd9TaNfLbv/8FWOL4v1VIOBrVm2pAbsyXzh1DuqAcGKWt7Y7wprlkUi2Bcr7
UmGnCb8wY3syox2b2wDczpH/9wtU0iXPJiOftt1Bk1plZ6Fk7c8xYfFWUnu2epja
b4hFWUkkuZqATT7fxFaxJsAod+d/y6VG4csgS5HCBXaw7t8HMuoo/qmP7SdYhIQ+
AXWU9vYpfoBs6FtH991/tytTcnNAI23Tv1QhVSTvVYVOYbSnpUTr1d/Kdgns3/pr
eUA62dUx8rNGmciHmwt2VDPUm56IQs/VdAwrQdzZ8IBH0RW8IMEYL/BdAk8kSKrs
cdoI95NAzcH/C/iux9Aq2P7s2Gt9Ft3mvSkctftt9kf0QnPI+d5cCQ7Xveyd48tI
XmWSvhWLWHEC1XMy2hPtEXykBSoIEmX7VLtFu6g3EZaTIre5ynfSwNQZSHc+tjmu
Pm7fVwbjLWiCksE5fhZ9qISR3KhnYBz5geKAV1aImmpxnqSUah3ljMe2BMyQ2yZu
MyxFAnq2n5FjOJOahsxDHwWNznaJ1GdtX94SmGvFusUbWB17rHN4kMlBagOj6xLQ
P/k0GZcCEW4ID27XpAXfs+KJ8w9I7yo84PPhxTML4v7wIVmRWatID12BQWmojnhw
ddtrizoRrMhdEpjqSadQAX1Ku8HrJ+VuCwfImWRsZGtHlB24bkqrMc+rfgcs/Mb6
ayBlnr3ZJkxzJKMbv3pzsqh3e9NbpX8zfhnAVnvBrSNKJyKV2Nn+Oi95TM65Md/I
QdHcfpwJqTllnzxERt+7oCxKKvk10AAKWPJ3sEDehUe6BWiB9aDIExX6qepot8Jw
VVb3g865Jl8JnN80/PoHmxeUlEyLJtpRJN76rDXdlN+4Gr2CvncFz59k8Z8JInLN
H/qq752uJ22YWbdJrnS0VyT/vDDtWSDqQqULmXN31TBqMerTcK1kJXV3br68qNPY
RlpRm+L2QmqZfWs5MIsab1K1qWX2hO6mhZweoF0ODrvnvVbOXHiu1zORGwnWdrOL
V3iS/k7huIFNbhZlTKOdABKMitmk8nljKMLGc2r8SOFNK8YjLR44du2cgvCDIcOO
Tv3B7Q9MDDzAnDXwVdnGCoIAR5XH9ZNW8a8RgA4sxFTQUTQUniQOTWth3eqhb1TC
tmrcJ7NcqSlYrPlHuaa+/BUC/tq46zz2xfURT6lO5jQ543gYBY2ayXqhgbyG5yaY
unv5AE3CULfKlnSsoPMmRU9D1s8sAfvHvZ65lZkZkfNgibn5w+y2nOdD7Smu6SdT
bCykbPs8NUIkZ5acfniz84ssPSx9shkmPgabhrLsyY1zt93YhwWxbZV9ympDNmLp
RYILDg6Vq63M+VK78SXoLrShzp0Rh3AJdiY/hpTANX3scbCSiUTNq/8mZ7YdXe77
c6+3R5r+sMPPa6egVh1R9KrUlHinkZtwgdXm3z4FAI4nhfmbKwen6lEMeM+O6Bev
1e0r/e207fDOQr4XRkvl1BxaImyT3N6b/rGtwKIr8DaT/VifeID9kguueHxVlnPk
mzctMQUnbsJ4Ak4ocM8rTx9AxdZQltWGetymphRFBIoxg6ppsfoDzx1I67Jb9YyO
GvFi00VwYQNN245JEZKOFiMmFSBRXpsgzQYHtdKzzG6AA8Hma4fWD91Ckqqs8J/t
ejmC3vQqvmUlYV6dg+bGJ+7fKezUclPDh/r2fb+g4CjWkmlftGWUxkhclxnsZ3LZ
DzAjHNNny5MeLXYAetimx/eoKlN44WvxkWr9tGT5rZpqU6q9RriL093+ge3NId1z
8BkEMn52kQM3qIHr4F5kpJ4iVm9JqkVaDr8DbTEpbslpS9jaZv2lMb2q5ANzqn0M
UMDrSd43NhMyimX5v75al1CivpY3hpO6VQUiEDo/7ZUuJpJCohsNIdTLSXqWT7QQ
ss2+z2ltKW5A4xVI2qk/qc50HRSJQTuOy48TTWI8aFF1OZQ+6cHytoU4HJrAqDWs
UvzC/B81qSPgrqrDZdndPHJ9og5p7XJRpOUJbkVBIoXV7cFHab/OGCWTRMTFhwUa
PSrEvJd+X5K5GFA6nOr7tbbUl3ZBwodIA+PHWi0+cxDszOwJ/AS4qjT8e3RD5Ibf
6/+3abZaEm3IoeDKiVuA4QOeOVYSHILHokLDSY3BcerjBTWXuTMON1+gs5RPwtFV
XtmpMNJiXaPBeSYYzIBw8wE1Y0ZXZ1SMXF0U+W2y4xDfBPDq8Uo7vfYxUEQ7wfjB
6iAL0G03CeLCP3PIu6Vt75vFU5k3Uyr4KVpOHETp5NuZPPaDpi5zs3QsvdSf4bSt
IxGtWVDwmRFcADNcRqgRKGI02cPEzZIUSYUXHqzVpAz9ZrVRV3mUVTEiw7+MA0vO
RQQ+1q7zH/tmtkxAm8ZC8xJzWsNag0qppIhUg6gb0kNlHOr1M2xdhle2CPqa+V2U
dKp/fkhJ9KdaEFukVat7WUl8/PORTWxGQ44SzZbfUcyu9AcFDvA0O2ji9VK8IdRJ
w76BMmwTIaqlT+CpMj5quG+inx1X8xaV4P1elSxH3jaoQLsGHrgG9Kj6JULy4ba+
yJ9a8HkfIptex9lDI7QNFQ6Mkw735HD7PBkTzfZzXLXNDKg28mYQ4QEgRO/v4QEz
QTky4EdtXYnzLQtR8vqO38UFwbndRHNPVXrR9OP+NorUkg60AR442r+Jm23pUjRV
2x7fRRjrxlsOrl7AaGagEhdpMMD3I0R2ZmckKTscDVBHdMPHAbvFYHXpKDEG5KMe
OSFKBiYkZdkPe1SzILZ6WFCzsnq47Pa6U/D5BRwGL07Curp48rWeBjcKNCs55KkN
FwMPfq7B6sYSWkIygZlu1U5tVTm2rhK96WEaGY3edecsxi3Pfu0JEnLo4DhU2q1c
jSxHE9aguzSaVyyFDR5rVkdnuUyEAtmunwmzusIYuHUrFkCy/LhBHWeRlu0iAppo
NDpaNCPiXBd2V8XV2Yva8J8DiAg5jMPBJsBgbeqpQT7BKOuMcGE8bhymn2Bq9FyV
+YwawYM7qavVxwfebVy4feSY+vDJ9tFNmyAZn1YSIBM8KEO51Vdu2PTJ/CXKGhdS
fCZ8uHPVAbC5gO+S5Tat2YIJNvCMnwUQGORyxAUns3pWlgfyYpXqk1bSNM4l6wSR
Ow6uiJbqAr6McPqPmAWDCbe5+sZwiU8Pq2j7TQyi3kQKWSdHBiDIpBOdmdZfFNPM
tV3LRqrS/QTtl6YwTkb5oS7CrkIyU3cS/ym3pr1MFADS3ByhkF+w5grhNAPXml3E
/DXyb9O/iKQt4+RwvKHo4m6Z0tQj5QQvvmz8lFJbL3PH7etmYXkTe3NjP0dEQeA7
KM/lZlJv9q6mgGu2253pXH6Ltiip1hd/idHNxSLI5sccggh8jR95Fw24r8exEwg0
MnJ3T4o7Sxc8rgdZB8v/x56B+1Iu7MA1ikPjnhLjcm0357RMLkeeHJnJNYTuZVAE
zx9PtJO+TQVC3BWM+gBxny2/hQ03kLTV+xgLDtPfzRuL29ab247OEsOqvJPWBJUO
bPRJJyehiLnPnr9iBnT940C7o74W+ct9H6bDT1C729ctI/bJK/mUrTJV5d1nXoLG
4E02xda6FUc6SmDnk041q92zzEl1L8KCCCGPyzjtrDSvvow6khVkLg1iKM+YmLy8
vewdl/R84UNqEYKz/TmvhaFqTiosTzYJLsRaJNns6cInCXG3XiQC5/WtUrtuJqfB
RdaUUojsjxnLDuH8YM3nFvecoazS0w9h+YLUCiK5BS0cmOmbhV7GYppV4oN7WlR+
nQCKoh04tCyi5MttSx5C8FBijywj0Nfs7Rw7XrjkPajq0Ti8HQYz1SY0vybieGsr
QFTtwTdUJ4Xdsjk3UnFuyfaQZKiHw4t5v5shoYG1RYmlSR/i6Gt01UEE68JEwet3
LL1uf5o7/Wjd8yIuPyjsTwUWsHCrJ8PGpTF3EYt1OdPcQmWLzPvDgnV3SypqOtHY
4ZoTbvyDI9fWtvNeCzU+9XJLIURFkjAYVI0XaLQ1g9zT20qQydNRR4va/0UsE/ck
e6RgHfgl7qCOCXRomCYy68Ccn3nOm+TTVTB6HEZ131+rOksa59EWWvrX1dxVPyQq
IfJ5QiolybAYvmFfQ90B9DGG1Z82vPSG1C0JU7V6Pp9Sm1f3hEJFxtnnPBSwIPZW
njIlkadKjLIX0clmAr5g/3AdpjQB7gewKv5BVzaPQBSWaLOJKkIgOEfTXcfeQG/7
jcF4byED9gLgaa+8d5dMn5L9EjZqPfXMECyCpXPqxM74u9cIdMkX5cZWbLqDT357
FjxzT47ch7CICOksVnph+swRwZFqQvVqkKlbG3PsMNiInR2cW3AqY5w+AO94bKcY
4KuBchhzp06WL67O5tVHdLXbB9u/9G+KPKQ4C32ALCh7ae8Zvi2jAmEq00rFAZro
uPA99JizNsMtYigv7BIRRMD91RNYkPEHi2oNEbThf5nyTHVlCE9QRiZ9Gl4+Muii
cDA9IEcVVdf+6VV0bSO8d8hPnoM2VchZrkwgpsqd2DDd8Gnk+CPx0jwml75eisnm
4VeWSkE7sHx68PaCliwcxoZJqVG9STxnVgktdqXYWMj5loEr1IJYHcu4BwgNkXB3
SPbRHUFJUFFA2R9Hk/W+qeHPD9StxTcMmv8LHl6IDxzQ7BpwSSgXJsXtoRXrMpJK
OaXxEvxI6VsU4kW3N6qKZY004wif5yLkiwD2q/g44j9xt7j8FXo0rYPNtw+IeWbR
6BgyOXT6nhH8NLxX7SzhsbH5u7FQheWSIxxZ9bgUhKtUiMpjCyApkioM64C35com
ocr0fuwPcCAddGRFactAw7b2DdjUa2IhAhzM26xud5J+VMyzXTNHDuC96tR0mbeL
NJ22HJGc36Kz3MWvmiaMpm393OXfXGbbTR7n209FbxTaTSj6dk4Ew5516xd/bklE
ptnsl3m5ufSJynWD0R57WogSl0cccwRUVEKZWSpMcoirrgPEy9Hd+nZ6VnKIpxFr
6CrF0XBDNgL+o7rZ7fWeRRxQn0faVPjzDjn+zv6OxNEfGETfMBfVkN0vB6Cs+ops
+hIdwTR1bSlNqUevE0x0WU/UW1jBDbJclY0tD8Xr7XiekN6FpbjP52RnaNFbKas+
tMW06CWHcL4+s8o02sYG/SM9cbvTq0uovvMJR4Q8VxXwlG24dBkxvFbaXLrzBgW0
ZXo0DSApxfw3VlX2xt81YAziTV9kq8mLx/LXWEjwjVD6IRFGOds+/CSIn8l8KTMM
LiDtB+9Z9HA7uFmGtJwES1yAcBh7r56wue1JonQpmKzmPSaf/CEes6kN5C18Vkdk
MYn4T3XIg4YIpnu3rLNIHw6nszxP+iI7VW7B+H/VooDau402e2oUfnL/YezgIz9s
VjDDjTcp9RyT+cWfUQ9sAsSmd4C9yh6WDdBdCJoYhDEm8bCJmZo4lnArlGNZaEIy
exf1wOfpM8EAsHHeKaIzV9yKxGEqm0XwpYufwVqRJlRnk6V9KFwyWDBTgu2jfy1N
Cc1oFRoC4Qy6dD68OuFb790w6k3OBjgoBLFAZ9u1YKN2qDyJUftdx69yqh/dVM9n
mMz1/jXxS2HPikA68daKXNxDX8Rpjt/W3Ahp5ffezWxoTH+sAwElUAXYHeMKNEce
u6YJFyJXjIPH4c1IpyuSaFc9hKSXOOWY1vI8D7/187hxTW3fIKbopEAxKInXC6Tu
4pZDpNA0juI62skb50qGDzQYpsjL0YEPQ5y44TCfnL+w3Umf0UNkcY/SnpTDJl4M
EeUpEnXTlRQ+Ju05DIemdlMwKKR84sQfST3pBSH8j532sc4uaqgu6axmDL7UJNQt
65U0dvbk/tEPwZVx6fjlqMjqn2ZEujpPt4V5dHAkLrmA+9MXxcAIRiiDLWqP8+Bl
sGfbtyYdZGujdy2dn/XTM+zpKQhA/tbYyEJ6OAZOCEbvdqHH3kkuwXDjGHIqVWmg
0kZ4nM8bKlkAEuv9eTTV6Y1g6nKzTVFKkzTVQondYkUFuJLRI4kcoeMA9Fqx9Vi9
4zvLq9F27yEQyBrYzrBsMvBLyAHdrGCrd6oX+MRUck1/i8ILd4f3Hl3uj9MEqqK/
SFz6UW7aSjmRdU+H8szPymR+kQiIZwXYCuPzXHcoW/11+lc9gmspRaNVtCnz/79h
v4SNAOklsu6H1HOC944XbTs2v5YaYcCdMHg0AiCHpINiHNlPOJCaZKveWVLnTL6R
kzn01+i9ReqdJJrhBvchOIedSHRZsMyZZ/QReun34ScABXf4R7vi4DDXKybqQRaK
IaCf6LLxBK166DdFOrSh/vV1Nw8qQ2BTE1SN/XWXck9YTmtnFVboUJmRVn7dlcwU
U9PW2y1oCwwm27jR51k3tyHaa7vYY2Ht9iY+kDJP2xjY/pHlJ7fZAcpcrJa1tgZ0
wM6OjszLHaFFMNg4OFP7MvU97w+IEdbxNSHD42GcpfWLJpyQG7JZOkR/1UFDOwJ2
vK/10biibLV4nHz9giiCd/gPbsrw6rguzqfMYR6iu6DwLLNz9TseNa8bfCHXxrRL
R0mWMUYrqACrBrjlinQU+wJb1Ao0mFOEn3HZrD2BK8D0vQZlmoMel3UmcXNB4yDY
tN4esIFQOY7vxcK/6gIyX3AgGwP6vXX9ioNHjxQ3JAzRXI4HKiNpEZFO0GQrdlup
/UeRrIx7HAHJS/B/Uji8PLDfK0iUQtvRCh8EaZKy9EkG3ZFK6uHIWyb2O9VnseK5
pQFjEQ+s9WW9Y79CM2scmBtAxXGxRP5k8MVMr7wJ+jzYCtAtuaAN6jWkROvvzkv6
2OZUL9ue54UjAx1CI7vrJzoP2NcZhXzkaRTBlHoiKN64xaXbA7xHklXSdzmNK6o7
K5Ry/cjcGTC208N0zID8a7eOPmcbrY0QT+o/Jm7Pfmu0ROUA4ild8yvFCBjRwdaJ
Pm1t/rEfLbOi1coeaAdeR+KOC9gCvlsMeTv7LLUs0JtYCbZgUKJenj3KkVD9pAj7
kZuOvTPhInEmopBJqifxW4y2Tn8NLJsKYA/dE4kuNGH9LnRDXSzY0WfujJGogCD2
P8NUrP4VAzUF4pAtw1z6fghSErvWTVUAkumzbqGikvrcD3ocrjdbaLYv1ydZrS5K
+usNXmgAYY17ObtqN0UFmkMlA54HI+zZqd3NVRk/+NEw11AGnYYBf8mZfsDrItC3
5a7BCdLneKQRWxeymYSMex/Wzc/RBBJmhtguWKWpSarpuR/Tdw0mrhG2ewt4g9Ir
Ae78kRTlL9rN0MdLf0lOMDWCwzsnKAs2ewLTr6qccXJb/VRvxtmAXMN7GbxItczt
XvjjGUnQ0DcFRj+EGEnZjrrjQExc1Mstl+ipZWimKwZzVLR0jKCMn/eENI7fWUEX
VKwSMQ4iLe6uZ4NXOOcI8+mumfuLCD+/ec3tHG+4X2kAR1xqqwkabQEJXnrddE6p
Gp3YcxONlKnxHeepmdD5HFav7gZhTBjU5hQeGGcUzdW7x9AZa9ZncIhxWbSWVcOF
9RjS5GrIqPTfLMCC/x/RvdhlgwGcmYvEU/KX9OQwNOjnX3wbHgMfSV/COSPE3ub0
2sGspYWHwnQ+qw6jnLLgNZ9HZ6zCW/wgVhJZQR+MfeFNPMcEfWnaLd6YReT4oJE/
cgwJ5UJzpLe3qhBBHl4TnAsEz0O8YPNvvFXdLejskC8wLpqGygfEIpf5umj6djZj
uybWC40ihy7ojZlWTtaPTn882WIgpxo/zfB34NnAggH16eFL9QFa1eHiah5o16Wf
iEWWwqroht7Kw4zVpgvRTYXBQaM4NI7evY+Xh+j6Hm0vP+pAymrg0kxjwWfhG040
WI9QPvji3bOmc7tM4AoesEJ8000rtcpa6tVpNtRO1W0LvnVNjniZ6Za6thZDnSfJ
L0oIsRX5ZUsWippQF9iyR5oJnRr0lr7XnnBKJ4hRh6yVZKlrKgNCUskIRcGs+HZ6
uTFwrLhiFzPE7YbwHfhTYgZ5CQ/ZdMAtku314F0Lw+vHzeNFbXwQnRthd2MJaQtf
9GOvZCceygdx0bkJHD6YLT1I5qvvtAwaiUO2vxoqVUtuBSZz0o4aOORDkE5+a1us
f/beM7S2F5RCix6GhinkHhVgCO6fx+DU/u63IjSywHD5et6fN32B6w1OQNusDJGX
/TI285A1Gi3krlLgrUW/rphboveZ8jU5Ed93KCEfOYmx3xrj64kVU1zazycw2EGb
BbKWJmJRIKzTNBaQYB01ojDmbLBN79qiemKsjNxiPPUg3y3e9clTIj/Rh2D7sbIS
NH+y4e0BWFLLMbKN5XgMgevh/yUtwAABdLX4QLYYocADA4B2Lg4TB5rDZjo4ZvQv
tYrw763wPgqj2EiNQyqwhbT1j8E6M9Nf4vyLin4hbqkdmjk37FKkiqkYXsGz4qW8
YXAosmGiov0rpD6NZvIQiAO0SLNo13IZmLequFsCT/qSgAt3rbb5rfWsVvu2PyqP
HLPPe2+btYFaKSKaIJ5YrMu2PqwgTxLagYwo9pqldRbu1XcJEno6pAEvYocVCYCS
1fj47ktdi4G9UuAUDiCiOMKV2lUK96DGmn+VqtGGWmW0GcZzxuQIMhfqU6b36bqm
lLv7DpsARTUdRAYu8FUfPgxpBHk09P7C/9RVdnhzaglE+XkLnwP72/vamj4MTwpE
CG5yDHuj+FRR96omKUPAD6OTbo3zAfXb836LuqXbP9nuyO2CcMwroekijukJO3yb
0PXsfYen4e1p5SpvGbZUm+9OzjxoEfebVHSWbfBHDFvfIg3y6iHyaJmqSpDBfTtm
Q32B7t5zGch6iUs6JLRNyaN3PKTiAqd3eMkz8T2iEr3tA7YSp58yUx8LTDXVfysw
VeMBo7GwWHWI2Fzvnd0TsMYmwklQrPg9Zxd3Xrzsj3HNENeJvTo4esyT+t0RMCo7
HaOq5+hZ9orpZ/6EGPnykIhrIAc6MD5QMwwvC2aZYJjDIzvCGJA8+BHOLzx1cXA4
7jaF3JN4zogLeipnYSXWS9ZSFJyXmzmhk+BeiX9mf4hVcPdmPmoWyrQwD25kIkgu
njp8fOICvErgFTFdlgMPtKdrOJTSz9ojlEQLW+W93wQA7VYfXiFRMW7Lj6DtlsHX
tg+Q99JvybSKIdfwhkh5FGDUrTf+Ptz8xqSfZ2WOMm0P9Wsf/jPWrACldGsrSwrT
b8JYBGgwVrewSeRmEP7RUfX5pfXyoDYwc0ngWjg+HFvdazaCFsvaz2l7VjnAYMb8
RJqtR7gqKp8QKXD75YgDF5xxM7pmYNNBTcx+/khb9iCrcdjkQ1rQKETyftyUG1Tu
+UdmlhPUqJfkaIJ0ngospe7/IO5vcTSsNI4wk2Gffj3L4z8Y17X9Owm+TsIbchpk
cmpoyxN4AtuHjOAOxe0o3kAUMTFyFp296h9sCo0gPkltEFrumz5xg861oyRXr4PR
WbuEdB/GrffYRoLDuVX/2/SY5yxv48TYtPr+KiRqn9CJ6VtgPotyBlnxaHEgUZDR
d28XWNd3SbyiQJeLW1jwKc2lQtLeKWN6SNNshMNu0ivg7Q7qCdMoWFr1B0/nPxeH
MsMPCvvzpCPjDx6uTw/FvreBIX+BmFj9Ylh04bUgLHXknlBbCSatK6gK/o2EzRZs
+fi9ftRzxOdaSk6ofY5gtsWQ063pu+PSwrJl7X/fLkepqKZ1Q1gKEmqwAqEC37dO
YKqYvE/1wDwo/R2rLqBYqFjjASvg9lhGh2bAbYaR17FcESsvXnHwh4IEDJKNfEer
88aAtuUIxLoK2JQjVOgUGS9S4VsbhGD/TTzhVDY7sTfq5RyNm1BWPMrlzwmJqVUR
P9JXNrYAmK8pub4ZtugUbvcagoawtG0WyYFncpXEQDg8DmPx+2HusTaJLYvYWyYK
sEKrNKoAC6fN8ZrgTNiLebOrNP3p1AcHZbg1pNFyqO9aywFCALlkpbwxCpTTlFYf
wbmxlJK8p0HH+h8pHaIQfGOaCXs695owkhbMbI5R6/PV+wA0yZFQ9V3OPBVvF0r6
fQWmTmjYgz9kbVYV4jz1b2e3gbdaj1ickXmNtEB+9LXbcVeoP8TQx3M/Ne3qeWAi
iylsJyRpkpr4JlxPw+s7tNSX28DMLrvV8vZGbXBBSoMddfEaw7OGCe3mKpymCh17
zK5L7jh47MTaxgHMi6KQVSTi8pnVgMKzNRSQqN/0YySZSS6WrDGcm8opuqAIaqqJ
8PqDhvyyR6EWq7r1JXG/LC9o+lH2i4JIsKAaG5ITdlAnsTcXuzAbrSsOMi5gPRA+
xnYrY9xpjgBKupMkb1RcTfwSw1jFD6Q3oc+upH+wKFZy5TSYPYbC5fl75cDjEp+G
JvNJ9yLHy8hwWWEg8PCQb5jq25lZaPhXLqz0mDctLBnO9ltx87OHMk6INf8I5CMP
kjEM0lAPmPonNTJLbo1AkjMU4gtWKw0E5DC5OuseItN5UmiPmBceWqGugksbeuoP
2R2kVrbZGT43T7asdUxr7jljTMJdizQM2kCTGOxdVKpKBN2X+0dws2amc/arULq2
M9C8+4RcLMDyt5EXSJCMUrmMT6m3jUn510aQ0TgCuG8z/POwKrxSk7ij2V5xzHT+
2nl5igGcVyawg/gYyIwrSojpeCcj93Hy5cLUO2UGzLW4AQ4PI3QkDBOZth5lAsBB
phbGeXlJ/adgRtxXqJpgAiavxLkcRyiumXcVGEBF3fOttfNBuXzU6K40S4GmA7e/
nT1MU+mIsaj7gWd7Ea4VbWpBIxpQBPW4Zl8quvwQUGlUKzdNq/Z/FJj6xvFYejzR
WP2BP8q2z2w+3NwZXrP3Y/KdlUprhFqO52IUTdYdcMJDSYRcHLa2GEGsHTjGjKS6
jBna7sV6xq9DB8TDBy1iWVCIzA60ccPVWt44ESHGvrD1mBWzK6ihg4phhiC/3mh5
BTz+LArAUFFoWAGs1rVGHFmDP2li2SiujokHDnFODuZwE92cE/GKQojAVQV6kDYY
yxnnPY/hFWeVD01K1ieqbrZQ8gqtUBLmiEu0vHkjdN+G/9NxvmaAtmdSR1sHG6gd
3UgCpIE8i1ldC8ZvNCcDr71cHjp9yueah3PYIPoLFwL4YDTmETSwg5k76nraACa0
uE6a2CNtRUxJUuO75r9gSkw3GABrGQD3ESvn+C2FwqCcN7c5bzb6mtORaTwWuOJq
O0ySw+2yCEPFpHtlWSsYaiBdYQtyPzvn2grcZoThNEU584jNfNhky78WKQL4BpLj
nkS7mwI76VW/ZZgFjKsXdZb9WFjLe8cTSKJ5uiI5IyBOkvgOGSpmI/Gv88aESqN3
ML2NtZcQ4tgL1UEWpIkd2U8bVZL1vD8dpBXFr7RuFhQAosUOwG4kMrnKCvghnyux
IEuPTsb22GZ791nuN69q6y21WVUICQVbrJ2D0UT6JDYMGDA6SzZBKDEjZ6gfW/lf
gStiiV0TU4N9U517oSHlxi7Ml60p1Gb5YutDjqvccnCmE7FUIXdkdRG3sjE6E5pp
EUk1IFDThOzs6aSMAu0li2KemUjvgqcFvaE1euBXWBIPC7PR4dhL5my+CO4XNx/v
OQk2JxH5ph1BIG/7oXpi/e1RB9NKr2Wh3Cczy+Qz3u2U+SjxVzLEk1xzJB4nKU/z
MxZ/p9q4R9YUCy5tCE7j7nTgzkoc5xBZ5UYFtNW4lGs0TF0Ig6B2HaQnowbHcpHQ
0PljREQvgldOuTYoPcI8ZfUswp6bTPa9n5CTylYU871A5pDgpeJNl+hGzdq0eNbi
ZkOSZEnzigFxbcziHS607dl/TnwAl3Jw4pVfkVHE5OfTDLaEdT+1ddXoUkxD433m
qFdPnHS86p089DsB+Uxah9d7scbXjY9gCZx6wGLSQfK749qo4Zn+7Gp0ShQYatmy
shEzkGlUVdm9FCzaYtlRIkwxar4KwcTdsK7P4Z0vZ2LZtWdNotgqBtq0A0MYyYL3
Dy2R7Dj3zl3Gb+N/Gicv0o4+zwpPewovYXfVHHzPhYcxy7DFVWs/zQe1ktQ9iFrJ
DxhYeGkB+Um7ZbpcIsLzseyjVTr4ckFtK9jeF/37dkjJQr1umSLDTzJ6Nwoj+G8r
yZXs38XSAhm4BKpiKhFiJHH/WYGp6vYp+na32pR4Rm3JTWbelT5ZqFMWB5a5QNup
9SlgM5xyWuk2JGpj/mfE/RbV+F+6XcZRcXxhCt103uH7PT5t0oVIB4HWdnoK1JS1
crXE4kVSsIE8bvmdBWcq6bSZvX17U9bR7yXR1U5blYDEmg5eoOj7hCimXcvI5/+q
UrCdUqzEmKl+OayvIFRag0miLHhFMagK5GJEw6t9J7ZnZxNnKj25QT7GFOzn01qX
sE6oZFxVKwBXVfonSIUvz6b3+JtSvCIqvSyynMvPZjM1sXR+C6RXiPZNfmqGzVvj
mTMvCAlUcSaGwGKJbLk64afE+dYRNv3y3jq5nsxMK7vh8Y2Zpx/pLnFw+9Ss2rhO
90qUOjk4xoGScbSqwrQRATS53lXvsvzr3JiDq+Yok2/oyrofj5tYZlaiC8aomJZ7
6wH9PbtMkra3zZCFEm+URy4vozfFIK6nmGTereZ8Y+C2LnxJGodhYIb8rfPChG5H
G1pgJTPmlcJDXlXNC2PAJyG9nELydiJQ3tICERWZZJhckcZYg8gGLJSwp/A7+vmK
iXHU1o0otPX+Zd3SSQJogt4gk5++c61fxdrvAnbRKsb02sQf15jmsykOmALPmHuI
HNNGKpHRdcSoCExXEe8VLYKLGQLolGPE95nWQ9dS15KiFM0LgfnwvKHu9UcstuwN
Wqb/tL80aNTiMXZ4e1FFjjSPt7kMu93L8wYUgzXy0SYd0ewyEfuDqDd5+Hp8FWm6
GSawrNdhPNZ3tVSebr4yitfyyAlVVC44HIF+gtjzT+558bbiZBf0WxMR+7umKTIx
DGPHhSMXqR6tAblaMyuYoIzrwc32yBBfxsALq4qUHxCuApyoqICMDwsxE9sNjVgB
NJO58CbGfkz8dMEtv7h05J9wmPkWF8UzxpN5WOuYVAEzxqEV2FoSqwfRQrDVLggb
qv+MKybgwO8OS1acb7uBFUxS73c6pCuOhmHc5bB7A1up7cRYEiJEu5lhnWe4rVJ/
ZCoVA+v/5mV6npyzUtYaAY77kiAQA5J1YdVDzwiaDb+/cLvbA3ewPbbmcKeUIqFy
hzUyh9htqlQTFyBNRYRxZ2zKMPmU5HQCgDxQp0GRkBKLu5ULSoVl4MNgzc3R96ZP
hdIraBmjbD3789EfLvxoWkgIkOns4Q9q/oSqPwppDjCsgPm5a7xGBZYkB3D/z7Dk
Ajacz+/6vo1J01lxKSH1I4WVn2457bOPAobi6MQ1HS9vYtGI1xgVV1aUfpLq3NOb
/x7Rxx/XBaqugkhgdbZ5J9YB1C5H1nCfjY6HCqjto3d5/So34BgfxsHWuVitLOf0
AMiVft4pmbsZpZgJNAWIZ33bYIZZUGEwi7x2Degxv7cEcIA3wvxs/mQUvqZ1XHrx
acXEQqGv1wh1sfkaA8OQzRb0P4fxweeteAxywjGbRJ9yYctIEWF2/yVVpiVz+Kz0
1zxBdmxy5tZ5XHA4fykGNSQKYiTAXPEcVd6sen29XQT4bFal4yMz5nrgk84F2BRL
5HiybKAlsSogatLMFf95xEWEdHfHFVXmXKmVLt2hCZ2MLx/IZRg2q8LUjjJ/FSsl
CcVlqz+OA3WRXfR2q8bMIWW3CirGyAx6hIjzAHReD6YfAmqH41m8zkYSwh3mqfir
To6y0VJUINoBsLj9Uzc+4WQ+wYpOG/6BnPMX/AsENIbGepeBSsRe32FPnrQloypI
pqL1TlKwo+ZVj3AhbDYibA1HCbcsp7MvPgHbmM/hqTrDxS0v7C9PVPogHdSNT9hg
bq8Qrb5T39ohTkXCy2FW42lzM15869wbbgIICidGBl9p+rCDaCWrGZjhfNMjOD/A
45OMnHVNzhYJDakBOtU9/rOSdOWqKDbvtPrf+McAD1OoEH+YZoXNgpgZggPQu+tE
la0sVhVeEMWQ1IaJaty9xulTYyKVqhdTQ//GZ/GWzQTbmlvWyCy1h5eK69MPTNZ9
XWrKTs3dW8rCotjvkzvTSZRxn+4/ctUVcIGhfGfKcNw6e3yyzI5QGSQIgLTgR3Y3
gkFX/WnqDSGM05WNE3qbv6/LcfEnXr03syRQd/v3nQpeA0wxVfDjImOmZldix9Km
5pUGA+kQ3GJ7f0XVScGEYW5PNhnE5kacfYYagOevMwwAOC/Ub0qgEq9nqz+HTo8L
0SWQ9A/+5kNKQObu5dotzPRSJro659KJeC+DQgv6TmDfNR167h8o9+VFJbRYE3lU
vWFHmHsalYKXIZmKPd00HPdfGpo2Hu8bQO+YUeNkun9diIaroeuPNKjwDrcG3aKn
7WDuVhuR4DP7uygFcetkvnuBtzBqJMGrnkYB54PMumd8qh42yZOqriM5MEu4BHmP
GQjodsVT+QU1M5Amdc3mISDo+leG3bKzaffV2ZjkXhPxPYrBfIHfcFU6Aua4Ml8U
uG3GmfnXYBqHp0i/ezXX5Y6B1UPo0b0HDH4YMmkyzK1kd53BQ65eQ91SHgkUfafa
aKx0FF2fTywzv+0QRZK5xvXOVTso1qkJrcVq2rlKGu2g/LpuWQWXJziFMigwii55
/NJ6F+n74r0ct4G+uLgvRZt4PITDBnEHvIaWwbwftau7wv7wgvEDO1JN0A80hdIC
GWunifIZYMXI4a7pdxqFfPDPFwtB999LGr900I95r7Z/NHatrJeNbA+ifFpM3T4F
whI3VfR7bD1E7XOF/06mFRT2IiDcAV8kOHES/3JSWbdVFOYSVxcGxPJy647Uh+B4
ySNpzz0pVNXjOY7pFRKlgJuMhKUHo0wPYFCRxuxDHh9TDaLT4PvLyEMjey6P+4Br
8rpo8nDpBHp5ETDHxVWzzxiv8dVT62WbxkowPoijAF5/slKbOQQygRo8v8Uc/Nb/
xiJQ6SwugEsqwrMudOwmy6w+9OKfqHglQmpHL38s8ZD9J51J6ZZ1wHu79crmTRvt
diE137AmqA5KL+/Ra/81d0B0HxQaTK5mLYRzb5Lj2UC1HgeUh68mvCltOJyIyd5r
/zSqcjpaKGcjg+y52C6nq56x+SRE7If6AzlA2FqBR8VOyrRGCbQUieVhA3xvz15q
Syq2reeWOei9wYNrVshW68uYeuq+Fa1bxsLNMBTcACsg/drD4w6F4zZvUqph6mB+
vf9WKK15j1yL9ZFmC/YDDm+T2DaNws+d8F19AEKzrcIs/tzQd0E/YYg5sFjXsyyb
wdonuhgG8V5qDyqiJUyeEJXr7D2htEG/pY987kUCEI99REZ2DV+QMUfI/MHNPH0o
jFvDmuwB2JZeRQRgD2ZhVViwKspW5+idSQB7E32fkOSb0ioTl1ZbkajZhdzuWTj3
awhK7x0YAJ1rGjM8EQyGW9GdJA++dEKhH2VbQLNzVmq2kD4a0N4Klq82ph7/CVKl
2j97U1MkS6cx4M+N3ZIGZH1NZw/6A5PCHSHQ2VONYUN4D/Zd74eQ99UEBr+s1B55
XCSTaCL2X3afGWsOT2k4t//HF9DfOIu5lb8wOKoVX2qJjswOJChaR7Y1wqD4fAdD
R5DU35ygsCJDg0u7SX6UkM2cCNzG/wbUDZjXGpPVTj7x085/6Xlkn7Ld/qge7xcx
TzgA8UojN6IVhNK6klGHXn7Tl0QWVMG1Mtuw3H4m2pXeAzbLzONZM2usg/y1KNb0
VzTLhUchCoafT7pZeKfQ5ZRcRaqIzrvh21uzvjZWgQeV4fsCKMN+Z95lLsVzgRt3
AylQ9vBpRwnlNCb9l+sDgSkccDjFjOn3pCCv1+TYQAPerXeCvhy1Zla+P2h4scBe
EXgzXf+tb2SqrC1Ox7UAUzbAoieQtxEkAXcKey5YdFSPG08KeejsE4OCmp3+dGjV
UG6TTXi/JUApzEOGY17mxvnY3OGgVBFlPCa6aBObZvbG3M4zu4swSMhwoV+ywaLL
Tm6XIuAj/mofU3Q8chnx7DCqs3ONsoYC8JTI/9q6UqPJypfwlKdeJFPAmugmJVL2
Cfj8XJ09/0e8HCnMxZn/c2yxVvKzVJv1C/ADOrtcg0Fy1VLFSDRGYUgv8ruTfInF
ngpCWbokyGRd2AVQb8ASd6DyegI2Itnx46gXYVQ28OERSwKOlQrJXaCM6ueRvKQ+
Yz0viVZeilYIeWiwbDpFqqRjmphIo8d2IiggwUqyo4yCscXNLiPVYy6JHc+mB15r
D5//YcQLbNflQHaXomYfzbCh7OOprfzkcV9flOA5T53J1btLBSTOcYQBDDMt/Ujf
2RfmDMijsWK94DMb0dlbcDpchHtchQw3J2vdTAuM7pdZMXahqhRB0nSdJq6/FdDg
TD40hzTwieM/j2kRaK4U/huJzUKsdIKX1m1S6PbKLAIyZAFed8fMPLSi3Ob8uVgd
nBkEPe1boD+P3XzXPZPGIkeFQxeBkw6B09vxzi1X6AZUAojpwTBSRuES+TGCIVMD
aJHnDjL4DSFd9M3iUy72Tlqe/IMFKU9zLThxoQ2A88qpH62LWMCBv7oYh9wlKExY
Zy8NbWY7BGcEHMwtpJMnNavhq5+R0n5I+4zgQBIk0xqsLj95buEKssAsEUegWJdy
nhAJ6Zf1Wo35sOn/BrW0Wir5pr3dAyWtdwx9n8s9QuukgABJwFa1iqdyoUinHoGA
kzwfH9oKEzF4JGHP/ciHVmoDmIwXMQ0CwTMJUtvMfZ6va+25Fw9rl16yzxw4oOHD
OYvxLTixqOzDlplzsv/LBx+c5ouAsRNiYTcHZr/bZ8RPmzLf+8iijw6NS7B0RcId
Y2FmVg0Dh4E4E7Z6QrTwkgHhAKl5ieW3NOIiq5dnazplpEo8BULVqAqgEAfjZgwG
YX/Os41nyCeMGQzx6jjn0oUPRa7jQ7Je9W54XNF34/MPnGQ4nMfxoOND0I1vwl9P
p7Jq/ihSZQ+GN/yenxompMEW37C8F/4npbrk2MxCVomfOveQcmz0iKjb5t0o1QbD
qICTfB62Y6IChekegXkGSBYG5XqZ53XCPO0Ad9C6u99rcXREc+HkeWcGVRZn8uSm
H9bINwD++R86RyjKxaFDZey7g6Osk9G4ljadwRTrApvRvIG4f7qMu5PRFGfaHwcM
YY6rXlrWP+ceBsErf3wBVBmTpW7rv/UQGcTwGmJBwM/wUiIIMN5/m5NNgTanEwKO
E7vygHwbjgoJ9dXUTmP+4HxF5z7ilsuxloxPOq9m+Jkd3LEu1ED4WN62ZcygYg6v
lFsxYHp9UNcYcMx5WhUmcinyxkdW2D1f1+YwJ1XlXm2H58fHjZ7QN7DMXtJwjmGZ
+ziyJqf0wzssMu944cQWi/GkX4uWiL/pQ8XLK7AWgga3ZQRv6LcYR6zZ2CzYUQay
XF+viJUkdRv/QWVT7r+0rufy8P04H81Hl7Nsls/d0RzH9+nytV+2jyb5AQ3ybR2V
gkRcbUNTRm47ffeOEMuYQM/B5krHMBSGnsae7x84e4YJDX3rCzuQaUEeWqc0paMO
0/QyRLF8VZZvmXXekszpokvEwcReUQmAXITwjHrCtR0Jvmts1lm154xQzSmylNiJ
yEwDM9Hy0GWXSs0hEPJt0gXuDpsz1IsAWjP5v38OKYshic+JaoFM6Y5WbEBV3CEB
4OQUpkSva2IB65DRA5I2DI1uFHZiYvKHAs6f9rTj9d7YPggDC6ryQWRKXSmialew
Nr4Oej2r75aBgKz++mcc5uvzKlZMuhwacOkqopVFtPpNudLeG29y56tWmgmoEWf4
bBYPekNMzdJ7BnrUozc8SITxrYFnADdMLbAmiJgO1f7EhxrY1yMReqpoyjk25rQA
OJFhY+Rf7vm9PooqTGb7L8dt7Tcb9P3ZkrGhnWEK6uXMs5G2swSpPemUSwlvTQiW
ul2SA8QTC525laETqfHJbWSVBlZA0utub9rv+Vls9Ztez8peh1oQMeSph6yZsaol
ulUUlIYC8loUFwh5CgNZQQmZXb+vObzwornbgntwaMb1hBKogFBAOmS/N39270x0
w3DDvk9cCqppV4CWdwPyXFGXWnPiQR1FYVWWvLriRsB+qoDbL6X3q5WxYgHTaixk
PTheqBd6MA9iMPt4JntGIVQSQ21rH8oxaMDJOq2qWaO0Sg1GQifM8RXQMe+VhWeB
L7q3r9vFO4uEtVtvsSLBV10HBWe0L7akeX40pDSy8aV+/Q5XUojrorF+PmGljriO
fopVQPeMgogCl0CV7LujOt4ToQnck2avOA/hE0NqCHCo8Zq5D2FfQQYWJLLBStHt
v5Zi5d+l662TlLN0IQRPCSyUfY3nj5P2ty4x5S+wrIo4vs+wHTQzqAJ6jd6wu7T7
miv77ceQ+weAQ+9ZyVjr0CmfqB8MfSLoTQpTfme0QW/mTYI8CRTHbMNEWv9oGKo6
bglw8pp4Pg/FKo9zJDTAFGti8xfcJEGS9C0iqflccWoIT/SJAjHDWJvXxCCG5BDE
3P8uLEmJxo1BSIygm9Sqk/opFfclznJkoY2oICvZUZ+Mh6XS245EJqudHS/LN4pn
0zeCSjoh5MoH7Eul+U60zpU5GYlp5t1L3pGuAMqbOUoW8pC5dbI+pXcBRJb8lHJC
DsLBKirT0+Kv+/qI/CsrYGDpq54SXPxcXDyXxieYWWCJXmWC+bux7dbVuIQBAOt3
wTsf4t7U4PrymIbEofdQ/jdZD2BkoksTmHiGBsdnDAxdlwJopXnU950B26FmmEKA
xcxLnDqtv+M8JIWRAyOFkQVDNMKKIaq8Hdx5HKPsJUTl5KHIav9khBu2+b/EO+HD
ug3gi5wN7RWLTm8fhY8YQYzlUA0AI19EkRZicIXjJ21b1cVKzSJVcDm0+k1dq1To
mVunA8KFw0XDTbqv+LevMOokDvZ2FUI4gwciMlt+YxTUa5hhpMxSAQY1RccJCLEn
N414vSyky7IPvIdtoErNE1DBXvEnHcPbm/5LQxetgoky5SoSWsfbs2SXRgtEhJRA
VItEQ0ZjLsH7NzRi+rU7s08nog/lQH9xjdinz/b65LtkHj2ittTaGWEpOYAG2Bhz
p8scwQhO2uJg0ruV9t80NY2glwTj0EWmktKkEoP3o70r4CjsH6wxi57gI/4i07Ks
IcOk4Nc05vQ81tv0v9UYpKJlAFoE3KyRF4dVEt6ToIJOfVuFei5c/GArDbQZ5UgT
5Nbjy8mEJMKjlhThxXbpqzudEAapde6K2RPEA3IBZvT2pyOpe3rwrz4myGJuoeuU
9HjlUz0eex9ra4gAI6d2ru5mw6rqnH//U8JyeJ7Sq5ARhhOQgE3Zj9Dga3MbD6gg
ojdd2FJtm5+xyAAmg0A6SnXbRhZgPhhne19z26a8RNYV3QER0tpkXTXRQii3LNSF
heUz7S8e3KmgmEVDoyXlIWAqpFzKOnwrMoH+rKNNGcoKoXDyV9PsMAHomWztArsX
qweyTUZ1XEcek45OsE3ri0eiEE7nGOV7IhI7I6CAqwSHvYbeeJUtCvb6XTTFukpO
ixKxStY4VjNRVtW6nMhjP+UzusQXptxr/CMHwZy8AjjV8hDoxtumSGFuWXzYbGw+
xrNutwZCxyOMrDxnm8TfMFLUUVRhcHKz5bUAaZM3jxEHDNeX5AL8oR6qOud4NN/4
HEM5PXhctUfpPVzUoUKJgebXoocbkZ9vM0UW+WgGkv+XWFRMNy2ScQWGn0pIsOy9
dqkQevNzJeQwGaHROl8QOoaoRV5TgWJIa/xKX21MXVYUAzxZNQctntNbG/UoRuQ/
2BxUIXAlDbhk9oVjylmByQM9f6yPKIhf8jAvguYJ23kjXsw0WX1kU8oofdvdsF49
TohBzU14f7ZNXYGx6ZgcYSQpLRXJKaiOZhCf+OUUSPqM2yTq818l0VhnEObRgaki
qpBaHcMXzm9mg282JwOxdoudxAv5xuv0p36zSe888f5LlICU4ci/JyQwNjLpCRow
5wL9wMc88Lda95swY836x6hlY8qghmlndGcozzqiYkChHtzMVIJXA9gzky69p/Zs
Z1khz9kWQjic3kVgCLoKYbSghee+g9kdsBcpTsnvbSPhm4Xkmaqm4lejHcSklG+5
WyZEpK5GKS+Xl5pszIV336v6N38KNbrKEg5vlNfPsl+Gko/H0THi/DnyzMYNSzsK
XQR7QgN9Li7aelnjZvsSYsRDm3exA0dEHfu0+xmTvZjIOE6mcPdYbT8DPBMkxUGP
Cv1XtSfKNTgrhfIugcJDLCRrtwPJ76bKIcCFnj/Y33OWcjc0da53KIsWrOua9qrW
rKOGtlWYwHjXLDCphbBhooGzICQZz/qFqxMet8R9lE7YynHfVLx5LvLLHV4BgfBJ
qu8ekjo40ozGNJRG5HbT4tylYHg02uVpDrC4DN2TF6YMzEOrNe9zqdxmRtsIrspi
dqPzHfPOtUrvC1UCtxp/GFMpIrlB6nz4QbcFdeLAY2reu6n1S+O+CfpBgjmMlx1e
Se0O1jYOJZXQ7CH1u8/R6qkkKuMWvu7eDauWTu7d1m/HkNrE778aLefMlL8Y+anc
aps322Uvz8W2fYDzh31kaFHLC3dnah01NlYgRyhUrJ5rXAPsGctB9v6wIRTClsC0
K4TnQ+3Px+UCmR61K/ASf/jNeP2278KlcSqO/VQn38B8bKfrAU5utBO9tPUby7cw
/nH5ln9kry5QscWfPCJMSTaSTezjb1uGWEAHNxVmgMSyU62w9f5sPoRMZWR6TuTF
cuQSyKsq6g3zTjs4Jv5dUhnCYUTDFCbnKhTx9eR3IR8AEERujTYn0xi1bzQsirN6
74Ue6o2Izg/olLKx0t6gHP7l3kvuC3rSP6K1bcsCrIcruZJaFmttWy9saj/jPcyc
LbdpsHVMAAyEAqyz2veNQO75PzBn3NBWVjANJWd4i1StpyriPwyugJjK2Y5A1g8m
X3TqvRqs2unaqPsOFCZtoYaZpaHMymis7/K2jblcunatrQ4BeDXIomInqz+0jvT/
bu/8JKP7EiXJLzILoFK10vd7L4266qCLazo3FhkHL3ZxRHys01i/fH7cpa6YRUwS
q3oG5qCNDey9Veu/5xSEzV20aerBIEa366lRyCcKZXiELdX3wVG16nKG3YzEIW0c
g1NN6ouG0hZnPZDZBNT8Aa6HL+363ZTufsh6ccvCYOUlwqtSPhH5iHI5YoACusEi
iboxNr40TzWvbCOhjWhI3ycLEX6ng2EX1U7NQtSoeffaCSmyGwyRu38T3fWb72ul
kEqJZ6ZMlbQQJqaP0ErxDCJh6gtoFFOxuGDVG0jqMehrbMCOopoW91YcLa0W0aO7
6EH7XzF0H5yd5VdFiDNIbwTXrqbJl66B8kgVaTCcpdE5ATPNV3/ZQXJhQal0bqeW
d70UB1Hu/+Ru6GeS59YfHJb8gjStFZiuinMOAC7Z3fscYGSAuUI/aavZZFq0uhig
ZDSo4rShUIDE3bt8Awe6iEIHy4YHSCc+MYAFXwFpfi2pmjVT2ajj0EDegeFUCAsl
rvCwC7X8bUplIQsrGrXaR1WBWVQuzNJE/zle16lLCyNHiIMUlxWS1xHoVNuzXprS
WoGDBNow6JlaQcVwmRMvemlKpJRHOq+LMbabcB3SXH6Z1xhHRTZcwaWT6H/TrJ4i
J526gLjhGrsmLM2+xay4jQiV4j96TbxnsviVaQuP+G4TfagTiZRnU7y45Utewy8m
Y7ahWEIgzWEYx1J9qsw8XubE85p/q2OeieYdrALeC0vVecyW/RqSJwVrkivnQCg4
S73TsjLQfX6b0AcKyNoo0YAoGF2pZN+W8WWTKRuRRMswClKp6YXZo4RoAdlEY5rf
i6JUomZoJKtuvmvpvUkNsAi1K8fgrjASqk7dnlE+zQde2wJiejbSY9Gtjj1GnttY
sXSUOJHPKm5jQOuMl7BtWl8/JuOOrnq5RDQZXuAsTjdSIJzhLRnLUa8gSK+/Vv/8
pGVVFA62LM/riPKSm8jsDfgoDhLG451mEJzPxepiQ+bXTt3fzP1xJVsPuIImxP/J
bery1ELYODshdBcwpmCUVcF/TXRHLibOnCcFTSS9GLI8FlmM+8UtunwGDYDY/EIR
Lxxc/8UAIU+EMCxf4DVgstggkj37E17rFxUuglYvfeHR1b899NJMjnfbVbmx5Pkx
Tt0EseuQ3SWJ81yUPBqKVKI8BOMdhmNg2l8BhKasrjgbTRIGinXel2SxqQg20yRQ
jMA8yIoXIXcruw7tT4hENlfcISWj/G/ZeNwUpCxh6BRPQ5ljn6gezKoID7JaguGd
L/WBNuoWNeszDxcs6Z7CysLyBYjhO8EDY9Oxj8EM1lLv8oYtMBieo+WWiGVAaohg
n/TYUEq+FRLMVhAknRw/R6GX5kjAWD6SMEHr2xAF8wgRY7VNGcv270RelmnnQBE8
1JVpULXAsiAxL5/71j30ir5gGL1XWql7Hag8/uNmzxxxhefc/Yg0bAx2NsUBQfAm
8A5eq5CLm0StiW1WZPtg5aJm2QDHNB/XpwtQrXYV+zre/oWHdQbzsSJRQXgkk02L
Ici6pdVVRqy9E32TcLr6RiRNPI60A0AAhLIWr7Y099oPXvR+xQyqHr71ic/8Kq9t
qTB2urXilkjAkvDChPLelRDlBVHdrsYCVGdAnpkulgcslNrIppMWvmMkYLi9SivS
+uul5mzBY82W6tuv3QNB8risV8gLCOciiMxlUXogGkHSP+y0f3bnnSskChBigJwV
owEiIOi2eQMX8UHi1pxXnYSAhLsn+tCmcYtX2tW+eufSd+IyuKT18u2U0Dq49ts6
6TC9FrFYqIzaOj/E4OghxSY3HnN83l/LPkgWPJTesvORlI3yu/lhoYMZUs0+eJtM
07xPsJqbu/Bil/15dRBeTLguNZNX8d5yG4V1a/hKdnNqinLG8qZDVDngPSdErhaG
6CbN+stM68YlyRcgjK/Nde1nctmm3q5nnEIHWsBb+LsOOwkVgLmJ/Ar6f/dPsMTe
4NED7pFVflS9pfJm559Mce2c/8XhecuM0B5aFZlc9j1BklLXhPt7BmdJUTrgGkP5
K3jwti/ly7wNq2QWORtX/hCanDkmuHAkCDFfP/XVeCwAIKpdDFEba2GHvnj24SZs
lWskygNomaDQJVm3mKVxYRkZrk1CE0WoOocKhyhq77KpYYLx8ZJaYq3o6f9u7PVO
gG/91zZbc5TlrVZScaojEKm0UCdG6ilKy8SZIsrBiqMLcma4yseX8EnKZ90ZQPZp
Yy9o2PGZJ80y2ba+j3hE7p6aZyZgS67nOYaoGi3gQOyuqQleqVYhTZydyX3dMlBq
8v7RVfB7lc3sT8ZyZHWBLMYGiSEsg0weERckV8rK2+Enf7jx7XjWH7q81ANi0bQF
Pla5ZTlfR1QDl1EHPEtXXjUjizlnr5qA3yOWa+oU64cSzehDP+QkP1LaO2SUyDoC
9bwDcK+jqBvKoCmV1RATnmQHIfijVqenmJITwvBuWFF4U2zXqYiY5GVz3ZxVd+p/
FFY0wWsFnDD39nJ/miliilqrOoKyMJSpIKERt3xFBBk2GFAUVS5czujIqxPSJHvN
f8NVznkJyvGN+W5l35tvC7jJk+fIt2qHiJnlmUa/raqXs5WwG/1zeu5oaK14dwd9
bfreOZICOMBAj3e+cP1me8hBzXHtJTEeC26LeR+UuK8CYzpHE9lKh+CBNaUKabYK
xZ67K2pWlzlFHsp9DVpslJ5c3SYc4g7vKxleQ2cwWIHhEkRfhGGtMWe4kHzd+AB0
u2pR2h1Ha5yVECqwYdkj47f/jyM0SgxSdJ7cNT9CUQwMNBupfDjVpadCPzp9FKsp
v23d3IhEI7df3dX/ONfe7Okj7QdSjG3gv8tHeLURk3WBocKDyAwo7nGvkTFTRiPJ
SZv01Zv+BZp+giVeXL7PqlHhD4OU/I3xahK4mNJ8NkXHk3guKynhqoco5GpeUTlv
fHflWvxb54ycDehNnuMGJ3uoQVXhJFjYYuGZS4r70WgjiBH5pXS3BErMSnHVAP+v
Aa1t9KQTK7W3KF3WDSe+ih/hDpukobKCoZGfV3o5m6Aur2ZQlBEiVlpgEw8YvT2r
AWt5JIVUhFN1xjO+sDNDtnc/Sx/Qmp1jZe24dAh0XL191msHIl8CvEnXwkuJXOdD
aX2nCqduEOlg7aHK++EW2jJMAe6r440yblXEkaql9ElG4OShbV09w3D8hourDceu
60p0vLPt5w8nphaefQ5mKdbx5Jtrp4OunnIZ8VW4QNrcmZlJb/NemCsA1Yshd+qe
qxsyp0Hsb25ISe1iKqTMp0TKVO8UBar1AkcMasSiw8VSxqBcwJgMeOPSsm93WOOr
bMuUpsAqHXiJkjHJzX4FkQo+MGVD7Q5GJu2Z0ykvFlSd3yAzdWgN+Pp77vmqXYKr
g2r7KzUIca7G5RS20yzMnZWr+ii1Fe8Z9kjmBbIJcEnyRIQ9fMyLI9aFqIM3W/v9
aOPh0g0BfLYxNG69v4IEFAAN93cly6KYHmxiZeVCmSC63e9A6H9Gny0m/PlrTxa6
mxbPqdE7BjV9UjwL//n5fWHEAaFhw96dD9SASKWYHHzSZI5fr+TfiYLFyC6jaqpA
lnm6j/U18fBevY9b6okqeRBZTfFvdeuK7syAG0Ko99c3betWCcFmnW0Eh+QxEBlV
vUOR6wT9p6zYS3QZkypFUkTCSxuYkLZIIWXItSczzxwZBkk+ZIHuuKu/cY8jtqKT
qLzyANDeFJ1QR6iVMtxsQQ4uu0v5fKvxxOlLTs/BmnXOajk7vPCVIMglJE/NXKi6
3kqYysRj8faqUFgzYtiM54H8IdefJ++hymVQ7wvMg00xQ1ftkpkIDpRXAvkIS8YS
Dhgatohnyb/c1f7NKTInCBjgvwCDDVpb7WA9QqXL76UWQqVIinvakPFwAtMTVoWn
5FjkMzZn4QLaU4fpVcQiATF+iefDotOJSb/WaIen5nt8Ews1xUoYS+SEDRVdGcDj
rGdHEELE3hjmYkJ9kSezo0HfNDGCQya0Cqj1Wa6wJanUk5gZicDSYh4Zxf51qjP4
Xm6fFi+K+7wlxxx9UOl2z/RksgCyJL7Y3NIZWOoWsmn7A1w54yDBaR2MEmVhpy85
Hf9+9Vq6qaiY2ZjLhYGbBO2vZX92YXcZp0o1oAYFrYW1vjphJPqE1JFGKKuyUrAI
U9Urmiun95sCKW3EvXNlFcN1PP4QkY1cWzXTfHDlvpe+9gZCaTyzIj1QnzQxtuoX
rnANrJYCcGyf8eaKcuFvNNNc8MG3AmTGpljIgC+N8OtDlKYhFs7o3BOwy7w10W8O
CuBVES/Oj8wVRA46eX4yuVALIRUZg6Km5yhn/5Bh/9HufmlGk1a1+hewoO0rF2FW
8I5bTTNujdUROtSlGm4nPYDA5G6mVYQfK5q53Msmz8vLKDEjslv2blI3XKc7vp6H
nlDQpyIWKK/QNPLiEQY2Stm0/fAMlC/jJQvQ0AAqsQUEcBUEOs+95TVkWy0HSohY
emmSB9LbQr2UKVhACMNS5fzr5LTnuNS63c9HPfztb/nhF6587Ns20E8eetKaqM5o
4BeeGF/8hGTVtNaxB1gqbsuQINJysJEX628Mwgpq/TdtNgoMSckaaOtfdESKbfBq
rSfhPoEbR42ZRA6o4FcclsFjc/PsWKNzuR69qx7uhwtbQ8QM+aPgcNtaaxxpr65T
yOtx0T+bgJqOYPqrJHcrQi3pCuXMhzDjyUoXY03a3OUEki42fGffFYeeu6x6HmPD
9dN5QQcb+gdAHKym6dom0aht21ZVkWimO4VlMrCr6Hanvk/Zc12zZS5pVb/0E5eN
pXpP1jtcZxn3wWcY+HtsD0EjwvqLYYQF/eW48dmGyOeASzZct1dRsO4YqvjgdAk4
Kui7QAxzbk7v2ceNEdaqZGnWWZ1lBpeFsmQwAb5nRYGwGPyj94beLmVhsyHBY9WQ
LykBhvVfrgjBRUIDXLGCy9WgQjfl7d2PhXk2tTuoIkXws4CouZvAHMU/UMWrvmE6
T/BGt06Hx2S0EvEp8E4PtWbLQ4x7/gku0SQICm6XX+mdAeuzmP7iJ3yyPdnkrgx5
95+7HXwa967F8/SJF5kaDtRrEoDK7JnRmP2Wafc3t4hTiQ+B9CU16SWe84Jmpsac
tDIWO8855W0xxmpIv2M3QlFqdUHRdC15Td6KZZmBHLSbc5JN41m/yuTB4y25zo2M
WbXoNuhxbZfgWykGoEoZQxkE4VTI7zxeQcscqEGDxxm+lgWmQSsUpHylewrTr2VD
bib44tzVNl8R8JVl9awWisbAqhpUxbDvDWr400k7QauwMl9xGyvtOtRS1aN8s20G
7pY/lKY+7Bllx0Z1Kytur7vpZ94/RAewmSlG1dTr7d9XguJVpUTUBt1c8FuvvE65
Guranm0NUV3kgeWZHcz9ZRkZucT1Jwy1EN7llsY+76NphHmqpr91gHG++vkKVVjG
8QG0ZMTq6Z5CZppx3L+f+17KbgbFPXDYVBTwH+78g1QFo2cdJHeNbp8x8H+RHijp
Y0XweVU9RWB+hga4ZNZYTVHprFt80af+9BvuYBwNMDLKGw4QGvERgSC1imAPhnoU
kl/ipPFuvIkkwAfcmJQp2jT1TEjuyHzR1+99TzcLcRj4rfsjlXkTILV00BCokhog
V1rxWEd32egmlckz+dfVCrvd+zfLa/MfLyyMkWH0UwjsvDvttt20vkG62gOqD4re
TCa7NYmkSD/Y7ebQQHlaEBlWAzoRTvYNsxF/evK0DLyaNcll17eFLKdmS4PJ++VX
PcFBLz+C8bzAk3o5vxCDiCzQMnWrnSS18hSZQ8bM/OhacHHsH0oxO2Yeg/2hZ4ln
Nno1ebupmPdlf2KwLNSEPhjkgXy9gTdke1/rJslmFV3Tr4tGE498MlXRgj3//qmA
3qbsFKCjlhbV7VE/KGBX0CTvqHSSdkf7m2YOMvlI0cO5duK+wmAri6XiZncyYhsu
C4KEPZz0ndFxbZ5uwSSYjmvWS6rlqZkCRp85rCsIieDpzUS9Gg7IqmG5N4GxF50O
dYAaXeOe5c4TEU58NfUQTxIMPwdhiF5rYyFSEzhyD0yOYXFN7nZ41DSyQIhE19dU
2Di1PudDGzIlzreQktFyrHvnIiQzDGQlbg1B9ZZ7tRx2qPwmlRrESTC94VAu2NCS
fh0dXn3nC2OFrKRU5Z6s/dY1dsL3dr4Z/iFArVKhrgWR9wPK/kDJQT72FUefF2gu
1Pn6L1Q4YHhBWHJQln9/cvMobJ1vyMYrcfaJM+fJoRvDu+wPcHcVMGviT7IaeTYT
WoXDpdeOLfHYZiCUSUOZa42Gxf17EKl6q2rB6nNawgqGZ1g9GWUZvguhkiFjmeDH
xe7KmkpJHuP4u+YNYtIeIws/aNKtMrR+dcfg1S+w/VKJxjkwkd0DpDbnGfs+aRIZ
ZaUOzn77+d/12Bd0fTcQyO8l0/Ywhc1goLRfwi4mNtiy3qp9wxtziIzkKdzFZGHT
m/HhdCfcWFtwlyocE9ChXf60ACk6dEqTtuFeERL8WwjsAgAFEHuPeatJ+yOeuzMc
ypaJr+pEogUW34QLiYDstxNB5pm2IwCAgCzyr8mKob1J51uYo/LG8EpfIfb4LpoJ
sloYfXlJym2aIVSVTS/5tS64TMSka6cf+H6aXdnDSLsSUs/UHmrNUyfos5fuX14/
W+46pZKo/eg7tIfJDbshPeNIMl2Vk5sr04rLHzA4vyecnGmM4QigaZ3TUDX1LHux
yu5LilWKuz2ahC79EX9AEtqYCgVTIxyyjj0lW0l86Lk=
`protect END_PROTECTED
