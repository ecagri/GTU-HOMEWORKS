`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TL3DC7D8QbX7RJr3g8MOt9avN4ZZPLRh6YA82MuU9izoWoRrHnTRWb7CgYbf6Pf3
T9Uav8y+Cr+P17e/CRen6e76CZE5lgETLgTIwJvVPdbcZTBog4Stw36hCggoODmU
sRX4oTLCAZE8reJi+24PYdze3fywQaCwHIzVt6LHP2fWPk99LXrWeWgoT8LtdfXa
kM6wFRVQDkhq5WHaGmzZe/8SmgqZczHJzgSRP/43d0r2w48TdfmnTWDh3zGWOhsU
AbuarRyyQxnzryEe8vxJx9/UtuVvRtxgRhx979yL2632INFny8a6EUL3fj+/tURH
ePUNto/LIj5Pm3YJhPVBF7BO/MyIn28a93q8ujeJWRl8X4MMIsY+kFATwgMhFCJj
Sz8pT6xvk+jKSfrUQJF6SMmdOBhL6Wif2F6MYPTKNqdIRv7Z0wdhlaHGJcnuSO8h
PCp5mqH/gu2pQ5m8Nh8ZAFzI6aavNELwsSpw3AA8ABzzfEpqp5Q5naRCFidz4pyZ
15bi86UbPyrEmmJ3e4GIeK9fA6YDmLkINbwuzqBGYG29RJjHrCMtBgEGrzDZLPub
ERRnIfpvfvgA/igBztCLWsG3F6CIHP/RN/5RFaodYisCnRwyokqMHuyqSIT9Becj
jE2eQ0ro27Eb32phdxkKqV5v1A0CoIuc2fdz8wnRxdDkejWv5VK64B64+UdxjJaC
QWKErgnBYbqrvYUb9MNp1UpYY4jEpJDV7rEgcGLk4CpJfvHr9fRZDMPwMlgiwlJv
un7YiEhL+tdnaGpNdrq+X3tl/2bndUXXYiBnYfuTfmLCBNVum6wpjwZGmOW+IqhA
/GIbjyRMYncS0fUak1hq8V4P7G7xpcAWGfGSVqRS/Flc/Hm8iPvFX4X5+d3bRPPO
LHCXknrV4o8LOyUmZLfDdScBJOKPCFcujS4mojB8zN0JqeiciyuyMITLZRLxZ/Sj
DWbNrHc9uq5Wz3EnQOwErhQhcbQfTTDPVAY8Q1caZlfskeaP/Vax8DNGtXNR7cj7
WTofsWuAre4onphwogx+QZ1akLr4yGES149lsgp8x4/hc29UJ0NMwscLRjicJuAA
`protect END_PROTECTED
