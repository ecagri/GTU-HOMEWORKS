`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mg9WDz3oWWnejZZ3/XFdq/KyTTvzoNg3vNqSI2DP9K+ObzKfgWz/4FNCdVHGinWA
FwHwXVvq/MZNlSmhMwNqXyIU7qgcws4wItqbPm69vFWVKu4bjO7cWji7job/cKhd
QEyWrhBsuV0cWy+rmIfWvrXG5+Y2icew7EnHxVsc+de9h8RbLLOFNws6wLOa7sEq
nY7A/Ekrlhabj8hYQ6qyHm0wvIt2OiEhi0jQCkXV6kCoFzfFm8aGjeiUPajNZW4v
lMnF4NXepCYvQXBi/J0FEDMwnWFPJm/ldXC9kVVXWPl2HT6ZYzmLUas7epmTW3i7
olyYmdW2DBeGrRf428NQzK5oo3FxkuoRhWpVhQPLcCt2S5xOP1k6xi8aUQJD5H9R
JtIZnaJAFkPPT+BPD8r3sKOdvjOKC6IjZJ7NTB7NhuDsq/PXkdptAxjvxwxRBYAb
w33CBVvlNcIDAiV4Jq7ut81SCeC2aWMAnLLygX5l6I6Xrjf075Zy+MQdxQFg4wmD
n3T2LDBezvpcJ4wnykmY8XvOb/MFtNoe786QyXUVvwCP2ja5q9vtVs/YSw9O+43K
a+pSZxnVQkIDMnMIeTyaDLOMeWA+zqMSzyxvpA+AKb4kWfTzgb2lNL0JemwCqqhF
H0gYPnHO+Z8K2okEz3lW9e7D+11N43Mtn8L1QR9VbTUYO03Pw3JuBpq3sDgLsdBz
mevR1049onXocbJDVqeHtUdtWslAekpvoiZzsUllOneiGt6l/LN+adOKo9Zun4B7
LVLXZMKVz4E8Ao11pJN1dB7DAF95Sg4jLoRza2Jv3Qg4JdMQPmW96UzJFFIC7sxJ
Jg4Ui/4PclQ8CD+8RpHsmn9bknp3NzLxz5Xr/jSLtuztYT46jOH7MV4AGJk+xQfP
sCtbr20rKIRoUiipWVf5WT6fZSvb6dZ7cG5YtD2GRNhC/VY9n9YyUonOjkGMwNf0
Xc2VfIjcHtpdiHfy87rN/8Y4axZTTBC7Fc++zxrHx30jlFdDrtFHGhOBL0lcm1ID
CLCADLYlKnKCCFMWMFB6Tu9OLiFsMvbGl4/zxelfUR9TkGl/OiAqwUrTHYhsMQLL
+/2/9Mqai/BSJfUWLlyOHFqanOEjkKlqPpQ1vNqK0a6Tnh7hY0xNT0NxOFmnen0e
HOmoqnNL5Taeu1J7mkOxDRzruEMIkF4WiCw80QkZIoCmSDoOWUJ2mLKtEgsU/ld4
lNYCXLdZ82uTQKgwUFeCa8susNWAMZ1eoBbQ2DRbJ9PaI70HXsSuCLk3HPPr5wLO
YfTNumOQ9GbbTUbkKKCE8BeatRbKXlr7f3XeUAu1P14nCVhak+18wUfGmXtOIQ46
o4lVfa9DZ4pGFlBaKru0V/1RKjPyOkIJFmXxZ9S8oOPs8ISnF/27y94ONMg+YYqF
wlmeboM/NQ5k/RsSUDdgV3/WviTkoxDle5RyCbhiMVOBEmaghUXn5feBmsDP1kwD
ZMAIrqIrdBZZzHkrqBJ3dPJSJlyhak7OZePBXGhMkrvReHOWpIZG+hFhXt+L/NPW
4atXWx1bt5AfRb9fp6EUw0Eh0B8qI4Mx+YolhVf/qAlimA/I17TAwRsy39oqF4tw
Bc3hzJgBLP9mayQ158hjhR1JrSatxRYmqTmRpTqJSOQltH9iU7fboLOkpKMKxw8w
`protect END_PROTECTED
