`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ek64CNjtz/HRUIDbiCcvXbJB+nGfti1JzQX3a7V8c8OVSbH7QqFqJwkERmmwutXI
L8SYRv1Sy3aoXco4oYsBaDHut1HDCq9VcDvzWoIozT/ksJ0y3q4KbAcBTQa8eQSU
nc7G6bqIuoz8fuAEY/ZMf50Kw2CqMibwOVfWqVMbV7v0oOZj+0iAL6duasZ8lAB1
PtXTKgZW+myUe/wDrQm1h6DNqXRARfTgvngoejK3xlTSEBHqG8JiRyfXTG23Z/0j
COkfh2jgspQAwbt+3iwy//mit2GMnQ9d1LJ2GXjlpuIPO5qqrNWYVoEgYz10MmHQ
KFWG5WtdE/3WotKWa7p+6H9oZu93PnyHZKZ5uh9cojO/1MxOVHNlt8DPbXEG2yF8
PD867Ob8xMvq9kyxHhR57VPsgvXR7mg9Abdif21WTfkpMXQ/+02mVSpxmLbiZhp0
9fCHbqs2DxfXLueshaz8P5Out56YkIgUshz3/a5J0Si3erHc7FZwrFiP0/DYNOnI
XxDkG1ToMaZ1P2nNI5njX0vqhJiSWQYwLZ0YnUuTZm2gw1FCQLLFPcXMAtPPd0Zv
NBiE+Nt5uaNfM4UgB4DYv1DLhBNDrLQ2VNfyzhljX5smGqIjYRYwGvYWA/tMYROB
LACwWSfIADLX2B0F1xy97aaHPJfUeo6bepWLB8uCVJ7G7Cwb8CXZ5ooS1cs1qeB9
o0y7ah8ay6S2m0Z2W0pAHaXbj0mPbQeKJhmFyVZqXdjvGUy3yCUpz4RdCegYXKJ4
3P8nrzQM83bECmQ/YXo/r7/jg45bHPYy36IOJ03WYMRSh8oxH47C1Y4dYPS0lTU2
TddyE0NDPCpcUVnPhaM/2AcqeDJdBMiYSD3IAePjKEOHoMEJPaKDjJf5XLw+lyr3
YZO57+UUnOJ9zdKnYwGjV5Ab1rwcUFf+tHLMOeI1/UTpluLfXEEvH/BGR9hlgB8X
DssT4rEAoxGODDE0Nmg69krufq/ch3fUZlWHyaxHcFUZQG0HyAAiSV8v7wmD70d8
NGmPm0SbJiMhrtPEFd3LzYLPGsTr9jtz0gK9SvSmMfvQCk+neQpjBVJlG3n/yxzr
kUSaNZm5beyKCDzMnFCFhnONpY/AuXeNTP9guiziZCx+GOOC70VgomB3irlcqyhT
0jJG+T9hxRdyVihBBUh+3hjsWWK2jVY+sIZ+9ZV/SFqd1wzFoW9GHu5x90ngrt+u
AFVrN2UKtQSgAjiBnLWhBBkbr39WF6csx79p3Y77lGh2hFeQnwLgtj1W/VUP0HPZ
VoIfXHkQSfKsfylCj4GPSroQpA3rgjOJRCnIPlOGkN1uBheXuYuT12l0HHfV6aqs
ga4woNgnvkZIeWGs5KiFT4A8OUO+lWofxv37cRxfPyXHrIg0YCMblcdR+hJ5d4V1
Gi5taUE4Tq9EztGZu6bznR8g/FwC96Fvso6mzBoii6mCYKNnuqBlu6x1hi/Zv/NF
b+YT4VcDTTxt0t1JZE/TtFJcc5DS2kC0747RLa7ijK17v8O00uRRLSLaVwZVnkjN
CdJBShyCSsloaLTJZ1PPJKr0oZfbt8fC79/SHbnsF03F4CEMv+XXN3jtA4Nhjwy0
LonSfXB+SzNyWZRSCe4QOjLnJKnlaSmz/DiwcBL+LkA=
`protect END_PROTECTED
