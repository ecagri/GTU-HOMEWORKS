`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gtHs4BnJH4PbnQy/edF/NFNKvXkFZT2hI6ujc4MfkACdoGxW41VhFoMhdPtXevLQ
jZEk4OI8TpXQyYv5Hk55a9p8CN6bN9yO3mhQRHRSNzSZ5N151Qgf7cl6dNbVOj8B
n4+NfLwrahfHvfSxY+vuYh7ReP1rp6xmUUZ2kx8re3biFM1N9f2dveC5p5HVqGBT
vuwigMvPb07fWg/KPVj8WiLn8V3AS8tSI9eGmPugI/PnEKrH884wuFFuc/gDTaRd
/AQN8KQf13jKXJmXDZCicg==
`protect END_PROTECTED
