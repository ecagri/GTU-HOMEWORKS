`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ekWJ1nRGuR0ePN414YpEJM4UwAqp7ZAKtVaexsgaWUTOdXd69rh5yvLWnT60l5HH
0qGtPkdzbYSss7+T9E93SqJE25tXz6BPqOyQTEJmaQO2s7GdT6WkxAfra4LDr3WO
AwWZf3BOIOf6dS7gzN/zIhDZC7E5LQgDWH0ckxj/3hlOU32NEbbUoGvPAYAO1JGo
4JjRWYV/WcTofn9NBxFZUSBzJWY8ODkVrCGZglGTmzWl+8uvpgNQwgQNoXk+lHWp
TluQpuWqrmu+pGOyVwww8pIwAIbWkKBgE1zzJimJYe0NwQx3S19L0aytkn3NYhER
//PSy1CyPvDIQNWHBj2jjrfUBxJ8wox6QfELhaTlYnbrGde4hlAV1bAoIz3RGW7r
7ndLNUhcOX6c9eRWoLkxL9hJ4avu+GNd4SV9Vfk5+5bQsKZx7XKfb8KLlk0NFCDR
7TX1iK78IS8YwLHOQtCEGJw8JklDDK/QTMngQ9jkQXiendLp3TdoeLBiTXykyiUK
sdM/dXV6qI/zz46Ib2qaMOdmNv1j1LxFypaWXeCBWE95WTddAlv3dk+HMgIL3xg1
CF6aALWFYXHZYOSX1WJKbf7uUl/wNmQ5czXaxjwBCIMfEQYfe1VQBmDo6UL6U1o4
P3Xjm3p4xCJ9RBIG4dzBJVPa12CYr8TxLFTxIXTLDDBTRnF92q219O4mrpXvJG0o
s5pr1I4ZXneJU7HpNYnvnAK7MofbK6asG1O9Mbsb9ysvp9xzfOtcoofseVRtfSIO
KfxAbaU9LWwh81agwXMYvg==
`protect END_PROTECTED
