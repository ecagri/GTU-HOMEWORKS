`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b2R27QLeLH1NDo1wTR/q21mvoSclO7Myun4QbkQ8A478zH67vFAyGeU3GA2mVUjY
HNkWsOx35+Rdo7WJ8JRmlbHgGFtYM6y+5ub0VfAGkxGX6Xul0Ezny5E2kb0NISzO
mE05GSahPvLkBZff8ll6Z40WFh/l4MpDv4hf+BoBs8hVVJFB9HAeP4jDUmfaBjcV
nQicr0qYjCkgQEs7R9mtCrleVC9yGqYuYF7DjqYtZpvedM7VXEtpydmKdYuhOcp1
zSJ/o05SL9/YMBeO09kijYOaNJ+iMAxjoC4+7b1k4wAFSvrSoNM3t+PuuBWE197I
zAeD3KjHSyujDVRnVqUhBCibhPFy8uMm+7UHP3rKrMuYnqDS3NO49ddiSECQDQCn
5zxU3DPQYOYIm+pEwxWj6wU93u2zWLLgJo/RrH7O8YEGig/2Q/i3CikMEWfcnmrO
K0WzZnLGGcWO1cSQvU4/lES4kjfZAQRDxMHwKuytTuE=
`protect END_PROTECTED
