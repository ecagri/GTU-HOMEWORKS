`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zE5vzJZtoXb35rk1gcjwSd/1ufQAGT08okoqJBExOBDZKVVuWaaaBKvf44qk1Lur
ie3eQ5EVvt79U/EXGcOIwLZwTswLSGTW9uRqgmiVPIR5ZiXV4ZWtGTCCsSBYyhgs
cv9jl8a9SEBAJa4XpwSuWHYlcvxTeRqn/jPiw5SHif71kSZYHK50uRMHXbZ/sl7v
FbjstF6rzXffQMHDkBnwFbiLWSON7qLiwZcKkTIinjf/45qyJoWbhVlwdK777wkY
4bkqRm+aYYfU7jd8zuKwKtBOXtty8j9nlGYlAn/NfMrnI+IYa1a+hk2MvSLs6CL+
V/RBhmojkJaAivEu1nn4cFcU+At2oIyOOZRm04AvmuD09op4FZZd1c72QksuTeNz
zkqLPZGs8iO5VjA8v3rg501mu+h/0u9Wu4oyKSMHE/PhiTIXJ6RclMn/wYHqvy5E
4GDeREHHQ/2MS085GKObnGu2fzoQp3h/ItdN8CMNUJ1jo2zDfTE4Yy1Z58zLE7CG
dlA0XF0x3hO4/4dQDb0IzgtMbg9EMFKARXtYDapCIVPdwIUa6qzgjj73aleGTg5h
3KopBIlgylimtcOOEwGyb6kOb/6zGaqxxbD7DskPjBADwrOeiE40U1iQCgRIxJZF
VCmUQQ/qxP00E9T9KaEPaqsawFShqOjrqt6zp2nhTLIeJCVs/m9rC9vS2k8Fx+S+
20/gBFe3VCP8aIcfmpFwSBjD1y37/SD1g29/XRObrCVnvYeISeKWCUopVv70DPSV
a7sZ9HsMjzX6FUWAoAjDsGa4TdDmeNmNiwCK6dXZyaEts3pNjofbJFEg01qzmZpE
25A/aGD31836mkue2rvxN7u19ophqLLZNrIq4vmcJsePEJKBei3z1LPpFNRW5HNo
txMAN7G8dS6EqwhXIrUE6uKf+PliFmyUJwipPGSIGrYt3Mnr+seS4FrzjAMkKUSi
3zw4s2XGfE63tWcCWsJpVvlOyuhNieRQC7OJBmUda9O78wBXOMnagofbPYXpAErV
KN/2yof2qoKSoy4eWBxjMKlDH34GHyMjTnuwB0DD1y58sFW0/1a2UVZXwmllGAHO
pCIzM9kxiTUaB9/FUUH/aFnuSoIEPRpxdGAVKFG/8Oo5/zWHyW80sZ5P/cBaQF7/
1cJOs70qJL0hepxi5IdrBaHfFSHJfAY1wcDuyl3oZ0WO9l/37pzKfoXjqTUCO2mE
QmN5PkGCgs8FPOlrNAWi1K6Y/yl/51lCAk37oc/KasqCQTjLX33FRVjeiabQEOTY
kDelXjqKPmkIyr5UTyjbqkHeRhbkUbaK+tgRmxd1zIZ/IPmzCxAUgTiZX6sdsaGz
rj1wgkMjEQnj7odNzlOsRenaMvnu19uNesLTrNu/2SOAwQ1WhJU8S8LwtPkeqIrK
L3IVadb6ay9EnRkNRYNbtTZoGFKf48loarnMdnm2tsw0oOkrmCtYYA4gBbmyNpL6
O35xgooBM8+neFz1CGa02ALZeDLp1PIswAQkTJ5B6veErXLsoLh3R+uSgsZnnsmT
SLO7TAqVLpX3KXPv4ESqvmcKGnv3iA+Sfsr2gi8PDn2/vOaYH8OORmyo8kSob165
WnDHUwlyDPbQtyjeY4VomawT6d3ulHzON+5BRK1xdT9BfQ3CYSfBRrDPzab++FPj
bP0twEo6R01K/yRVWsXqYJNFou9P3n1aNNwaHjUmrXboBEVtsIfbTYjN7hWXNe9E
YtHkeE7cOK95gdwd8WiKoEXmUJPbm40q7t0KjSYeVauHXaLbAmd+OwVt7g0orV1h
akWJIRIX4rJI/9SQyNjdMnA97B9DDmDOzIowf8J7eV+KmqvsDb6z/8fhYI61gSca
gwzvT4WOuOUgeDZbeFAa3JdxHgYPO8nw5iB4RE5BRZQjY45414zDa80UQ6p56LjF
vZFmQ6Z1cFlP6ibvSX5jgWTtYMKiEWqofBrmhrmgh+7QnzLWKhDp2NvCGteZKLrY
HjysnAXL1/X7v5Hk/+EvO205/uRfiVuyw4vD3IlgIjoKpn5EabTUuyDe/kM1VW/E
Yd6cBllJOOIy72Ec8YVbomGhmWPyx//THMabn0rzPr9XTZlC54HE0YPXT4f4s9JG
cBol7waaPa1wh8o+UjeMBg64l98V75dFfBpTorr3yEa/vo3bDuU3X2yFZZTOao6N
2IiAKXZnW3r1Y3FcFGJGqd/aSsX7TF1Lc9HfkzfFgn5Jx+007URvyMvhHs5Qg7nw
ojK9l27jGk66SowN3Yo3aZMzg1fNrbXxwpFoFzI9FH6o5B2B2V3W/Kq0cYK5g2MK
002SShZ/gNAk3I9lTipckaQ1AaGyrqL9z+ye3dFFPDrjAfEVLAze18o/x2+G9Qe8
d2TxUTLYcIK2xTj1idjBq1YGuG6k/VU3KBFKm6JNH7QLemveOK+ClM9AFM67dfk6
9LXH8HLXyhFW6M4zFIo7+53+3DAusOoWGYWsLpqmuv7acI2EHOpudUSwzKZROxvV
GoAHDt+UPrKJT3U18+rMeYMqQ+5dNI9hc7dODr11HHmoWX0fWf1mz7ESkE0E31FW
lABxh/t0MqqkdkCuEvvYchPpBWazen+GZ229WnLFKXQ217JCjdNDFfaCIQku1Hg3
Ybdw98kPYUQwXtPLHoRTNcrolX27VzdMMYJsPzLfBVxLKPA/CxKA0v+UKfVlT3iP
8LW+SsLoYyfjs0iBK0FOejch8EqtE7tRyApOdO2+62M0tHajyoJWpr3No9I1MSVk
g5fGkw7KwiZMnV78thAbeZYFYbknFRAxKvne6KQk/VIbVUJ7dEFm74AqrENXZA1i
2CcV+hiZ9D2xLqhOBKf8PnD64womniaewhj2LXVaN04KB+lmrf+7R4KM7nY7k8o1
nINGVmjR/i10Smr//gsl22lJDp+38ZM9kjK7pPi1akFZhIUSti84m06UnBYoSCsL
QOnoKdj/Q9WSPypFhmZA5XtYRPKKzwzmH1P2nnJId0OhKPaCUY1vC/Ta/TTjJoLA
Jigiy+KGRILhDtMBq3sqc7xSzVuJQUKAKmMUDUdEGBzjCqxCNc320WDrGxuOAZW6
eDMuJfiUD3iL5hdAwjX1JLbyvPb6apPjqoz3jZGINZGdxHWLjufrGLS5xNvAGpG/
VFR+MAS1wdUS1PvAXTfS7Qqf79W/xD9LHAdZSj75xXevIpU9WMNqYHKNDDA40/Lc
ysPymQSZZNv9IhixyGd14r0B6GPtYhstWcs8aOUKHkjRN+VcgoHiMn/eTYWCQ90d
9JOoruLGZFRwwoNLCXcnEI2zxhAA1ZD9qrIalu/kA56IJ4SLZBhdZSMHviLH6e51
YTJN4sbpygGdmZgdMB1XNWQkqpTckT5VsDwxHQumGwKDMkay8rfwGBsDpR1MQj/b
6px2xdwRy6yEloy/t2Vj4YT8mzngO0+q6yUMUoWAOTw2WJog8+ejf01m/SOFJNsf
HEYWqDjNvG89CBRbfwKR1RyNL3dFgqJ00yRMlo31ZU+e58lhp4ojw5EmrdB8SuMV
F/rwUfNfNBzxTLgUbhoAb3YFwk84UiruJ8aLD9wPItYB7qyaoEK4kpKyAep9cGqA
JvIhuyqLPdWQ3/s1IjFeaWCmAlXgHNSz5kIMjvN9Sc/sy3COm6Q4RtsW9qxrTcjK
vuk15z5VQeToBQyoSkDe3aE1p5cT6ieL8ChYuASiU9qsHcmhAZWJLLdTfBJOR3nO
IpNXE1JnLZnAX+YVtOuDrik4XDSsPgRIxPXRdImI7OHr6/QM7oBgLbkQMmeh4YRf
uZt6Ecm4j7TWtYUaQ/8606Hosh4LtuIKfbk8IWZzqiw7yas5pVepNnHadbUewUu6
ZlB+u7Y2mYcIK4buEW7HS6uuCjCeYrcA0C8qdvKkEMprxD1lJhMRhs8SJLqxQpKf
tAylM1j/YTQqEkh7u0F3eLiMw08mNMBQgvhsnqccKnM47vNW9aBpQVHrJlBemolB
ZEQbsN3mfYyRh0VgFDtgR8oX1zay/+yHhnNrMj5jEa3xsVLIxmQJHKTUD77NPXyI
5knGcbadwfNlsO5CFufWIxOllVcz/R75JS8UlrJB2KANN8Tj/A7W7+nAxkm1ddV/
KHc8P2gkzC0lnYxlxGQ73M6axTaVdx+2/v4clHty63ts+5QWYMThf6UUsMoHTvnP
UyAwtaTINqM4n1XtXQSwQA3lhtQG19WK3L8iVwJ5hTbPAB012tvjfyHkGOQPacfJ
8MqwIxz+mMRcgivf18EtCEbdP8tm9AlDoZnYUHoKErpzDVYQSrGQaC3dpYDiFUAy
yD439LhspK4+rk5rKtEIXMnnvXxAuME/2c4tPlkNG9+S7riHD1MUkgIGGAGaqrXl
6W+BYrwdQZHtchKCydXnQkhzoF0cEcmqw6FtdSDIJaWqnxYXh26BgiXt4e6FVh0i
ytKOeWcQrZDEcc/5fAGQ312JDY440kxnNWezJwUgnZSfZxD7cqj8cE5gQCGROCq0
Hv4o2BN9CAQAAlZ29ERo70oVAufYAUHH8JU8qKubxSx88owr0CLMbX/tint3GNWl
5EhrFsOWHq5kRMpVNSGKbu66Dq9aYeUvHu3cTq5h6r7qCidNIc4Xo+pih4Fp9XIl
HUzLRA8TxhXJluVO7MD68ZGMmnDpUUQlHmS4p8sOMHs51KBf4QshS/wiS8wq7R14
hsa/ZwldagfYaI4uuIqTrXew/Re/8vb+gr2eSgEFj9VHTPN7Y3nSgt2S56HKQ3SY
vcJYtEDJCSQmL+hZaP6jN1qK2ooBu077eEyuYFGxE0XJ3E1TkxQetl0E9C28Cjot
w8ZO0NHzK9DJ8a1xChRaLPW3bJKepF2wC3D1jRzvVgRW0ZIUm0fuRZ5FFqVtMJl3
q5DhgDTuFFr0PTlNtjvfVY1buYGXPi0s4qHeeytRBatO6Iu6bFG3zvLjIBFoHKet
tuTKTjNNldtQs5QicgMJt8IyHI/PUc660VjIG5LpjKCq4GQfIS7bW7BM0JHK3m10
mLfvNTnQWjQ267aLm3p3XU0mxUBPNvngGEu3TzRWTJGsXztHLqVueuX85NbhtWMd
+Ziw9xy4JG8E1fGb2hhaIKIZFo6rjrGBWBPv0OyTM8GKOuVMfm5oBNGlBOcjzHs5
ZD92pZbqkhEkCWaLz04im2hhh4hJDHi6iFW7V3Mzc0xOuYxbMpnZKKGSnIMVekQY
J9Aq9MbVHNoSN3jed5lGeqExPafkeL226nY8BVICsCSB7VyFm7TsHi+7X4W8o5a8
GMVsAPDQW2ApLEKP37qIIczib3NhVZP/mo4KWq0vnOlwQBMWYVQPp+PKjnDvOt8f
mlHqrZqeMqeMMD8s0chSvzqsxjMIXPc9mdiHAaH/7T/7lTLwDEgYtWdBFHNV3vsu
VdsWgaqKGznRksRxNTp3BNzMgVDwEPs+VHUYacAk45987+ExsTMn3Gdpbngk5Myw
ikPnYjd6SVrlfdbQ8U7Wj6Js2dlrvTp9HjeejmGl2bkCvMiUx1420iC3vAWVCUTX
0nwNgaNZVznR9tZxSxrl/SEsKG9ZPP9AR6Ac59QNHO2ZVG2eYhqeDbPN+oPqhOlA
4csUjWQcwOxFA2kk6WlHl+gSdVDl3HJFVPJeuh4i8A/NwZuhmPrA+6mEuCjq8x7U
l4QvWX6EELavcTKFRvqYOJZwmg53vl/aYuEshbGhMdXLTJazpL9ZWvX2rGFRBD1Q
AKwOYCAzPTubkT7kHU2Tjpz9whgYR2gpeq33qK95MlqgCZVMz0yqPuzPRX6acKaO
Q0lhANhnjy4Vt1ZCtUSIkhL1wtoInKr61iZ//yLAOx+1mSWxkp/NPkDoJjbp3oTc
YyKdS7ykAPp0jEP5Y7uabxE1Mat2Q9+dADnMlieAG2mygtidAoiZ5o8RPz5D5Y/P
La6DVIZ/lqtjzBCIH8BJOFdgX0D8L+sXH/+tON78GG5AyN2DMPH2sYIEsv/tofQ6
bXepJhmLssME6Xi3lnduTVJ9z1BL+cUxMvGBoyTakah/kZ+JKklDXc41PUyULifn
lbZW7g0bLXK/O94I+oVuR5gwU0+i1yqy7cJy9+kq0bGuIJbEzWXILs+SBhIgUUPM
oT0EJzm52utdYwq/4rTirdQZl7VeumSVhw5dwrC0Z8/9Debx54oNx3csCXUMkIqa
FhZbFz8abf36JanQEAQWa1KFNggbrlNUzUMQWVrbjoEGUsTyIQgHdIbh2XtdTvhf
j/Lgoj6x96dnDv6uLbWt8b5q9ep6mXBKfMdq09bQtuIFGmjhNwk4O7bcVJRqVGJ1
gV2i8b2XruTRWuXqRQ5h4t1p0BmZAVupJNirtT/OimrI68EuQzufx0Q35eVhYPgy
ILEYaO0G4lknPw2tePDOHp6Zob4KF2CMXpP9ljSFUokkMBw4desGfaLtzvjlqKY4
ravIeXWRlrSFZjYgch5NXgH1OISPSmYveD3j0jNjU2Ztl+ok7LSk3lcT4BbefgpV
IaEUlqu9h7duF8OSlkWA6r9KqQ0c9K+KZNUMWG6sYiJSUXtzGjYHjtewqib+Cwuh
3yILrBhIifo+bRhKEFOUeM9O86Zk1oXDXwVKjVnr4QixJ1hX4xE8l7Ab+aBtTcBr
WyjTxTsILXpZeVzzQ+6DubQeK1af/RYC7w5vHQ/jrxTKfvmqeCFsFua5ZX6YgbUm
KrV7VXlxvWhfOKq3o7h9XzptL4ZG0C9jPZtZWpmwcCcZh+hNQ/i9mNVk5dPj80ww
2WbI/syzB89wsQbtMDmyATuHFg03Io3DKRYfsc33kLKArO71CQlPT6aBq33Du5w/
uhugOpWGMofyt/Qzj51ZPIVv0VZtxU8uiU+FZm5T6MDeK1gmcQjoDxMmIBi3BFiD
Fqr9Pcc/EsRTSTKg2cFgUvLYYMGyNqxXDnp725xSKPrg7N+yJWruPbrl9IhYNgJW
2rVHthfbu9unrf/zhLrDbRfsKj2cNSJgPBCxaluAC10vJAgTz8w5NFmqsJvi8OBP
8eMxp3pBFv14X/l/cbn7FvgNLDou9qODbIYduD3M3OBpZLJg6XIXdl/HaPCtJf17
PC3S5pVBiMP+/cFrgBEhjNa98DvZATn5QaD6T3EAZ3byU9dl1tUD+PlmOscQ2C8D
GudQ1sRiuoxHEVQ0pVyMRQkYawAQ2b0NllrCHEd5L/HFvacGs4eQ0y3QbEKPUQkU
1L4aX99sjYEenRiPskAmoOVWnMpnEXClmLURYFFgw3JEH1g6XaoP5jnhy1MoNeAs
lNUpiHJmZpdP9mnup9IxpEvHb1/AIgYLVKsMsr/CBJ9KqyQ12PORNMwnNkFrVT36
vH69EdYDjTF0LHStMi+I5sBTcdInqPLhSMBU928l1ce2tH3a/PLidOKUTKJgC+N5
gjIm8gQBlPO0CECAWnRn1M7SnVD6RA73XuTeAKTAhSXRq+sEA0ap45moe6yToG/Q
A5xKFueZS7NIDNZ+fhQ8mqe5f1jXcXDdJ9AJnWvGtwesDI+/4TDbqqJbS7Obw+cP
Vm1+OYWyVgt4Y1sf6xl8aFaGAGT9V733X4S/9bns5jn8AbN++Z9H8lc9EnVoKOTy
Ml0CpWSAVrCtrLaAuGa5tIgEf7pp9boAJZUdiksV6dIVybkY7j+WG586iAbhUTRF
W7S0fpmCSTAkehy4PzMpkSjp8VALc395fm78tRfSW8OlSYNCEul++XGvd5WwYrvH
o5L7tXOvSCIuPerxfQ80IdwZQD9bfaJBLhc1HYdX3eF8Vmrwx9QjAaxM7/9zY9Fo
h/U4oJMm8lm1K3fRYTWWOH1BAZ3HHJYqFuGBOZOIRUe04qVQ160OLPjqprEHRkCA
R288UJsLLN6bpl9bHKkllw9sz3RG5ifi7A/P7jsMwRouryZbarMuMovcmI9J2riF
a50nHe/GjrrBXcWkWyLrokA1ZAXiD7c9g1NaV9sZbzZeoYSNHoNRy4JfEmR/pCa8
t227t13wajwxOiIrsg3jRKXgVjQbwQwKh6X87NLG+YQE/Iiu/Mch1L9okPJxdolr
jwmFFY67dxtWXmDyEMDHGrQICJvWR02a3vU08MZIOsAa93ZiE8q9vq/ZWXU2V+CP
Max54mqoJ/iAksjIyNlHGjBha3qONRAvyBGryHgENlUJcLsvuo4AGtELsnJa8A1X
HJeod+/fg4/W6CWMCUwYHmDm0LiCXYAkp+kCYQh+zMPK+K2s6QjlZFoxdFalmwkt
ep7pt9zk+OToS5vWSh06iXQH114FCzCKjUZrtDRy+Y2dGudGtJ03HsnKmb/KSTqo
aPF8aWcYxoxNQg8Y1FmKY1r5Iuy144qcrrCddKWnMkSJPvXz9ZUFe2GKoLNlo/US
J8V3ekv5S9A6uLTvjeB/qJrdDGcRP3jdgaPz21LnpgRzMXlQfGR7qdDiurnDLO0C
uH3g53upY0VyFtyfVN8B38HPhfSIbVo2fCuJigChq/VA04tZ6ksOLzTo3pObxlQq
qmey8GsEZkk5q88pOsq6Rn2fRC0FJnqTLOgvYiHjhWbezdvsB0M1KXMjhXmss3gR
dDI7RQY26Oizr+mNm79F0J4ejVIEJJ2wJ0oDujDfEriU9ElULOl7YhOhZeZW/Gtl
i8HE+/68Klpczuge2Bt1zjrYDPJKliwV7AADLQy8jmcvAy0pV8wqt7smNWRQCj7x
aDuE4TmoG9bzO2Kq1NLgMqIEJ59OYslGmhTAUsy2Zd9Fn/WK5Mygmq2IyBURH+qs
YRtIK8UYHJC8u3WCOZSZDbA7S3LueO6elfz1ksOv3YgBBhKusHjY3X+i/cUdOoGB
EiGdJOUB+P88HkXpxZUrrEzPDukU/jR9Vrg7BjhuP9ZQr2IrM5AMAe1PTwQ/qWxy
AOkgElwNG90RxwtgLfhvYmef5yq+9YHlGseAwlIefJ0sBMb2IbCLAS4Hwoi+HC7H
KOnjt/+7u/2zmYufPEsBvAVr7tStOmPiMtn2/S1ijolDAGVzki+IIfZpHpv/8BqL
KjK9frabQS7w6U++6DolXss1iu6nDCYt1/LA9IY6uIQMqHPQYNB8Ju683b5n1GwC
C46WbVJSeA1go4leh+RV/85Hp7ouMfgmGizW9YCGlGk9mo6tGLcubMzPuihVvMgR
t6Oswh/EsJn9RKOmnXnu6EldkVB/OCVKa4hEXKkhPQmjPbg3xDNHt95f/tCPx+Bb
l5j0ezqDqqKQWAgudwF9pPE5tpX0zFFVLQqzljEHxiw7lnJQ8XQAsXSKBIwbjjQr
J6CKGmiZg5qSJm3BoLNP7ULiYeWeSW49uaqPav4iYF7OEqTQLFs2EbbVwXe8RO4o
QS3v3/JqXw3yeg+mo8oK+PJGuKVHxCea24AcRb1Y9vSK2QWbiRT4TsCyJDDS3LRA
YGp8cwZQxKdNTBUxScvDyOKxkihYJzFrz4nMRT42tYowXs1Eufhbpy6CfRgjqjop
7YlgilSF2iqC0D+JPQuPfB2tRJV7+U+GeJawJNh1UoFG53128LKDtOlgJ7pn+rIX
HPowWvyPKRoNxBtUzMIrNY8eJRl1OancF9FyeHGphwOVqQ8zAgSEI5MTKhOGap++
cyNYrHzrgfEUHrOuvPAUi5yrRnYxrgzQY1GcsGrueXjEIq0hYrNYku6peVTtPH0n
OKTbCgoNQOXM+6vGTes6QuPBZFFHS/pZ4eesHX+66vSLBgGBpdO5an/WH+2/R6+i
Xv4PfYNj6wn3DvQlGD4B9eYq88IHF/AG1IdKnchBIoTjwjSsLdpAzU/idl47I238
f+UZlHX6Z7fyq6zBuIAGKk984TpesqxW4JY5oStkrns6SCH/JQ9MT9BZYOlM57ox
/0UEu0rZy0LB15iRwD4i7buW6THVOogOeGZUc5ETRx5Kj9PbNG/QYViS0l2WvwH+
CLVbkl+fumbOdFqHPPMmQUFOx5ohjwCLPAlAZe9H9gxS9OiSm2QUBjqXkZoE/4LN
PBROKQDA8+Rgpiw+o0/1n6qaFlTGsRp9JSgt0tyG9B5RynopzTp8r3ulIg3jcAPF
jJYI/NKqTMYD7Db2LRfLwXuP3aftU4c/zy0lEqJBMyYUWlKTjmHQmhjL9qsjdXa6
dk1/vwe7bytt0c7+uv1WQ81picm0tB8xV9D1ysZH4GalQRchxD96ohFGQttEjNom
JGFetFjbz56eDnBc0hau4efQ25eIPkrK6h2WUE1th0SomMwgAYGDDVN3hJtxv9Tr
UJ3iwFRhdynhRWPB29z9AVJHF7tQbowmcnWpXwdmgbVWv0VXNYq4MU3BQCPyBfy3
dwoS4erB6zhCoavYG6BS/zvDgSRFdblgb0YCXXGL9T+e9wrkFBJUfE4hd4lFvy0L
Cb8HhkyTRntU1R3mI/ikp+gBhHWKQKp9fjXl+N6SnI/7ogsW9qJHQpcFXs/u0AAV
f2kx2ydB1xU8TWoGIUDaM+gRhMonMeM/kWpmuBExs2Vx7E+q6ole0mY1VSfUDkj2
uoP1TJU8HkJprioP0W3b1DsAJm2gwAmtTkMJZrvhRl/6+EgLwGwfa9bamfA3fSp4
YwYuw5QblLKe/13oMk/LnYx/dql+4wR/YbiGH0o3zv6t6ltY9YkOZHbwMAU5rejK
cvUj5zYM/vKSfvPISWaNt+e1Oo9CU9CMCxRpqdOML2yg31I2MdfRhncCc/8GWjlh
5xRIOvqmqnYm59xjqaNGRz95pORAKSfVZftU9HMk0VG3vxmfCy/FjsL0hD/XTc9C
SDgMD6FosJ9JNZIUTL5xCUkPVRkPIEf/5hNRVpykhaQyiz/OCmI2kvufsYj82uW/
w2wnjVP5NW6/JY5ghnajHhhBe+uoF4gWm39IkFPFuRaF1CaHn+CfXBrBgaMC5s/S
Tn4zVo9UKgSqosGhR2GM9Svo1Rr3tM1h0t1xUZZYf+RHzOqt/kKh72M/P7mkdNJa
lE8qEOpMTs3v/5MT6V5h5aB3HT4BGuNWypoeNn2bSXgdrtXgipkQnuGh4Gs/ZN0Z
QSf2ffFYNcSD8b0UexwKvPCkLzVwAoX8dWE/xYNww5mO+1PXem2w/UA7PLyNwldr
8u4Jv0I0ln42mLhFu/thur200fWxjKLqnfdqi007GhZWb2YEZTC5ec2Bb3ROJH7z
O9WNLzELNgzkStfy66m/9QFhf24othAOyonzeHFq8GoxJTcG0badh58ifQEfi1RD
sO08b5XS8f8aZtwkpPyOmRO7kwhlO5LBY2ODTCMUb1wbO0i9ekF/3WaVTJ+B8Edj
MFjkd8jLECejG/xdxrtL9hBBGfF/pp9AcUFEH5Bu8z4ec67nkRko1Qiv+e2ET/Ws
D0rJWkZIJw4EkUzFgPU86il4qwP38KIx+TrWJzGb5qmAeJANV9F9fLaarLq0V84Q
VPWwMI4IeZdNMPK2E1HhdbBPBWAQVuLP6VLUbs+7Qxus8GedZbZX84bGoqbPUc7I
rGixRL4Wvg6qErz3q8DwCDIpwAaYQErRfw2QBuWWQ62T+WZEAl9sA53CPcgSiJSz
uKhnhnpq1a14VOQCo7Z5OPdZi08Hqscf5T6vTRYsa6D3EdKDaxOAL/hRohnMunJo
P74YK5cnDU/JmFAsa+Q2H+9GKyKh/yKdm4acgJK186/67k/E/PefFmV6QdZm/7R3
b26fbOaTx08ROjZg9guOpLIrOXhjqKf4rNwPFhaJXCRih6W7ZL9YdSV2pAnTJ1NQ
8LiMsuYmXxVoYykOM1mFnDirZkcoWn0TZebUmhyWehzFrUGHJHIIfuy3Yh1cy2wn
AbNxzgTXeIoaSROXa8YBIRkUeurNzieCIZjbM8bFVAZg6TUEgZDIJ99JVSW0tAcG
4LNeJHhEKA+UePfEEVML+hOVi3GWCOIgtZC3alS+4PxORzGOTK+8JKlTAXQmiutu
cjKq8lSqdouESpBWfJZIN+86bpT7LVi1FD56vmt26orfUgLrJwGp54nC69Yd+2Fm
7wBylRnOowp5p5KEGKhkLlD4v7TSuVqvV7pPaTWuvMOSytwTxYNiCjl/5+R6rlDj
CaWZvamVWCV/dkZxJEo8QuGc9xKz7Jq11YuVt4iTmj0kC+3nxNzrvfpWvK/lF5UW
bjUmpRvJ9RMsGD9EYJU5E+sP9Aai7WP1IDOY0qaxa9RdUTY2lowcle4XUmd8dZkW
4CfYpfz8IJQ8PefAQXdkj+c+ufFLprR8JzBicXy1laDFWUwc1VHtdNlrNPFLttwA
MKAwOWHrAkPFVKz8ENsyCiAd/mGn0SMMiLDtCYi/xy6hSNPHEfBTfnFYjHhT7/RC
1/qOHwOmEB/9N7J+5CMdyES74RJKy5/7vPU7PevxkByOKm5VKA7iQEMXR0A6TkbL
OXof0iEXkGCAB03ZKyKl13djbp5IQqu+UmcsvrWKQifDLV/gWKK5+6P/SOUUZLrW
u9+X55WZlRMT4uQ9CLSPG1sUPVeXseJcC58radf9pvSA51hXI/XbucRKQbP+UBOn
QRzD4dF83Xt14JX9CEonXgW5UXDJbGc0WTd8S93IcamE4APjs6iiUguFGmUW2s0t
ggr3abyE5ES+QDN3RWm9YJsUOVEaWgXVA428iMrlbCtr6Z3frRvdFmTEG5jagJnU
QDSx2pkJ7lzHK1MlcEpEqVkGGArPpXLl8pKHb7d4+pk0gW8KldJANPUeaCQDO57o
oGWwoxqwAD0UKqd9NAHHcwHu38DwsPXQnY2kWb53WG19neXhwbPnrJIip2lxldb4
+WrRxSYRD2vmAHB22Bzj1c3AbfNiuDaR450PtsuOLATtwsNaemDSq9Yd9OJ1Cs1t
oo/9OA5/1StAHseHaAOf0FWvc5SQf9rTD7+UE4QpPWXQ6JQVEUsF2ugMZzCkf1J2
T2cOrA5ZjDtr7w7uZV7rCj4Uvq0bSBR4hEeA/WhJxpPSBIv71iEVT6CWVEhOkvhE
OWDWOItAqkS/hOS9WCWp8/RNLJ578yKkmQYmOtXMFw0kg7fBZu/3SdCZsi8Slw6v
McH7ZhY1py9R5xBim2SYe4fY9eOyP8kxgIkNzBlumpt8kHd0UBYxTk6h0sOqNPsy
PAh9jJk65fA7asC62YQpO59CPXzrOCb/ZjKaNbeNHJmZtVreUTg1KLx1HUHs8PE1
iwwniA8CgH84wHlTfpTX5UPa0N2xtLk7sjGBkmbAANwhRThr4oRoUu4o+CoMO8F9
HULreQoBtvX41Q5UiFV1+603UV5Xw3rW4vJJnv9lBHZEcBuhAJkJrnqJ1cBy6sUp
I+JtWJbDtEil8p/KdQ8SNtAPfHfkiSw9iCsOV+4QEk4LOQdi6SWUQAPDXfeKrykW
PWjLUjN+z/ZQc5f4KjxBTCB2s4HpachkXiZQsnE93aWA0Xls1Xdxd2L3X0GKX1Oh
uiKzoPHSxlVFUdI4+Mk6U6NvjD16dE8mVaJOjymvILqc5i933owgjS6IFngyc96/
yjWOP46SkgszTL5TuqN5qZLOW0vIAWjr+x4DBRs06zSj67ylmzGAd0YxSZWLIO1D
VTU6f5Vt+kDgigXSJxVt2Iw6HOhGSBSRLHwcvNWQu5vd+Y/BOLNtdLASjAFF4EZt
0BOO2osfljrI9gTI+3HkxLepddUkn28l2R+Rf0d/LXQPtA7kP9R+6rPISt6v3Kw5
ILh84yYvyUgSj5Fox+/pZjy3inBKHnqMtyLw/dt9cobuJyLloEfskBhPoqKhNTh+
SDry6gBwRfhUPYLR16F3zinmsp41sdmiLxIOwV1x1byMdctOslumwHgH2rStu5we
aQS7coMjl7yfQY41qVcxXSCd1SntgEoUZpGYgSvx3qkn3QLAn5XWoqQUktrmf+R/
PCtawiuRL+bFLvshnq8JfF+dAMIE2az9pWYkbYj0BcM=
`protect END_PROTECTED
