`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9EBVvKMlUmLdwbYoOIP5982o6OuW4wSn4x/ZQet3JkZV7IDJMKTJcjMzdzpZoQ5s
8yENaSgu4MQerkETTDwrfobQLZ3VIQxmXEWDECupWkmxALFVu7mAEyLxKlyDo8fj
C6GE9r3eG5KPHhq/PJ7iWZ2UG3aitipM3RduJrqktR4NbX+6bo0TitQ2UBqUwAvu
ky63CP7iyxOtdIEBTFGumSgZFbZM7al1PdnxBXl65DBjEbvbrJ8/9XehzULtakeZ
QWlozmMyCdd6HqiMmPY4eqkSfwu3u2iBQkSjD+D1P8SIE8L5IcSyfzsOXZQBkn3W
eBIQr4LMomu1BUERLdYjFi9FgKtFRvefjNgOKymsUFp0gOKnUMjtMEnh/WDG91H2
gRqpbIqrbnpVStfrvNUMSK2l4Rxn/93hbKrNG1+jkYRRFVPq2L+UGpKznDHrHBCl
4abqO4uM5zeU3vDMJD4A/4BFaDT6bQ6PSUpbq3GcV9VF/Y2Af28mZoT6/uP8tMrt
fh921RvK8NY6pHvRm7tZF4A1mN/aLOcXVDPH8iitNYbUzcPYTWzrTWSizgWe3Bpo
HfRqBWxeFEZJ9vpA0g8SRaBQtc3qmj5kgUOuGRPGiLlgCf169KEkurVTi7Twxz47
myq3NCsxyN2N+ipfAh609GDRWJg0/YD17cBXQ1kXh1GCcv8XR4fKFQe1nr9cL4UH
236Rcp/eRypEtCFffFYHYXkFnpYNfsXAhUiCmN/JnrG0kIWSqQEFM9PB3CWNbod6
PB9JMyjpqBR/69ulOWy5o5Z08QHCYiHp2BjAVXMwC842MG7P1/hSIItKG2asSV4N
tMWINWqSvurxeeVWWfwSyY3Ui0+wPFiS7KATvXCqEGGCVqV57EBK7d9gYQBCReo8
Ci3X4of+ceeVO/vybJd1RgmQC2fSBHnL8Al1PVWNF3fRLAtk7c9Pbz0qmtNXn4yl
GPZFcZtD8FdMcTPiAhgU2pOD0DmTLT6yKrDb/DIKqUTbiJSK/a9z001T1WW2r05F
umL6Lh5YqCZXXYp3nI9TDw/mCbd2d8cSnzkBETJaCtV5atS/LkYJ5gmKnsubkUGE
tk5iaKXI2Uhdbpl8dPKN49YbFvFAjw4qZ1N9rSvJjJd6pma4xLPNV1O/zTsomfKN
PIJAVhUdv6VZMRmQcUiFAJvl4VK3yLUNE5VH0byI2h3KYp/ALLLt8ujktZkg1mPM
IsmqRbibSON0DuRWRErEN2m9dAr9u5UTax9gMouHf9eWYCHgweRakcVeJl+PjQWj
5+ePsw4QJwiwbFERaG5px93v8wUIo/YEkuSTO7L6/PwTjsdossPsMiT3FGDG7mAc
nS5K9qGfEqInV6v2Uyf8XEiC9Vea8a1iq7018SDvKP10iOPZldKN8Nx8wTybsH/I
aK3/RGlNrGwqnEa4fmA1mssKY6ulQXXMAyLBkcF79IedlzaVQ3GbbkMazM6lNls3
uQErZGlOSI45VRr9ynFmysHyLQCZqTlGWOtNmRzuz96RlKpQ1H64peeFkTBwkNhu
k+tyhMnjEom12H26wuK4OgdNU47el/3/nA6HpebuoevxZLl68jbSmMAAN8jYfGp2
hDcvtB0keLfx7DVxanEPuHjwdpO0eMNIuW04KMaVJTfnxqvFO7V97dyLXADwxfec
gzNsxd2OkaP4GOwrzVPZX1cLx7Ii7WA9ZSWWr/zOMNYP76bl74kRocj23rkGCeR6
rvZ+H+Sy6dLRvMAe2jzucj/60vWVVrHv4xzrPb+NqRZ4wWvMvF7MA3NeoqvdoBRL
+25RW8k9/CfcApDmml2uzuDWB8aSxmyjdYtDyp64QjRMBntGmDGn+E/XZrm3RWId
VrL23CM2zabk9rCwKjrIzqnR2KW6EYrLmOVjC+ulpFbzukhHXL0BcBYwfe2K69NV
rJN0btoWgEJ9B9XZelnUGRq/FJj9o1ha7bDjub1sjvJcbUNXAQzII6P9JqwT/5ot
U27M6h6dvYYsHTsqk796aawe2R4pT1RSrj77vPFsf5x+uH39hGV/qV4g0hDQMiMx
5hT+o6C3x/foMovlHq+wrMswhumbyhnhDpRHbl1sCZGwZJ48OzRvXuXaQsP8t+sr
Pn0aVA9kqDuHNe6//4eXq49OV1fdWrLQohPtrmJLu5EbCuw1Evo6OQ4zuaxYmSg4
z8WLLJkUCWW7Rblzx6ZIlBCO4qs7hbTmLIQNwIpYyVRkXEd4gSHIo5n0PoIKUJRw
iO78z9a77nIhWgA3o+7e3Vg6b48ZS76Lr+JqOzl4rDm3ad5pStC+Pei+Loed4YH7
LuShmYD0lTyElzGO6F01E/p5v8jrc3ogfBh99kLGlE4LMCKgmpT+MR6iXRf7cDlx
f6jJfm0nzsms48EofnJkS3+X1U+dwXR+AEGYo31s4Ijlh8das6a7X2EiGUVg7bkE
quwwVRYm83f7Pj2styAKHdMsYllwoNvMvXTAMJEbIUiiVBnDuOMudQoXZhDfq+Zt
U0N98kpp1YwR8R9DGqve0umoMJGLoh00sgOMTx4OAYMv61unEeyrA9/9D1jaqPa8
LrCC8+pke+A5CaHWSa5AZJVAzD3fiN8XQlEFkGBHsP8ExvIkZivdP1E162KBESjw
bYMDK/4AmS3MOZ01vL1sb6bHBqNpAd612VrGKc9krVnVevaWT+PcbaApeFDEQ8kd
j1lqOvyoYGu/P4Gi+GIzkuurWlUr0tfXcOoPQ9jjHj7AzAA5x4yn1zAacfuP39MH
wKdjxfz80nGRDMph1/kwEA7ksAb9SXmiUW+n9Q0oDG0kySBibXRWMeCMLLj9nSP/
vN/7ZZqqczJQ18d/NM5Ts8cOLtsvQwk/ow8nif1DuTNKbtUUaRFmr0SSyf504Dh4
rO2Btt5psYb/V9wVrdTUBEiak9ZCb8jD4tCaxZmn42koYrAQVgtW6nR4bXxUfsnf
0CuZUMakjMrqHt0xrfxFFFUaE0W80l+6ve0i09Jf+CtJIPEsznX2TLnGVKZYyWBG
VV0aLCRpbXawRaH4HhfMtMzZi7bGEyGgYCchEOiIiYwBSCu4hz5lSjrygscggPIf
sm8JCydQuHkQ+XBmf5X+QCjgaz9f5Oz4BHdLlF7L90aZjcS8AxGw+Q0+0DZby56T
NzOIyWuP20wrFMaeh1uUB4hxJtbXaAtlJvocmH4Xnrr509LFt9ma5j60ikaCbfrq
bJoNnYO0H89ivy2vj0ksJsKEXLMJ2L6GyfOQ5vdBKIqA2PGGoyAk1hBmR6wzFHRP
fMIMExnUI2ugb7vHZlhzR8RCqZ3iUhXk0/J6819SjpPySf38Dx7Cf/1Y8hWcHmX5
mifVBPIL5JW3SSLMqhvf56lgylkti/hjrF/iu0gfz7Z7AEpuXHttmvVlwHLv2qIn
BFWtPyE2bpebyb8NBxtkZW136FC2iLYAcn+opfrxXA1eyzO/3yRum1Bsn73tH7Si
vflcnQdbii0a69XaHmyDC5J73xghz+K6M0HXeIZY4URFhdpnJqWxo/hVC3IpbifK
ALyjlvtDWCeFoA2oLTB39IVNFE+JDavAa08LkSgtTUqgrzW9DFkA4wBJrOYytk0M
wsOT0kqHehpqQM8ZDO+zJOXbhAmZ/o6MCiq//A3UoZhX2+6ZLGFJ9S5N78WwsKmK
3YGhfLo18bx7eplgOFdsOSQrMQdtudxwfIqH8wg4AstNGmMuLlZLlvuH+vDJ+g5n
Z5d1+p80/WGdOIbpYcWuf1T7rS+rXXORE2eOrk3d3hfDcUKbyRqtU7YHeCT1fkCt
BZAG012Dp/nbORzvghq2pSN540oSmQd+fq0qVaBFaSE3fnZgnFbvEF2y4rY0SyWj
OcNkI965bWLuVq6Lzxj+BGLwkTHzx4s129W12oRr4VcknK//gZMkEADcILYQzZi9
8eX9k1zLUEi5ez18LAsjhytP+cDfP8Fxs/CqD3BEk4XSqBAh9/k/Nm3jrV8WTWYU
3s2iec7LdDWEhRcNxQdisbijFuo0/Y/e6btc+MIKl8M+sNUOzdziorimISlXATyT
FnOS23lkHY4guA0/eeMNVq0tKKdwopLN3F/iN+uylzsIH/i7dWlAmq8SrU0wgLhk
5F8R11sP6iY+mzjVzmV/Ub1CLGrtBWEX1/VW8MAqNlaoG3FiE96W9rqXT960ozBv
RYR6lt6wtdGWul9VSMvQJ3SaWuGBC2krOUGJjsK6kEGT5+t5+FqDKzDgh6ab3Rqg
Qgs5tXTcL192gtIkPOprA20qX1Eh0TyqQOpywt/0Zhga6Vu3qL/pyT/psLprlhva
LJLVW+MgS4pGtJYDSmMpUSo/y1COJKxWj8Oz2ezoKVkTBQpTbuvz2356ZZHb+Lpq
I2qqoK5KTGCzEV1v566NnbC/GR2rElWzQDo2VQyBMV+SQoy7dx8bTDFEZyAVEZIa
73WmtnM8ycqY0xf3F0mPUh2QeGYEXnwLw6D37dZ6ctsBblZxCR5Uj9CfmR7HWIPY
UE+6XZUTQ+VWDvnPCi+Xphg92UvpZCedEBL7saDvznUwZNWyuodQ2W2VekQG0RQU
p2yZSbofF5PNvTHrb3ICT99hhNpqCTBVc73Yp2h09NZT6O61kTxidaheL1lOw6c3
kuPDe3zT20zv7SyFXX0ShW01OkoKsrwTGFHvCuCtbm/RSNT4c0KpGmum06NlWNk+
fWyUQDeVRRCrHj2VQB3/jPft6Tdo+a0AAJkEQfEDfjF+NSZM2+PM7/lltLo+91rB
PxTLtBeQOXlJDrEPuIliuc2XQNmM7ROeIwaf3gUUj+NiXdUi7typxN6DJle0Cf7u
Yfxhf5Trgt5ICPlHSov8f2x/+sAwyyP52muLCm/8laeA4D9XJSPY+Tcg8EAbeDIP
3W8J6BF01jTj0PHa93TP/sOEE5+sFuQ9HhuvjD6u+o8QfNtN+XyobyoNhcletrjX
Uw5QS5cmO/0gQpS4C/VAUjK3Nu6QtubUA4Ryj4QE4otCy8QozGkDak72kc0M70pC
Afe1MxQUR4NTXy2og68DGjaa43IpgN1s3hYIpVmN7bXql9qvMqS2daLGKev9RWx6
I9GM6qCORnpVmTjz0VVHnDfARXIx3tBl6c2pFgKJOhJAXV5l1lLEz5jLEEm5mF4s
O4zMEFd9BbFLouayRa78M4cPKPqUmohXEegVHeQXNB7/U8jMdUYT3y0CdKg5yqIO
yKvOT1fQ9/LZWYwDNx7yhVa2+hdEyZjILKOPqYly/gW8n2tUO4P4DxS/W3d6+RfL
1waHlVVhaMVbN5RSLBaVTZlZVtaX+El28kKSPCvsa2X5H9NieNIeQBgsOi7hv7Ri
uk6h5G5WUuQ75qhRRrSS2ZBjpprL6UVmAAiT2JMX+nlaRaPsbUnRoBj+Nmyn9JKJ
ApRPIvaLMcfU4R2dYuM3IV+45EvIfEVZkPVRzfMzvm6t8IOpk9bhOQ1D5tFtMdxX
vDV0+EdLzlqpmMG+nxNvUhnHauIlh5u+J6xgq8zn55C/qFvJDF8IEOPMfnEdIQn5
EG7s6RY0ydIRjqosmu7jWT9t9SjYYQftZbgajeicMB6lF/UIx/qNlBdEIbMEdei5
puSYezEaBaBh+xqTTzxixvwG6/IgpmFqk1bF6s3uFM0J/dDfB1fGoiZN4ar9WPPK
1vjgzSFQ566xtSerQuHsfE5CHvi3qXYaVSO485rtnl6GF7SRr00/8HgRm1H7YRwc
4choVN9jbcidQZJMuMaMhMeAMiulGoHLhMX7AegQpco/dUkRzHIB6OCtHlFS4Agz
0HM+JE6kNBk0D++Drm8Xkerd3OZnjWi8O1xlwnwJ0wdh7Hlf2HTnGyDHYm15AxhD
vRTZdUxZ6oI40QGvTNJaanBnLe79PllBdTGwt3O16FMjgDEbV3Kb3j4Ir2aaTzT4
Buy/jj40SfrmxRw6d3usXx63MN6KVCb3IlO0E1rfVA2mvEjj5BqrveRa+v4WEIa4
oPCRsPPw7KGolGIEpj99Xq3MApRq81rt7HwrZJ9XUJdDRDtLkEfY2vHsldaizZMC
mmdOsqRtPbGfHVNmHj+fq20WN3HL5fjCL1Qvumhy9q4=
`protect END_PROTECTED
