`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8thP34VYO3nWPjXLNe2WrGiOzbAkCyWbcm85E7ProW98eAB2rlb9bW7ljJmLpcT5
fPFSo/xzuqgSFzOk8A64NHzQS9wNsQ9+XhnxlqRfKfCkgnPxQlOIjpH4li+q1jw+
JxD+WRLEsoUq8lIOtmJ5fLXCQvvYZDM2kiZwyB5W6Bs6G5PnWY4tZyWKmqflOXRz
q5FEQQe8giGH3YOyq6RfV42FN3ToWD3uZznZTFlIz8OZ280uET3U1kFiw+UDbPbP
uCnIWpHBWo+AOdHBv6TyTnLDv5HPVH4ilXtFdcRwYDca4Qyplxs6YDw2htWcgcH/
dVgxwx8bE7bFOC83sBkAB/v6QdNFuUDmlT80s0T+yQDLl/E/0zeezmIzsP5J/X7/
qwgC1OykiEsmGTvy8qsdZSUUiJzMxYyEfduP1W4KT1QMd920XAs/hjMkBok2ACtd
AFmXCB/8syFnogczdzJZLzt09u53h8QvyMX/GsZaCwOtsB06UdfBlm1K8wgtItxY
o4K8Ei/LrGrurdDez/lppiioq+OquzRZ6pF0jCyMk5M1Fq6Zjv0K37ysfyewbIAD
mPSQkaslCuEa2HKffasJ7fxpQs0qicXqXL7ALVbqoqb7Wa7O11R4AhaFsC9POYNH
JOHxuxEb9vsjxdSt7KFd2BBW82bKgP+9ALR4G+9ROapdvG3jG4yezB/eviUWp0wg
eR5n01G6UmKbtNJyz7eFwjXEvzERf6kOMCnMwOnIyNbd9LoCrzP80YvU8+/eu61f
R5WT/kClvTXjyNCbuqH2GSriYJqxsy2nTj/ptDa9QN9r1kSgR9qijW1trLnxKkfe
TAO/eLlaLdv+alFdQjjqSwdkaNTprOTXCqVpypj8utVHbGeKucuBHX6nkLMHfm11
8InUu7Q6VrnbOBqBIcX0mJIv01oAqj5ooQu0h3oQ7Bxs8s8WHolOefAfABtlSV3R
kFxuLIOL1qwVDTjChQ5V2HQx8LcENkl+z+smG4TBZRxrgXKu9XpavC6XlKOS21Vs
R/kxt2wFDt3mOD/QgKkXH7j5+MKfyi47rTvdI4fupC1ZWZ3FENEPdybYcIS2QAvP
1PHLcuhpTIyhil+AjXNGKB5GMLFzpkAG2MENYWHxv/Fz0cG9tPYFtDByCle4kqa3
Yx4AE74gH25VrkZNyMYLND4PEJ1TOg0zsD9llYJIszYkd35EnJPZruJpt6jgVRaE
K4POF7qODOVWQJhu4UFLwFxtCbALrfWrb6e0pdE/z754bscR671mBYrkxSaXW86V
AhjFIfldXwGS8lZFG/ijZ0afWuVWSs0dKOjfe3FkCORV355FCyhSWm0TbugNXNWQ
skbLRAidirrpd3pUnf4PNV1HIo+KoyQKDNZ4Dg+XtK9xYe44cQRI4yJ3rwTuA3/C
/ivuCUL9BZTCh3spd1aQ4gwIf+FUNgl1DfaqXS+muSZO+9gi8iqWfBzpBb+6gNBp
gaB+HQ7VQHdhun9n8i0StNJ8ahDf/vK7UDJNQkxZV2Xl7iBah4qvNdWj6nKiF9r2
qda+4Hu1YdSpVjRxJgWg6yZ12XF9LBxchi9UN/9PdTMhLO0TsbHR+niFeegJsy6e
5XpcPPbmpyAVQV/Q4GYXuP+FKqnolJ42zvdVL54XjN4HUHbLkRdKNoTLF0GabOc1
zozDj67+lMuVhTNS0sdQokkNNMVY8SJVzF+T13XVxo993vU2GtMgOlrKSmrd1oci
gsip6TcFN0fQuPcHEfMPuRTPNxXcLh3CQ51WP1KYaVxfzht4q8zj/KDDSPT6jK4t
HJZ4M/6wu8xeOpLiQ+WHzIPUvvDvwk14oIXeHUMA7Lsj1GtkTmdAFuzKFK39BMG3
oIQZxLKRVvw0VXkS+NdM9A7YlxCaVkfgNdgLbTzAs3T/axMeacwo7rQluxEbvbKo
HorfbiSmIfRikcLqnWJf/1FI5iC+bSwft5M0DCHk/GiNYYQDOG8IILeUZSv4nyPG
Ut9jVR8pPmEaDeR6IPp+80yuGXG/xXPbHzvKy64+nodmzceL2GA7n8p2hQFHbkRG
xmZNps4eW5oWjAdUG3hLVzGe31mU7EgC3QRYJCdKDk23btT3oqIE3pYwz7iVt7yG
s0tSMQssHkw2sGKH1GcXb1rDQrVBJDiY6iM6ja5nk4naD02Wmb6Ef31E96a+NMpm
C4bApmBeKl80LH1rUtenfnCNIaYxPWc4uK/5/3LKdWLCL527SkfUPYf1hwXdB7I4
QZ8srg0t+Vjib81px+EkTu7ZBc39/2UtQBllxZ7X81PC1gF2OmS9C+97VAFjDxul
J8tb56u586ZSYwDNq6WrTrPnNreAG3BEvu0qdDV3SEH2kiNgzbNZoDEEGUvvOgIj
xAVzB0eF3HPs562tMUSv4l4BLmaIB/ld6ntc7+QB+U7DFI+ILPE3SRxsVmIQr+Ue
ciU5hLYcJUJyox2QWTDLsmkzRtKsyYLlJL9rpbPO72xAcDRvCPi6TFYmwfCq4aUs
3vUHTPxfeMRHXy6+3v/+6VsCtBCEyJJ3dSOz6KHiM4D0I07jP8Y3Yw/gSO/g/IYC
loMytvMuxy87Qs8Y6Lcd1DClw0Tq/jvJCQwfbGF4QUo4UIiG2pDabghQgkaixOQ6
hqQeHzoCqX4IwzqBY3gD+3MkwBBA+PYAHmSMZ3yshON3igi9JNwWq74PbO+t95So
zSTsN0WtTo/75s+NWFyfV1nRymkZn5Mi3Tj8o4Ef/CZpZcIoDZyHuSLKMIYn0dR7
gSbNJmHRiuBAv0bxfvszbp8B9RZPxG/rb/WcTVYt2K2JQfu859W2BOJC2V+RefbB
C5wpU8eW28x3Q15Y3JivTLHPw+05TPxoLkZd3ds3IGm1LJpOI9Mj0UYTH8tgX86D
Fd5XIqmuHC2V2oHHW/MT0FBpP9MGDAWQVdn3CFV+84NJ5P0ncxEanHg1tf67mvTm
owwZPIe8X7PNxqOIfGob7NV1YhVck8WLEi2VdMykUfm4MCRmLlD1AHTlVPUGOfzi
qBpOVsBL82G2Qu9fTjHgas8l6ejYxK8Eus8PuwXkFLP0QW+NkMn5JmsV/BWIfvp4
0aRLxsLNh0lZR1xIRQPmYbAhAym4C4ejzeaS79/h1KV2N6L31lN0TCXw5jp2AOpQ
qa4aUul9FY3XJwGDaDZRbDZsfJsJseiE67h58CtwsqnEJgpg+XUx9e6Tf0TUi9AI
qsh+6DvjZQsvY0FY7rCeYcVg45HrntYA0PkE+dAFJurx1kpqJkt8CoTvFdld5myr
a1jsyfIMbm9xJhd3QSW3iDkbyZ86/g89tiadnM1ZWZkWeN86IPF1HvE/Gl3eBW5Z
QvsiCcLss7j9TKZ4PrH/w9hEXIg5hv9aDn4zkhdn4Y2uOVY95KTALymZG2LS8wO7
cJt9N0aT21UcD/Rr7E/rCntSYvP6+y5/35+t5j5/DS2StHEgFj15YRs+iYA0oGtx
AvAvezYTCZsSSi0HSOWJL+xFwi5RZzykeXS/ihsSqOkElhv4km5njzOWKVNenEgg
5t7kAkE9y2uQ0Jg+hjoXQUfWGBp+3mcTzIC8ZgzS+FujYfs/2LTWATujUSvnV9Nw
W5JI/vn2vJBXpUz1g8MOL4zTjwqOJyK3SWeYDnkNsQzYZ3+AVb0iKmyw9w0jORyv
TTiNDDI802v0Tpd6CsgVOCSz+I0633HPiTGfEZkBx0Jg0xxUkEwFcthQkvA8gzbg
ZMBBE6odH2QYPQj0s46lqKScHL747AUyqBEWVh+uurB5wRhW1po2nJElTe06Y/TP
Fmb2ZqmvfmYkTeWkrqS9P1G8RcR6cm7zhG6bOie/VQwGJWbmDk6NLbLQhrK+4fqq
X1Zj98AdLUrDE2TGSuJMi4SUoxwwD2j4qjB1VWIPDKIWrSuk1M7tZYL3/5m7Yymn
jN6JH4YBZ1YbYgV9mwbCRbcQvlXhuURf0SmdvBVRrwYbpNvdU66z0ZQO90QTx7Vc
Rw3DLyelEIH6rT8/FXzljqyubwQgNnbs8RzN2jNk1A1fglxsabcewFlziIaWNFaz
RFipxlPtCA2CT1wZNFWk3j0L+vXUVnEA38t5Qs1RJsyVwnewuuKk0lLBdg9qBn4A
Mfcj1Z8IUIE7KqFPxyMa0kkuDvgax83ZTgv0UvlO3QyK6fTYprPlwyvhstPD0LIa
rNE/YtSGNV1+uqAoByfQA0tYd7KNmeJYYgW1fBnQTo1ok52HEdAmKcyb0kHt8J8/
zAkxEi/hjivMDG0fM7ykbIGI35YaxLzwyunMe0L2lzLheajjA6Ve+h9Ltam1zoy0
B4nCLDnDklQZWxEhMJcAiYBw+ic03NN9p/1lf55Os2qquGWMODN0eIs0yxSofjhJ
+DwnHp96J1n5HHWmg6w8Sj8hfKFHjo/ABUcerflytdiUk48/S6rZvnE5igU9ibyy
DfdqqDt+IOfr0hqUQKwU+AonAeUPRj2kmPDXXGWrIR1pIy59hzZnIKLkrMH+sCuP
FGeBjeeR/9MTamOQQxmv0PjKTAQXQn22/U57NSOD9G/9QM4wKTJUMYIWfQ6pYPuW
RsZpfGM9R0SCfnXo3S9lZ6MIpq+S3BzskqpkksOqBVq8P/NcFs/oKvjS+kvK+Hvs
mam6Uv+JqxxpBaXqO6VTSsQMKzcgnyNC6zT3TQVsaZpzP29Q2VrHm1UkRiBL5I55
z2xsDrOl/06p5FDgkvhJJqzR4VrNcv8cZLZr7FM+tzUFQVUxkWfqmPlwqkk/geLe
OjuLrV/4Z72A00nP7r2BudE0N5GOH+NLfWclyufPmdgq8ICwHqc0xvbD7O1UZxAC
ytjgoCXDElOJ2ZcSjEfjmsKIZwJmgvKUtCPTioPqMqn6SajUpKBTeJvUVvs+XxEY
V6RZLu/ELSILg4cwTUuKVeIWuBxNQrQzqF7082b7a2BBQoYN38/gasOaUsud/YWp
L3MP1cOAZef5tsssgaOeNWH8+2IcXmh6tFnLIq1772TqqHepIMowNYD8+r6x8909
d1zfHQL6FIKL8zLa3rOs4i7puwZqd2HBepshFXkNJQILi9rWAZ3jP+ob131eS7Ql
dgcula0aNhS4v/5f1MIWzLSweMF3I4aylCWExWXRkeVLhvm19LqGNPi7OrnhvnlK
WbWKwAgrJnruDV42HkJlMtsxmLzZhHTV6NE6UFqWserRkGJmMDlp2AEQFieAENgM
Rm8+RBHAS0yVMYo6JXa1LiaCgmeUsHd4H6oxTFQaDRx241EyNlnov6FrJuv06UJo
YM6FHVfbzjQp6nEG/trh4+Mbh+zpSVHic4fl3R5wxquQX2sioSWQkNl+eer0Saev
bGwZDK3vvLZmwGjuekdw3pMX/LIr8+9WHcVEO/2LavVrWByIDscwz8bhBDNWjm7R
5O4sz8KD0yx0I4zOHfMypvY8YHRrLY04L4Qyu1EBDG2/EjW3WAKJ8trVz/0BM5cu
FrtdK5PDqg+Vx2M/d6TBM8XOdMimIsRa66En2oN2GwyJR7A7YNNnFTtt7QiFTLuB
vecceptOxQ1yDxJU2+wC+qIVJMYp7YZylEVDiY1N2c7eIQl0Tj5+kD6cOmWyKf9m
un7eQbHZkyWJSJTwzoC8R+mlgOdewot9NDQBSy/cMlL1CNHNxRtVdvvkl9Ebl4tr
8s62O/qlKHbfBI28v6OE6zNeeLr0lazdabd3kDocvaIVoIVXqWAZ4lAgy2H8USK9
aKWbcIk5OBHbMBR/vIsKUnG/MU5lzHG0/4OPnblValEDzPDs37IUJ2uWzklnH/pI
+UIH/C3Ras0tuex0Pq6srRPNu4TaRcAtsWm1rqQwF3cYXxvZRMThuFHoUnH6gBni
67hg6c2ScAe2cdQq9t3EQmCNapVzv7ARO7DwjqrjyGahMXF865KdxSo8a1BeCbNA
ZYd1BQ/flTdwRUVenLZiEKJ7mlxg+2vwjhWNzEKIk9dgvebkJ7IVNvsK508Unjp0
dzGAHJ5tFmZJkzGuidkkDDIFvUO4d7Kf3iFq6YO+Y4f7c43uSo3CPqhaDDvKp/Jb
lpDD/B/qaSMLykC237zYI7/MX0Rx5wHS3NO4eIocPqAIFhC7aeSvupbBlGZJ3ggE
P2kopzeY54VLT1PySaLmOjUtCFiwyrx1McQ2LQi0qKYY+Hjwj6aQOphFIdggIbAF
aIEWlFzVKjcXBLVHOT69vjCjP0oOFZvhmXazdD2IIFobpXd1Ai0VfHeg7wLj8Oz+
BN/MRb+bdZ4QiCbg83lOb6xHzctD9AQ98NAKmtHglLc0b6RYFXPmcBcfE6xy1l7I
Vv1fTgvr6LslofDXLZKByU0Nfx2TYzsMsT2sCJ0S1ydUrYD5I19pfRTNDAouDh4Q
8L6Tld8Z+8jv2bGjppn/opDjOmSZRtIYLTHZxcdlncj1KSCP98HbjQ0PFAP0pNCR
SEEO2+8cUb+R2UvwU/yktnhG+NOGCPp5vvXWKjmOMeAwJPjOPuXrmHzigg7eW7M+
U0BEiVd2REXoK923ufCaYSD/2iRTaGhXKjhzBUqkTUxHeff0QeCKnalZ4AfXqy9D
gyXnvwkQEWjuA6SsS3zCuKwk6rHQCfnL9/xAFXOU+JcGhsI4WQU7Py+xZJBXQ6Gx
4YkVlVx1pNsdleLCpnCpp5sgeDMrw5dYGv6Gv++CL4+dqXZsGn355w6Uc4/4DSns
yJpx2W9XswMbtzNaUepzervZi+2g8HoX8V/pGyXLOi+UHHIX5a7r8K1aCX5KKG/s
cpOT8XNC7ITplFQoV2CRAcnH+W1rEpD5EGuOI1nWrzEp/SHexTC/X8m/ue2izonA
ARZaxcHuLfi/QPNv6K9fB0KqfL3wPto7UbAlQVofv+X74QvHLhtgqZU62QJsIMtP
9W4kUc+akMLEvjIZP4fircKD3EqtvidGkabjva16GKop7EORaM/Fg0yi/YjAuTeI
hV6JPWfmaheUAhumeaR+qWT1Js1bl1fL1V0yCtNorMrpUelSmxd8xUrEDZXN7lk3
HOVSuXGH7TqhQO3yBQxCrEqli3ddHlLwvDF0gps7/3u/pbFFYl4OBd9/RNNmi9vZ
8wTBtNY7CBwaFHxtFoVBsJhW+2yr1LbxNhbXtXXesvAmmXPqAgypHTcwxo+XIxC4
9cgRJqO/QgFm/1iIMe9S1ZlGueQ/+QFkwjaKHOmrqijXS+nTOhyo5d5M/4J2ILnq
z6aHzqEb/ZJdQMZGJo5pHdGuL7Zd+3jGSlkurpVrw6/zVPt7V+I5WIkTSOzqh2nU
JT2BYHm+/TQM6sQW6A6SknhNkNeHZm33fg5HoHVV3+yOmsAs8dD1rRu/3qntD9vL
t7nfP0OEuk4mwdhIt8IQJtss3sTjzYUNIxXZ33FsYSsEdZnLcRzzOnrb2PZPOiPV
DI/1Lhi5bOqLlIfJdcD8QXm/on08H3JhWk0uOuJ0602gP533Up97yZq7F5KbFnm+
kJE3bJV/rBmcjF+Ync2z40KR39bm/PahkrxQ7aKqWL0H+nMxlWDrpIoX6/Y+UcNP
axAZABr1Q/+kYasqbTAFyuNwXaCG9Azssw76LO6TqPB4g/5Yo5MuxKewG8Trn9rI
W7pwScGv4bGAtJnhAOMDGgYdPr0wfwNdX/Ht4/685jnBJ/yStmGMM/ZLYA6WfvEy
ez7t/gRJaSXeNnt3Ve+ZkJc7PzgSfnRbu1cKK9T3SnHAqPTChuMVUDlQfxTf8pCA
Onunu8Kg4+DiAmTBByHmLC4I9CFe7JUH1EuvkLkchVgvITiUBgCPT/bjeKv8fhuZ
F6R2WEL3zlcgjZ6C+4RV58L+piiLV5SO8kaG7dv5ea9sznbGgrR+BYiwreiiwmBG
ptjxL+0q4iiREEd0Cdt0qGe7rB172CeXc0QL/pf+/ErOkGKYUI4lgQYppoU40Bp4
xSXrA1AmiqAvnrzkKbIYmguzFzVTDTxOhKiRy4u0zl405FgxG/J6QpF1wW/cgrmw
nd2HCT6R0a+RuyGFjt1/24LxVPnYHY6drCy42ZwNI132DyXgPF9ZFp9Rt3++jhNM
QmB6TfETdMW68c8NSbsJ1KtjUC/OE2lJZlBSdt75rmfwnd7LB96kYIYWv66NkYoy
9vk7o8JXPqPesCq0sJ/ADvB4foNQFUldzzDwSxOTmPpbbM/X6/sunQpPi18HR3Um
ph19t/CAQiSnKLjaqKqrhKPL5fwf6MvVBCigzWn+nXraUxAl99JR8eyAxVVJXoNs
J29jz0bccrghpIYq5N1dpLTRz4ekeaIE7F6tLWMhgSRY73B+nA3j292jZcej6fS8
/m+N2F/bksDoXdzw7V94ZmBF4uob5QWAyWkc4LRtPNGaQ9D3qwOYe1sKMyZ0VgwN
psUyduxKsAsxZAOZnqi4K1yyseA7zIDj32j1ctQ3r93chaR9ffNfDAoT0jqylwCT
ummhRRTtoQBVAbPwbSroNmfVv3RtXqeFKrAYnp1uCKCCiPXBHYufQsF4VaFFh3+1
5tVUNjn9G5hYgC6JtIF9mzm9nS67VFjpuTYVAr12jwIxOKBT+qrJzBO569RS781L
KwcU4TFIVwSVfTYbWfu5f89+T3tcguXYVOWfX0zPT9/s6kZaPKPJjJSWvyH0evbo
pcZLT0UpwXOF4Ye68VwMMdgH+NFwWE2lBvMgXPtCUYXtLeV4RJ44f1gdUgZ14VNk
JcQlnPpFSiWuNLhYRdGCJLmAMxEg03wdzI31HbIba8Q5crT52Hh60AU35nL5LZ3Q
AX1rkjLIthh8u2KGAUlRCcTx8dEPgFKQviK7nk5LBYVR84dW3uHOXveywVlhEIBU
eEkRV6qObVw2MlN5DCFIEsGQtbogbjoD8TvYj92tH4zVaD6sekmBTDUWccpvajFQ
RbYjtaXMqx+XDWhI02Xc7VRpfGCOxs5P2/SnSlkTYxqWG/HNaOjPOa961ItHpjTz
tIIaaTryvW2wecSY/y4TX81/kMwok7z1otnxyf2x2oJqVoX8FNuzGMvepoH53mQl
p4LhrHoa58P5bcQcmx4iIzTIslJll0w6/L1B8zBk4efK7W9GGt12KA0UHTTOIEX+
uaj8ZCYVrOg+q05/6xvNHq81IRMF9BE8cVuXC0UWQQEbefHUZvxDibIRqJn1kNzs
8RlfuXaC53G8qLk9Q0BP4MCr53QYZwHPmcroFJA/shCFmSR71b9jdKnFGIBhlYHg
vrD1RYTLxtZPnlFQV8+VI5wk6r0IlUOGko3S6e/BwoBjSIoFSe1GeGOmAvMp3gA/
SzEBrp/UKxs1F4WMFWW7jZZHLuWKF4D8RV32n2uTjgux2Og7bdAyGmYaCOkS+TBa
9dxjrEmB1it39KQS8baMVxsdXiYQFATgoVWnM61owWJpUKTLFouaQ+lkOhL+DLC9
SuN8ByYvfNJT/AChofVKfy1pTfpYppszNsVDPAyRpaBmuQvWdBDyWGiR4zi5mvAK
M33XJPupu+hCZ/XUtCE0jMfUW5F3oGiP7ky2NV+MpP0reyyAHlS9W0CYWcgtHpup
gYFPMdK+A6NT1owbQnXQSE06BRb956kGuViXsDpvJBfI9j4hS0yqherBW5TWEVhs
Q1RDenUHv0tNHDwFMMH7fztwJRg5nj/QvICI+S/0tDuZXLjHbWSvYbv6hqcj0G/a
wQ4ST3ZVTGtoBnwKKOu5xJh2kNV/dZvgHW67GIpwFHW3WnCB8thBjdOmDhGSHY07
05ZDqmxTxaqrZzE3NhTuGyMJmguom2dVQTYDqlnk5KcNXDRCOacZ1BF3T+v4dot6
M9rNbneJW+T4hFpUrKMGzD4SGfwLUsJ8PhfF/DEDt4Ff5sSO2uEDNU35N50Stx+w
OybCka4omsHE3bGfQxQ6hm2azVA3de9+Zia5Iq95VMMxVteqZ8NJDNqtHDJAfgO7
OI3ppIiYt8AoJcFkoJs+DELMF3/7Zr/1f7WaWHI0/yu/bUNnJW8NfX/JgAVTRMPz
tkG8BPm/Sgq3xxogZ7Sm0lhUCbCDKKuyV/l3iB4SgfieKsmX0T7Yik4WzKH1K5xB
xvF9X4KSyraeG6GLYGCwxNsrZNzi86EQNoxs5gTOqH9TEaR8yunhcu3NbhS8ef1v
4B90r0M2fXLQg99Wud7XeMRnZLXnUQjy2XMRzFvVbhkHAZxr8ZtfdmhbIuRLKZ/u
ipXrV2DlWVx2qPGLSheRvtAESnEP70f701IN3UR3JHcx0oGo+/BrFY7ouIhqY8fQ
B8Ck/uRnNeN2QW7ez8bPeCYDDHbf3NLcOzEEGKjZf/xMO+LpE66q0zeInMU3ryVk
pxgMSIC/IIkrlqMQuj3bTb5EDFaqDoDRKHlANrOT81p/1fEDaPQzDiEZGLSmpQZ1
GdSJXLAimQrpvNfCVhr34Y4n04ew3t/EMeFAvJlBijXqJY1Gwchkyqk+iJ+zhg17
jwc72AFM0nGEjHAdFAEhgaSS/IpWRZiKGZo8dst+znkKSj3oTBRl0c0P8rY8vLuY
J/w6I4MptQRyQJbVN5eimcUVi9ZhxZ0HxZbP79b7o4Q3TIrx+0rbjnqJ+YjwIjn5
3Gzj9GEE76TUlF1Jp8x4SNQzqu1Ccr5IQiAONpvowRcVfMqSxGMw30zMty1duIVO
xzQ4eWavkQIcb+qCry3icirv03qeVvef/0GVjk85ipuKC142clhe5iC9c0ggJGLU
N57OmyBfXHW64YDrHY6nytqfTV1BA1EKdmKRrYBkAIlqhCjI7BPiw9r17eXThtiP
bTLjkqdl2q8vRLoOIka8FfUP4cAK2y1ErTNB8Bryi6aDNndjxgMqXpFYxg7WFvMw
3SO4VUrCk8yHXMX8mKh6g60OgLVMa5yQAetSz6shoCqBkOxYC0wPt1UvZKjFNKkU
7VPpHU1gV0T21c2L+4iEyGdK9PrcyMEglIytGRz9jXKch8xU/Sd6UIdhoVSRwIuF
Id4I0rcX0WTA1vvA4xVpKXxIIm0qidjF8rUFwxrtyGzeFmMTEdCcd9RvCRKa6JC7
s5LJhX8WK2Qade4w6it1GJ1ds0+kV4kkLbROQabrNHU9kfunoempAh656Q3ya4AP
MNoOiAsGcrrNW/IJ/Tukju8ohlOkvmXxC64B4GcgiD4i0Xs1Wlen/RDo3j1M7JZy
FpQGJq3OejqssKCUuK/wYX46pTtuKU3c8Lt3LE0cypt6S2uuUxwt+mcNQb8EPa3X
d6RIFQPht/D97nKk7kvP+02Qec5robMUHO5/x8sS8/KwgZOqwzrId4OIU/nr6Sin
sJSzFIgVzAcA66EF8THHNUX4z9Oruzzqo9pulCyquAco83rjkcAQvlYTRR+CGHJ9
j02JO/Hk00M6o8zc/MAQ8iVYt/qSLpQHR0JA022VYfP3hBeN7bigsroypKeX7u6U
6fwKS+mFFvf0SXeIYYuH6aZ9CATfGnv32ccgjVBRYckuA6dMkPZhY5hRunGqVVuX
5XcCwyb29hmwATMzjLv5DWqysocXTQe/GPgDnFJimmvNofAfBuLvh2VqP87ykLgH
g+cnA0lAuig5chsqx22B6nb72zlF1/hK45YNAcH/Jmgn5di7EF83anpCO0dAgBut
nKcczK9dOlFrOO+BEBuvn2zwqBmJrClh8Iuf3+U7IZF6gwtVbV0CUxNWvKvELUCP
w+Uunn5B2PFoy7RcaB4uvemQkZIodfl55F7C7E1VcuL3GolcYEWxQTZiyvB12cCG
XZ5B3WXotNqnxfffME8EWM4ZmPSYU3RzOy0lxS9cngwPeHTxhtcQYrlUGGZQtirC
1P8YgGr8globChRpSoxewOhMFpGNZTGGpG8GUS9gC1ZEq2h7l43LfnPy2/a8TM5q
Fu0EuKUPYkjtMQ/M+W7QA2z/BRU9xMQgyH/TM/j8m1ERNGBAYh2PcUmSRTGvx+dj
lsYF252ZDYqSr/u7SPocIRx/t3acJ0xrMC19+whpueQU0Pbtmi4WfRrpZz/ZvRMV
Ov/6udWW3UVSdm45f3vz64JQQ8lbN+9X6nDpu7HIeDJUHcYP2Y/LXMCAVj2Z5yEc
4n+2K/JWPE9sI3BrX4XiTgRML2dzKL+Ez7ZBmrp+Z9njHHCM+Fjvi+D6878kw2hw
ck3cmLN6mBIrrJ6DKfD39QXVrlkgcgZCDEdg+srGZNoV514tvTEW7ktNDncFu2v4
nZdsvDNw7vlf4nei997WRcEdqplgR6hJsRxnOtHwRHiSPqlWsieCkUAU8ZKhJfla
HSAinySpgoc35hmXvd4DKUrwD9xYhAfzZMcrH/TowRk3WdTgk0OMvZrVQBhd5mo1
zgQdLoHuhLCa1mk+CBjRwETTGupyTXE/8MgYhZNPILLQHXDdHDrIbzWGRf2Q4DIY
Y3yY2yR21iCrvtDA9iiVJXaOPir1CpchCtVwOyrvGzCUj2r33kkpZCJikqmV6UFK
dI0obq1zmTxkTy78VyOxM4OTzBzybTYIwxd1Am67OuhlYJBwRq9JN6cN3WJCnZxX
vomsjGlsGxDODMGS+ycS/4KzgF4GaNJ8bCwobla/Go1w9NrE7DF5bQj3IkGscwPa
W/Z8s625r6niQJRnyYh5ZLhuLDuE5cWZ+T2pEmqK9RQE2zhDFvg28CxQfd3jDY/y
lmNIGzHHY+P6gkysezeeComNMonHi47XrMdKN0JroXZazzJH2FaV0B/zChm4WtQc
T1OTqguGozB1SLx/pW6boSNN1LOvvcPqOnUm25KpFsN/IUqB7NAQDSTVOUyX5u6d
9mNGw8KvVOfD09RuYCB5yqyXNudvI5L1ZMG1IwYLMNFDc4k6t9qGap+EE1XUJFTz
wVzCtxeQY4WTCzImkexwiSmfTBbRebMrgWnU0sy/aI8Ws4ySKy4ZH5trJZ6eniix
J93PFJcMDAdRD1A5uZSyb6GS4k0uqGk8KeKzKZba6Hclh3m3f3GDNi+4i1SQtNQz
W5JA4lVDYU8XF2tO8lkU0CaYbGjB9t0eeMZmQqzSV62STUjPVEHtWKFvkXBaaQAm
7DnVOOx1le/mABeHE7SkZ6SU2YXPMl3aH+7YVHvH/ksqCUDI3vXlGFl8yRximKwb
WQeAp6HsLWRsdKe+BAxXtBkTVVe5lH8qEuVPqsfnV4TqVZwLhv8q2RbgccIEy0JU
bJ0gNUSVQJ3zVqsL0apxiFYfjJGIvLGfP8cXYHUys/DX4L2c4ophz8l6Ll28sqdh
MfOiYZt4S6v3VcEDy/AsqHoe2rdFXb4ellg3sZ4YKOhohcvbThY6FkIroN/0ABDN
C+P2X65MT089s9H4aBO8LxXOthtgCzgjXCRel+vAYUFhnIvpcDkmr/drfcLRR3lV
DIUftLNY8+d/7iP9SlhqQ+k901EhDQLxQ0IK+k8LlQ9CvOyp7bxjOYzQsiQYJz3s
GYLwAGH4yyli9Q7YrnXuaXEpfvClIo2RdHreC2HPY7rF7q5BEKnko8aaPgkMKsOF
Trso4xR8ZTm3LLSkjijo15cGA++CX1ck11ce6MNzA7DHJokyZcqzfNI1AUKBUwo0
IeyE6WOiUfqfYwDrVkW+8+iAqtA67PFdZPePwmghiTwXAYb68btyK8HD0qyYNrvz
wvlbkHlXhg2VvwsdKKk66prZ9uxSCXvrEdnHFR7Wgtks1qwuU7GrmdK7+Pxnbfnr
vwbs3G+EUCuX+04XYfFJ++DtbdWgoPOOse1PnX3RfYXTUsqArKTbhkH6J5Q1op+e
Ji4tnNm5vj9esI6kQRBw0o3yY7Wbaw7IEr5UVdQxbrT0qI/gCpQcwyPENRffeBA3
C6AJlCcXKs64hEbnpj4eydvVnw8huJpt0lF2Msl82664+svkrSgQGkmiD/LG0FME
8BYuxpNyfQmMorverb8NfmFlHYV+cffMOD004cjHjWkpB95tARbncrYKEVIL2Bki
rkzv5g61FgKQfCbqCPByadI+MMgbqWkjBaPmRZsGbDEIbAl+9U9iDI2eHXv/4Fr5
v8/krVz4dDid+WOP/4jR+/37Qi8ep0HQFsfr6al0j8OJqEpOPY/vr6kbxkHXLzLh
T+a/HBE9v2kpo9bRW+/qtg51lE5IS+k49bt2gzLa3a5+YMknT1/XH7MH5b9FChir
QO38MTUZ8DyBOK7rKHAjLpzAMvjEnxTmDoc82kkjr69tX6or4IaEbJwyGHr7uFyq
3UUtnVoILg3DDZVfS8pqqNRvAN0qBBeJJXVMFUlqF/TFFi/Tkie2Hi3AxDv8bhHG
pLXqGL9AyWD1VXEGFYRHlLAtLt9e4CIxXLFFUkbsQ+f7MHVT/kcQm6nxzjer0+8F
hiieZ1nyCOdfHwYgkrxebYkqG8QNEBKsGJx1rvVTOc0Fi0baxi8p/uQg7O9TMUWM
5B7dQEjRgTrm8oqb6156YZswQwa9NyIlP0LhcS5hdM65Yi30lF8Di7GPGkzFL7iY
kOwwB+PQEF8ch2JrUgsirUzdLI2mHSyJfayadT/wp3MaAmNLV/sDPtUfQ7pBVqPf
ajmZ/6mnf8e2+ds9aE0GJeCMNUWM593ywJ8lQ/oWmezYq6VUyez4TWVFJ+84IbJk
sQdrh+MaCrl5PC5e5wNmkhEilFVtEfFJtgiYhFSByauUYojSxaXNU/kWXgrP+Q+V
1mhyK17K/Gm7Dqp9bJt08IXkhO7sbC95v9FqARVQHWcp1krChBaCScTVLQW17shU
m3HoU0QOYXXeBvfIINTtKBevX08au9VUfzaTU/Zc2ruLioSRDmvI8KK/NbX/LFaj
aPnCe2vI84kB6uX9BkfS92RonIzlaeGCReKkojuErAh0M1DDqbVQCjwySJoz5uPR
d+Q5R+e41YEiv3GFYIRW+MkK1m0jO71dDVsorpmZdBa9GkbIfuU6HHZd9Hokw/BT
6bnkJlITphj8uAkVerNUwW7t+Hh92lcdlSy6Wgr+a0PIEQT46IqCEwr7abPGpCMf
MDEsfb1fKxEslDET6Wq92Hn8LwfPKfHDg5hcGEDMf/ZuuR7SpkhU2dL1RIDdO73q
b4CivAfnmzcScKQAXaZcQkcvG8UZRjXUUfiuY9YQy4VpicbbHuvkKqQaCh7Ux1Y5
iYWBtxY904oYusBnxi211y5H5BZbKw4o3g16yXOmfFP0l332D7GYWDLHKZYaW1BC
vtwQ9IzlR6VN4IQmD64v7oUYthJcJ1Be0ufOImgU2g1fY7Joroe1wbvxebV46T75
8sH9YKwNCRRO8dLDuP0IBbAKthPx/Qwq4JLx4bdzmoKNZJA0z/mVMGnZfGUiqpzL
USdRT2ECu6zek44l7Yb0DbGKQXAdf+5KibrFdS1XcfDEPA68YOYaqEo/I9V1tUkK
k8HkTOrv6YdWELkrHDyylRZPhyVBJq0/zdx7ck3WfZzHMccCwt88MO0mUh7EymL+
wibJUIeqBwPNnjTAgN3INplQrdA3ZhBtTqYl7M0vXwTgLsuWQnF0CUHdkfZkwk7f
lxAYMmA2uQJLPg8JMAaqRWNjBT0o9kFvbL/IJBefV0GHYJEj9nELoou2yt9iy0ZV
KOwq+3JPW+323EflX+mU8cq3iUd0Tx6MuQwbGeIVwOLSSSLxooz8x299LXGMl3kT
DkWqPeGdYj8x+uVskx1Tj2KV/zhqd6BL4vLSFsm082+4iDYQ/w+6lKjGTRi131BS
5bqC4DKU81K/G6HQREkgG+90s+qjsopDvqL0kKo27c1C+NntrCIgh2y0W67RXDNN
v2E/45vkJsdlCGeyn6fEi2ul5lz5hahyMnlakJ7ygsE7c7AKdpaHOhXc00Zi733H
FjFnKjLLOsIbNFazhJqYz9dE9kgNJdv5Ma8DATV/k18KKEc13/3HCqhxC7ORGdwV
oNKNH2nOIDHD8efmZvtalSoWLpz44Kdoar7aBTf6lW6Uy5i1RoA/XHw0V2fFzvSG
P8V8M+7OViAun4z93rofO6XwbuRckyPGyf1CftKFaT1OLmCxT1TNceqj1els+HoR
r7l6Vk1CGhqhFQYmP29cY6rYuOhG5QYXTH5I/ae6y42UPp04Vvg8EmIaNP44zk++
6cPCTa85z5Jw7J4q7x1H1ndB72196t9dULztr/6RBPHSANDsZROuv/sItwgl5O0a
NSrqbEI72zHhL3CBZkBiB+Tj4gsnZQJXRIavELuumdPCYH1ScB7NstCXa8EoP2hd
h0jPm8z+V3SGTsoYW3gNdmrt4MKxISdkX/FVxJkMrugjiwADtne+W3PDb6htX4at
Yf2EbuKg76DsT41AhtH4/URJTIz9uBeWPBcR/2WXVzHwseNtj5zp+iyqAnqqgUP+
x3r0j4JWWISiV62Mi0eRKMbW3pgz7NGlB1O6zFUaNNPpQJ4y2cjnIBJ7TunoPTae
3UKgllp+9h3BKhlkHbssT95Sf9Km6ot6Iq2KRBhVHxQ69Sl49PqeMsQGCtJ3KLOl
4eWpnnEuFcDRBMazXKxh66C1VDBNt8EhDVZCqhHEePPOUv3qmRoqFmbXdcDs94yq
a/t0+ldhjMb0tJFk0LCKjA8y9NhOQVIJpt6iRjKROEP13b9ItG3nlx6FnOf53sSk
6yfaLK/8KgTLHQxrxfK2Y6r934DgkIdeMHkOgwPNHiNCK9dbM6xq4XUzwEjMq+vR
vvjFf+gCDEEv6JvVPH6EMWSIdMlP1rjkW6NRTct1T+AGR07AvjEaSi46qK5bmYuK
GHPVzQlT8hvXpsaErKQUujvO8ybfMKu58ZWaaI02p/XoHsG0g7KnnpSb/evJifXx
HOv9QoyBy0LQ3+5WVMttj39+5qUy/8gtQvvMIYnXyqCL+NFLIhbmbMCXheICmlD0
zi/l4aq/n83URLKW1JWwHr6E42HrUB9R3QXnPJ+GHLE/pZ1rvBRH4OvdXsg+EG05
Hmz9mERoaiVEDYrA3MBot0gXVorPz9YVtxWOrEZOzvSRoiZSeNj9Dl3pep3A++Wx
KEKFzn3wzKG7NSuwp56zJnHSs5TSflWnm9+VYBGV/igfTmcZLfoEmD/DwDQg1jE1
J/635Lv2Y29/h7P6XclF1aBU9GTjrYGfGRUlQTV2nroV+OOzPGBm0x2ENapcmw+8
LzSdncvE3D9yhz7lFmBHrreTaO4qYeCxgUeHqW9cSxHRvXQazdbMaNKczGB/i/EM
kbQi32skCk0EOLvjGU2fyqnTRJNUTxmKwRSKihy88x6A/EZImPEU8NhAZKLQD4DL
beyg6YrWPSS2xFJbdJAadJRcLNO1yflJy43n7D6BEaFyDHvji/+4WJe7/UBxWc2g
3qCKiTQNbGutxt4yom1XwdFRPvoIxOqvpQ4ZTHXzR6L64pC4rNqFW9XxLJctO+gy
jr5Cxtb7OM2taYIOiaMEd8ttCmUiekIGjpVCgr7yt5eyEJ4qcxnP2HqnGJiDcei9
9XwnMXvMBckipWmDLHXmShvSqH1oz/S+BOWsod+Tm2cC6BnjxP6q185lBrptLJGz
6EdCj56iNxPnIx+vtjggWA+bdzxtDIaITmlVUuWpTYOg1PgIrW3Z4lBjg7EMM9Ut
xrgb8pXvzK3MRXh3md4ln5g+6osMT8jo0r0NBtywYo/+P0pnLDqitpCKj5lnainB
amRExpQIir959n3MTi/S5tdAggmbG1HlCxS88U/x9jt24v142S7fj0tjzWvtNbXY
nVmwwz6oqWLTXo5VCdIIXFWMorLSYqKI0k7oJDABm0xbUCaLDMi9Dx3wIjrdddiM
ijHRnlYLpnqv7jcqquLr5cZCWW/iVFA9xyATlLtUyHo6dyTZXE2gbQ8XQmuuGUFN
9C1Hj/Ntnzj59QA0gA+aOPWX9ztgebDV/Op+UHIWRUvYtxT1Nw4MpCIc/cq+/wfp
wBzh58uOBlDccAy59eE61T58S589or9Cwn2E0gLrc0vJSCmxYa7JAWJ9uXZR97s2
bdXV9ebGKzvXNSpBANTCikSDwht3aDnVeDAJxw5xLVe+8VB4JB6o6wHFvGmTC2T5
Yz1Chs3tz0tzSaMXo05vrhVQz1thlJZg4o0jICbE9V8HV5m4XY5BbLygMSn8kclB
6oWuFWb4YMPhd7v/Adyho8NQs2IMPOywMUrfEPR1ZLxc/LqBB06fsCY2chIq35Fq
+hrcef81CRszmUDDzl6oSc/ELERU+kISo4/l1X6OS/sqM8STLiG15d0bkZcOxg4Q
tvRpT4WZIFZJmG7mmyHxYSAsjucuYN9at5tO9dWzfuKlUX7A1M5IOv5Z3MkTddZd
i1f8E7Xg6gNQesrj4lV0ZdkoLB/1sXrLGXqQnCZJ9rak6pj0+VUAJis/ctPMwIdL
EuONJCq7JHdOFoCSZUrxaCyWxH7z5x1UOJBfRwtNgHZa1krL+x+AJJ3abHRzWoqp
M7gvgXAtoMkYYJfjf9/UnGrz+Fgs8dIDsWdaoaSVZ2++7OE2pMfeqHvq45VTo98S
fDekjRrpaIdtfq68f3tuUlikRlw/HGvdhpGnakDZ98Z9dx4ALBKDraIsLv2eWDsT
kJykjHrxwQwX8a/rLMgEF06pAwNIVsLZfLu3uweVuENA9wIN+NwGcBKmOesFjVII
HjY7L6u5bmfFL/F3XQhPBRd2TkkWjXyeWt5TnI4bF65/3D8229Z4QFCoUoAWdWbw
bgGJkkRWWiWTlwiArdUhl0cHWhrmCBcF5REPRcIhJ4j2jqb7LJwLh3HM27Vjmk3V
VqeppZtDkkruuTDQ2v5GgJXrxJyIKJ7qCcAzGUFKFI3w28VNaFSHCiRwpTxZ+k1A
PrJtC/gD0hdx1GdXxofX5/hZHHE8IGfoIUftiXSLrVKnznm/MsdZynu47Z7mb0Ok
pJ4Dz/DYQvOjI9Yp5OpqecoasY0HZ3ih9ce10bPCEJ93CUapCyTJRJgAjhfX4BaV
8zXk3NQbvkBKVJDBJWhaMZmCKFNJFh2iOuHdS1NzHdgyhIOaVOhQarzyp/3K5f9H
S7Yz4OMe5D20I3evNZm5us8xWRZX+TXdzKrgSLJV9qb9JdAO5ld1JJChBZFXzVbO
jqErIj3mJ2XWAq3DSlQzwHH54Tq3LyFqWou8LZwCdmgXmDaKrGhcHBB1Dm25+qv4
5zqFHcf2AIML28X1Inv0ufOKLUfOkNpMxzeF3dJ7dWqbt5JldLQJvtgtRRZU990n
OrJs+mJTgygf7IBBT/+v++KI3rZv8mIisg7MDChv8ZiD2mjHYujeqZAB0Wm+d6b0
zSqm6Ux/2H0ReB92xKrGxoCdUCNVtj4W9YaI8EVaYlQJk39gjWAix/lr4h1tMXgv
h40p8FyLkQGbEhUiytxMLUeNDsOsI4X9wqhInRZ7UTy5FGoHHlxTj9ny6mY3phlU
LLAnix3ApQHpU0V32OIL/akWOH5q0J2oXLtkoA/AFpc+HdTYWost3LEWFR47GgeQ
K+sdMFb9v5GUQRlP4lA1m0PIMsuZrRfgPcV570j8CkLSrCrHRC8a0kXMrT40BNCn
iMHA3dwptwTMwKzqCBIYSLhDIAfuN3RXRkQ5oj99Pu/ouZyrvelDCd3AGroCDB/C
nzhgXuJIHG1ENA1n2QDaMXp1x5dqUSyabEHzDGdY9/z5axWoF+KaVhk0WU0rBlDB
FGsv7OicI5ACCOOJigs+ntqIKgXjeGN9mhqhnEzQ9nqHRHr44ElviWXgNY2KExyT
37AFsRAN4EAySXriTt44nze/QigANDzu1FxTCVF4uPoABqv9gD/6+9QxzbEx9utj
q99JOyYlrn3AB4vBLcbRjUZwrK4Kmjxg0J2WmcRaNE1iJvEkluy0LZoAsSLXFYVf
KDtNuy6iALDg283WiqFK4uG7XqAEVB/9abBrtahhDziUgujrPb3qbYggTuoguejI
8YCLzBVcjyvgI/L4qMqG1ROk61ef2zlKKi5C4bVDKNvwdkYG7ueJVJ+636GO9P1/
i4dibZP+bJ1cTnV7KqONXL12afgQdsYoAjVRgNoNqWgDkL+M7I3l835yYjb4LXLw
qv4SfOKEP7h55Q+zhusJDHAAw8JK8Q5BXAMRpXJAoTOyiYGR5QWe1BNvoQq9Yglx
gIG+nqL4aizb5uYMcqFubu76JvN44jC57MBV7S04OWDi/wTF8qaGAqnN6M0EYM8y
l7Bxn1S3XkLm4mJbizUSwivs/s6CUND5kbS5feJwrDhfAbxzHehfusztwwaDNmxm
DlTCw/m97VYscJhe1Qjb2R5zOAzFi6vVZZPfFdKW24qy+sIKm/VxRQ38eOOCZPoa
B4SqqB0G+hrynfdjMenjjMHcGkHp9eAQ5Qku0NL4sQ4UHT0g0PqHX8b2+gI46nNe
r+kkIx8jzjnFn3WXM/n1GAsB1REdh3eLssqG34/pCH9fxm9LNjMdGo+/7xjHJdf6
D0I6c2zhjNmZT6roj3BehyfHHXn8bPS9CeaXt5Ef/IIbZkKlAQzIRaR4yfVca4Q9
Xk8411NFF5PjxDHUBed/7MSRFoYyXAf8LXNPIJ7byZKpqpkYAkWInIbE/fo+0o1m
V+o0HetfxKmxu5Qpra0ysnSsqvGAZ53vvFkQ75LfYRVWOJ8tptLaFaGqMgEcOMY5
c8Vdzzz/3i4uM6v0syCyB94tA3YgedNQQA5xB5miq07uooo/a+64Tnqot3EUIPGu
Q2URT+uefatqWUnQgKaEG0vDItO3vMeB6nf1nil0/zPV2HaFllw0yC4cqBD2YLLo
OVFeiqDJfkaxzvLwZv7z4mgXnzQpsFxE3kHJYxL9pzFsy3cIs7uzLU1O3MC0FvUB
1+6aF42vI7sS/MPEhfFdiYW/XNEhMKVykCQa+URUAeRnjwFvFqrvQ0FA936sf+A6
+AgooR7cwYO8uDEln49YvnoV5N3PqTQNBouLnmq2X5fQxbzk7oY0Kh2dlqEF2HRv
QjGm0wEDYHF020NSt5+2aA8hArBDdGqMOjeeD/xZg9KE/jGNHYCIWVsL5GYkXQqq
iyb2QYHbQlsOhPSQBjjLKrLG7IkY/+6DlrBrbXdzHz0zPYJM2z6o/SDFHNUAdLL5
g7HYAxJ+QdzdCdeJdJxkhPH+/gvv07CCgDXwIp0yX6ijTCNyMZea/IR/OBeyR+aS
Otd0NK5gV12BTApkcG8FQDRlJ/aEymh8OMrjirgnRVrIp56PFaNzaP2l6CDY6DvS
9wTF/APToIvegBzV/HB1aeq2mKUZXZbIMIehxdZR127gseLwbFrFh5HFxJfvQop1
mngoRbfLswufUuwWmuY+rIULMHZdZFTArSofS9g8HrpkI+HP1s0lv3Lj3E3GUf2W
rtS5Hi4y9EUE2xa+YlYp8a1j5NtcbWhFXxTk0etxJP3ru0u49mp+i+puYh22WL34
c+OkJQlMhBtgFxrnJuSHKGx37zB0QMZToQbBKPPzPpYjSg++SP4jQr6o9KdqgnM7
q1o1SYMG+mLZlI7f3wGcg7DpVPKYzaxZ3yXXbnzy7B/QsD/1ryk5gWB76TNSax8W
5jrb40l61QzD+FV2cW9CuU98IWp6iEoIZID32jURP8sE+/3y+bRppD3gLmDeTI7b
laRRgt+FwVZD4Nna+wj/seVuX5bXYdNUPFqAW7OrQYYuwLdlxcYoruWooXhER+aK
aW+2uyvCSUVmTX/tWYP/5TVgpC4s3jHiGFvvJLqYV4QeOASvkem+eBCHZ/ubXHmG
888YzND6sFwcJsWTnZPWYLHt6s/T/qdX7yO9eV94WghPsa6AaA/JydRGi/ntM8Re
ZDAe0UkzzxHuBCNzMYTdNW3Mp15RKI5tSaNumcltcPOwFU1qAaWOTnwwuTTm5hyR
OV3pgqqIO+ErXAiozCksEd3F7eRyY9BfQ0D/KfPietdBsi/jeKPyWq/Gw2UUgxZv
8zgCA0TbcfaqZz7ZdmoM8/IpbmqMCKwiPpNg+1jQXPkOOaF/cbHgLCf+G31mSPJy
DuW6pOmbhE5lBkd8DO2mtvdUgeooSqfJ90qSOInjFkIEG+sJe7pulH6qjJYxoxJ6
GSQmW/nH1i+Iy7pqX5ORQEuxm0368XfaNUeC0xTL9BsIIeGWDUkaJPSEhbZkbroc
CmB53gm9I87/FRrokj5gmN1i5BAjSH+FjzAibP2J30SccpUESiolAlasFpgqE4PN
g+i8u3GMikRislIU50h7VOJ7hamX3XCeg6yksk506oDLNK3GOGWv+SMaApBa3jZU
1FMrIgimVGJaO+AbPieEC9+HVRo9NIEpXgmPOCuxZtHmlSa6J1DeBtY21CnpgMk/
1gaY8wZUDLhsop5CT6MRudg+JbVsYdawkNjXCX4zESRMe5le5j3A/8w5dQQYuBhI
hOnMp0NMG/wGNcnWXpPM2IZQDK9GxYW9rm3B5rf4mvEM1S2hL0O79x5yUb/Z/hc8
SmkPxzxJ0L2N/n7+8J5ZcvuwIPln5YHO8YC7EmOvmN9TE4TRFqLZRZPS0fpEZPFQ
pdMu+wsHqEDMypRzEnRJIuTeLbL7InptcgRbbKQhuWGM4e6HSeQSS8tB0nhme0sW
gJFtkPAWJzfkBn1pF2npcBvIhckD2+lxS08Z1QUqH+8VVsQw88/t74rpdj4LXp2x
uGurXgdGPHDiboGrsLRmgWGzJXjsu6RkWYDVAPBUNQXqgm7DcqwjIl3B707hVkYQ
d3iO0Usxu3sTGTjCRLLC78kiyNVgocJF+cru28z4yp1UFs4btM1pyFOcdhTm2kIi
7iwtUiL0xU6NhoylyxbEXHR6SP0kFdIRlLRClu+H4PqBY37iraI0DQC0Utk9zpqN
EjsSuU87OkilTsjc70mjkSpuL4+u4CljVqkCjnhIr2X3qfj8/sQDq1aL3uKe6y0P
RbUiKDKVkqHlmA91oHFXSpMOkIs8YgzScmNJ//D3bi5/gZxeYkcutJFb4021ylty
UMspxpJD8gdVl1LAO6eIv20ps5HfHIrienGa8iOkXt9yemZSTarn63NVDi6gqizZ
38JdNjyCiSMU4DHP76q26nSK5TbV4UrU9w+zqOn6p4tSwytj9JfTaVpcH70vdOws
YgmtJwbeVdsE3JJf/4zOX+VF9j8oKZDfYNk+c/Egke0YXJt6O3fCWMRyUyRmg8+C
vs4/8uB55AssvBay12co6LExDcRmWojL4U+KYLQFe1LBXmKTwoToizPAjKA0m/kC
STGBoDpmw/VixqUSdUB6femr4lvYHEZfFmEogy9hG3S0G00Cfe0LJeSFUjSLptzj
KjkrKEfqPEwB5PgyPT0jAhx3r4O1cgesjCKSVbOrhHDeJHqDuBwSnE7ldSviuoyT
L2a/9AXZ+/BWnqeWcvHtKxdCxBfGOZNh5HWvX0LorIslma75Ou7mojQpLKyqjEGM
TMqXWKL55gnifykxXY527s6b2OrJXszK0W0mkQS56PprO7mI+D6iiiJAJmIzwDkf
sfTDO3l6sdGqqmJfjVzy45d1zDPJRY+8RXXK+Gns9hVFpVL4xNHPBRaqXktL+q23
jUBBCEQnA9IH4R9ggytr0ItUqGfMB7cqp3fyC3MXfSTexsw+m3CNteiB5slEfjZp
jMag392eLsC9vESFs79S3xlLqXUDat8fWym27kvX2WCSz4dFjW5l7ErUfpGahQJ+
KR42MCcNVj6ADh/nALaj+Xt967TagIfdfFeob/CBlH2Mpz6LII7IboSMfjaCyLIo
0rCA8njzfMCqnG2Fh0o6HIFgvMGAZpTTANncz1mcybZO6fGoR08gBsgXBmwV0BMH
HLeeQy1dzTI7m7U1jG59uvXM5UrMtjecNKAHAXdz/q8IiSgNTqDZvOA/ZIp8Ar6a
fCFR143VHmtQzeI5eDZ1Hj6xm9pUWV0V+e3e13eXMljXIBT8/xzNkWT7wKpcUDGU
aiPwYziRAeoBr+HrSPwwTYBcaqMFh7usQpLa9W5tfN25zZm24SAcmKzdszyd5ikP
l3PDdSStwbIT4Y4AlAWex4kpwj8JD9Z6dOtvIt1GEYEVF2GlqMAx7kfxkonzya+7
VxscYjKMdcaBRIMCQsMO3DdWzBZH8XmVsnXCcCna6RKnX8rLPtE/s7hTF9hE/NT2
pj81bazM7y44Vq1iQQKn5tAl8qD6Wc81pJMJgjlzLrCtyXujaK0j1sJtlaV1DLww
HtLzSJB0rZ0Aq17sMm+5mL4u5EhLsIUT8kt4kmO7qSNJqqth9RWxhsjB0hItMfb7
bG14HjXYOlNO+hFUiSB4/FzKMqxTegqu4FPE7t71OirenGIJNpSrcYmzz2cuXcVF
wwLLet/UELc5E5q4C4vH7i991vsA9Qx0cL9Wml5Tv64YVDJ6VuzEArLefYCryZIB
hbhkwvpBzzn4XuWQjs9g7XrAIH36y0liGcBxH7p9koeJUlk9TqLwEEK3gz/1RDis
uwfeRogmvp6gJ1yiiLn55KhV5i1gLytod24ER7nFiYmMjt4kY4oPUeiXgyb5aE8M
s1DpsuHcIuF70i3gpcGsnbZlf0IlWbplDqzaPB7tztwtULfmVFZbFvU0sZMJ+qIt
b8TfJukdGUJkGJzN9q2ZW9KcZojbnfebRma2RqAVULPz3qSRs2o5Ed+3mUpNjgPQ
fHMCoKjQ0BH3Z5tIkgR2j6bCLrYe1vOB36tR3WAIiER/W4oQN3kMlCMhr0+uSeDo
/u7+bhYqxY4D3IpiHNAgm1LUoLApfq4df5VCFZ56/NebMvVM/k0pAyxr5mFKZQPm
EVStnuzt4QnZZlLRLV8tRtt38W8gh3ZQ+ZTri1HINQ0UIfGnkR6uoDOleZbl9hER
Lp56vOSf8kE5aYSlZVkkrSM5tIO1xtZ2eBrrsPVuVG1lN7AWtym6qJJMOXmMI3cq
A95SDRusjjY4p5afsMDW4ytXWBtQtNvelf4eEF67kSgYRHR58Cy4grdDlmfzJ+PH
nohHqg08Mtt7tbfj1EUNtPsCMtVlATTse5IykARn37aVPbAQt/+xSeGHj6f7wpCC
HofjVzESHjX8bzitwaHE5eHqWmKK/PGiyEUX7ffvXEuJIyMqPnbWfJHzhAozyrh7
a21yGVAUaKFu1CpVszbB/SPugbHG4I0wd5zzMGzuYaukDH3hbbFo7jhF4UvFR+UB
+cWemuipJ7kvuxK9fbWyDkZOBLeNC472hV+h6XzqzxQnDYCZSAnMWNVG24X9uvKB
vmD4XiMtCjvULBJaZ0P94zCimV0VgDWXqlZUoLixGxNgiDloD7EuQt0/jWE7Epwp
6ZDziJxdgOVSwnV7isgaZtbAr6Nbt9uFrn9HjFfcefCP+8u1ypfajPDI7RDFzemX
SYCJDeZnvw7EagbO1bdmONJDLZzVrRGnE/NU/qzWsjJ0Yycj2bWcf/yYTlDmzLAG
2Yna4tf2W8E5T29Im6PYM0F8lePK8+wLno2gfFrDJMkKynzkmxXjlDBHhACHAbEQ
nJW2d/6djTsSjNjS8fVwPQl4DvrZn4HbShnN1+V4ttTwqhLmNtWNCC6i+tUuxuAz
esaAK+/SC9oNxnjvVP9nHPcjQ1Jyq5yuemBUUtC2rhT72rFNzIaQRamKL4pKPpZo
9pYVuylv6j5H0ShR7ocp5Bwqgjb6h8m7NfB9hSvkWfXdvJ3rjxA60TmQzFUtbRxR
KAsYY3mAySflogLqy0TSge+dVsAt5iE47OHCVWJe6XmgbZ5KRkYPDCjh5vuJWfV/
bALf66qY814TfLsrtbuNZSi6UcL2j+vUjFedeZCgenj7bK4qTFUauaiUVyYPf9ZJ
ur2EfsDqjUssiyWizvFVqX+dxXunfFvyJXYwI0RuzB2qYiViSQsmVo680vBeD9Ha
Y2tJRibfCVh2fZkKRgV3XJ0yKlNViw7f7CmlkkhOW4cH1TWLfx5fBL6zOokJGchQ
RczEmE4CDuQDWqIjKz1QWRYs0Td572xJtMcC81C9EsZHIc9p58ghIhD1AJoeluuR
4rVMRagHCtkj0Jorf9GoiQ40FaYbwhGjT/SP/SqN8lUpPmAorzhm6kqN29jODtGp
WUjWqKKaMHswgLY2pnzU1S3tlIcBoSCaCGhL5GGtTHXmrF3/CPAs2k6AQC8fxVPG
3znczuBItC4lN+ndzy1f9b9nV5iZyOh1d85PPolFduKyYLjWBa9jBZL3OK5qU/7W
YKP0G8SrLZLhoIBKLbUwDrVRkSW8fHDpKdmADGul5M9XSwg2lVIgvfrAJiqtivyz
Zfkfjtz66HLI9MwEp+U56kx7EP16DjJg05lb93X7WDbVIXCAiLlSc4iiWftMXOnS
y0CYOYXRS+REcg3RADhhDKWGlrGDb9kaKmzYYZAA+1jLWdJeleidPhPDKfpL/9h7
m2AID8brmIgQUup66QVWHpzIwOwDNiu6Q79+CkN0Bcks9R1dLE7ea2KFgdU1JnLE
r+BsJPoLHQDfcPX3mGBt22ICJXRsAya1/+k+PaY4lVXPOi+JeDJg5Xt6MWQqgyVn
5hvTce91QmZlowCRvJqGgjuXd+A7Hj0ekA6oWGtlOgIlc3VKqiHntG8fK5IZMfYf
2axOQ1ERrAy6MMke28//NL5y3vFeudVE4bm7Vt/+UyWfut/VlnfFAGxiU+gLnCC7
BmBKBSydg2lSgpnHxHWZM1NG3AH5iTD8dQLQrD55CRGuk1xaqtE9c3+oxequoFjO
tlQLu/5a2jfQsylpMlXyIjEYGqClI+MX+2l4rfOo/gRjfT3dHsteKV0yAfQQLAxA
uBbLNSCC9fhlH7kW4AJJBGfMZBtNVCu8BtXp/bxhdQqtP8skwpsu4rR2Lt0UOIi9
gaDKeF4EyYV95a5BzanYY2ldF3rK6FaoV6AbJyjytLG2vDbOP2s1Cp/cQGQdvrdv
JIIx9LLLehqfcFHd/7Vj/CtBBeAk7ozVgCallLd7P1GmNrnxSrgs42mNib7RjCSb
s1pbcoDF/UoFCw/YODawjlbtThMF9KT+ffLeDKjU2AR/pDPXFHJLDHefdhswXZZl
frpy2rnS99bYPZ9+6HkKfq8XiYmA3nELUgx7YuMa934ISjdxOxQ3FyDqfGbrzoyu
TuABmp06b4Y5Iz3sWjma6mXEEdv8ehgb+de0uqVHxP7EwufT5jt9Iiw8rFd06jow
PFe4dBsKQ4HTN3KlBcp9HLu/q0O1JUVgH8jeEaojoaVbxgFvrzXtZDvawb1sgLAj
vACnSwJ+RCkpA6hlFLLM5yT8qtRoZV4U09qv7DBgV/c1FzaO1qIF3jXjdy6iioeI
cAPtLwVWxLoyEWtfFvi2LWn+x5v+RZQ6QDbFXg1PtXiBbT+vhfRzjknoUqyBShi8
aABFw5lMbOdA/42Jy4+LLUUtuvLyM4xki/LFyX7CvaMEsaEHUqVXnN0UDKQB7Dp0
7N5SRsRrvDwt/QFopJMa8cUrb44mCWIkIv0SlotCOemsaeQ2HPImQcQVBmhREcYc
f7jGmY4Q7ny1d1Cu7uh2wkNlGss5BsUp2LVOgmlInktOlTEPKdfzCjcHc5o9Vyyo
ik884eD0jSoS6pQ0ll2ogL2IHUItfge2SwbT4eUYKP3eZiQP0fOcs+Lh8uqAkhAo
HKmAk/MnisiPHlSNu0GCy3aa6NIZj+/F0RpvZzfvkrXJ9JJq9SVogy89nXNFW8E8
enjeY4TBAfxa4mgcrmAlhP3XtA+bcwxv5APkDW+MB2JWSjBUUAm++L5sJHdNOpKw
+q9FSucFvEDXVmZX4p0llsD4YVcquYMCltoEStWncqVBzXChDGxKLtk2Nl/aNvDU
BHoqHS1jBBlzooydt9NpEhmCWIPiro/ITYdzJufwywoKU0GyMaUirTbLQFVcZ0bw
4LUmAf/61jhWRtTy1SvHmvTZr0BiCQF3NXPlVkmgD/6ZAFYhjsv0q23vSuXwDcMK
6Q2Dlpsed5TY+6UERA9j2C8HW7UPfSOYQy+jDFX1RFwCk0qIvpyVOtUTDo6sgyEh
nW/GgwEMkudcfwTOwiYVtPZ/+0BOMxRCZzC6WfYY3arPK3vPAG6zIGyB+q8uH4Xy
WL2oK/qldzyquyPQwgJCVDq4AST8yXaKoG6YBvpgzeBGRcNvVGUxM+pWm32DKTPd
rqttqHKExHDFsmmcjG5gwcukjwyfMT9uenrdt8sfcuAZ5hcrlnUMPk9otDW1W0eY
MWIZpdSvruKRIT+hNVnpLKkF/Mupht2yI8YKaMIfdAoWIOaBcVqvz47uQwguw4Px
wIEK496h9J5ThId2O5gF26pQrTYoAQshm39IQBDDRZUkmoSy/7EJWowxyu1O/muL
X9WOhjoqjpJK+GtHzeawuQ5vrvD9DjW8zDE9f9KTr1/4+fxoCqHEbCs5PxKt+Uy3
ci1WVROaP5GKXGmyL/zCzMkRwW3PY65C19243jXB4nSaGhwhzsi0ffX2dHfQtRvW
OfWzGjV7JOeMM3J2OeB65mWZ5dnz/Zbmz+PnEWfunojeS+dhxLMtPIMINVaNc8iN
O/JJOh3XPEmUgt2aTgRGXVqKUol/8RbPQmRIr0bYC/jjE8KBOdiIwQ22gIPx5fh0
cwL/1jqS/F1Qh0b+Un2PkOS7CarVaVVRG7uiuWtKHjE73q3vies344MeWmbms/Ig
6jnlD3mQKEUzONYF7Hn0x2nKPzcSwfPyWvnGRTEnUxZHklwiAtPe6JERbvecOB3z
6XxWjg/jooi9a3FfXSBgp3iaSq8DbZwChrt2vG7lkoXhUFCMKyIPNvAe+KdvJPxP
o/Myp4n3eGWBww+NDyQyO7JttjWZhnDCGyGNC1vNAxkZoInAh05kLc15F4ftYhQD
eiHM+P0pLOEUrRL3YuSxvlcPn//uxbXs18QdHb8c3VylMLfQVr4QyIswnktk3S3C
IkbvQ1V2iv3WWpbIxht5Xu/rH71Wj0EbKXnwrZ5sUnO8TmeWgFau49unL7a8f2vu
5oc7RImvDaoZ+T2q+lPjlmbvPiJtU+HxAk1QYWKKG936bw6tUqk6JmdI1gMvTFt5
rNtP4gOXXAUs3zqJUC9TSFp2K0wCztbeiFFnU3NX3cBsI3dW16ZsCbtQTzywZB3L
6f7ULTvpvOAXB2GlJUJg8Mv4axlSW0T5QxqLf/7q7jHrVaQJNE2t4zxSLS+7HaAl
4Q0GpLbu6Xt1rEOkMSw9Ufvu9oMogg4eSGAbKGYP7VMfQk/NI1tKDJzTHsqSR6Iv
8pZcFRsM0KUIHNY+cc3aqEwzwQoeSFlgQjOpzaoUrQRLpDYukXN+hcjFnympQ6Jq
4gm941kSyr3Y3H56xw11ZRGQHqmLLkOtJQEVK7FZWU3VnKfndS0yqsgOh7Q8fPQh
vQyk4mzaJm+pJu2Wc/ns1bVlvWQ/ci6vTVfj7LQE6id8/ksQRAmDVQ2GRmjSFYov
ki+sfTFuebSTprUb8Cy8Piwsn1Ayj+EYXOoB17RXCl9V6yXwoHmoEI8c8mncqY8X
Ma3f/Z6ecIgTvqoemjVwgQpicydIG8tFbiBziWVLuchhbHini3rDq3ePVg2UfARz
2JE0IDe+dcGwmF6XYe0kQAz8+MwhUwbS7FHYosTrgGNFG0+MQaVcT82b3QZJhYpJ
5/weEve2oljtLgXxRPFFd8EPAHKxexnbhZYglk0Mk3bzEnUq2XfV0YKmdbS/PMEe
GsfkWnMLx1MaTrEL73+FKnDekMxi8YdYd+n2VngXNUhkmGVAmQuIBZLjYWHItg/0
5V4cKPc2xfXpWscq9clh5mkedkBgYJU1OOJqaq6Vb06TiHXlTIRMu8ay6IPlJjqr
X5h+CR6KhL21QnRqU+/RO+rdLBHsZgUJGtcpijL8VF3Tj0uozH+9yUPwkaILwbJy
6cnexXSGWSCILspj8hvZ22Tp0sG5naRG1uvSLtEsHdhWS1U7NR67SWersmhBhS3Z
rj2cnVxx4B3fd/j95f+2HfsTFWf3HYR4ayEr9MgS4NnQzvFyQ7iOEphm/dwfQF8w
Hue9AxMQhObCYsCczSJYqKXYunWmRNUejTHGo1/dmt4c+1/mPfm5BKsvumtSwwW7
00IMvoPrFv8KZgEtTb6K5tOBHfayW4bxMkDBsWUmMc6S0/OMLbH9JJfiFDBYWllf
VlrUZ4O/uOTTfwEGwGnuLkYZEGlIeWG5ZyvE5OhGZvom+h+aNVReQD/VKJkRUyZy
/1yt6ebe+DFI6o3mW2Vj/6OQUKByi8pMVpdv3EqK23yPgHwNsieFfP3Tk0Z27UVM
Libp8WZwCSyir45HudYw2DoLMozvt6p0EJ0+2gVT4Gssdcntm7zb250hOR9BRH75
68jijAPaVpxWRnZIPlNjq56zXT9xSn2ZeSSM3kBlCawMut2ViE0VAWd/lIxOIUHW
I9p26UwDzpUHKJooRn9+TPGMm27N30TwWfjaWps4JsEgyxhlXa4IgFCGzW1sF1O6
oYJ2bEmxFhN6GjSg3VotWrtC4FQDJ0QMa27xmvL8Bs8PPaE0Ojvj24YTgekxQEmQ
VpBTT/bOyTESTRzCIb/rIqfJKvFaHWbp6YpofJQ3Y0g+8XU/XLGwHo8xGeLYHT0a
+ADoXf8TwclL4PLeoOCOA+4t+ljAfqylIR3/qoeaSgm2i79bVVX/SwKPHyb0wkzT
ssHJgYaoaeD0WvJC6Wbwic3p++CzQnVtQsJnO7wX46Ql6MBb1txVkal09GYcOOH3
2TKWdgoVfZJ1+Sb8IXA90PAfxfKu/xilkw8EMWfIIw3mM6IAT6EqdcrVBFr34SAb
TXBCUeT9LyO0q+m804H+24qoQuL4LbBTZyJBoRW/5k4pHfgSM6sTlXMdlF10WSZc
O0+mUCNreXrsvvpf7aAJi+XRxRFmT+x1G6FQGpRQmFTWC6N/kqAj8iVIGA436dBV
q4Vtl2tKrqgXZIyAXswrN+a5/zF0WyXlZ8SYjgspzC0c+RqvQRYmedKbP5Oz8iRD
qSu9bLzbkFy0FJYrrj9RjQo8xB/U0AnhqLKbdqDkTFxkrou4tuNnTqeZvTS2SkBZ
7F90ohEjeSNiG4ezdiRgaFt4kDPCfcZLoxuNK0DI3T9i+jYha4pg+jIHrvt77RNZ
NQC41VNq+LdxKp+0v0Ydq546xABiRYDcuYdtF2w5YLI=
`protect END_PROTECTED
