`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8EuIuWmNJ0q0mAuF/E6Hrd8oIMThNMbDrPwIq7/4gmQh3Jk4clGfpdZlYpQ23obt
uJ4Dcmu1dJ/g0KfmRPd/CKbWqY0mYINdi7PtkFO6Bq3a8c9iLoWu/zDVcXACYAM6
2qbhcydqPtXNxIcfdnGnVcKyTUc7VkNWS9izEcMpxDiac74xvHsKf8wAbdnfZt+u
oDRyeckWD91c8ZG3MzEefYdLTlJT0RUm4elgUEoY6//9ItX+DHkAq5EAK8MLu/oa
9kXXKnSdxBiH/CdiDKHN5E4bhmG/hJY98Gl4dR8YioOXVCCXXDXUksSlNpZhadRN
yoZ/y6m/4hxbjWchjyztAaaKDW1VfYpFKIKdjPKAaf4QE20btgctjU78AtNnf/fj
XiaJ0yUOxsEPHfZJLGnhNjmFwOlHeZjt4ids4/gH88hgDi2VEBkZLpjx3ahdGQCc
NgvUquLygpEyR2jPz/fZ8NcmVDDsP8XNCPwZvW3Isgti7uS9nc1LmsnEsUZ9srBO
GyjwgYBDy2mDX32OBvF149eFJ5g3zHf3AC2zjzWBNwCkDrHhVQz1xPy3jUKvCJZu
oFZ65yo5edVSZe+6LcWzR26rOVZ9KsmVZzGAspnYLrkRapGGGKitYkJ23XZZiCkI
lu5CKEn0ZYZ6O2E7PjVa5sEYKdaKuHJhxb0k1dBQw1ORmyns6qp8FkXewX8ueFDk
QZMRoHwq/YScSkmo4Y7ddyE/0VMPNQ5KJs+Jskjq3/KBtPwMeHD/Uad+zgu0MYpi
tD5xkowijiBPs9faxTFrDKWwi/vV1syI6igAh8K5MXexS8C2xohi7vNgjW8wfAs2
zJcMCs907ZbLlejPaMQZ9Z94fYZSIJjZJzlIAkgcqQJgi27I4kkNL0pOOqVKyNF2
vIyssAVEJK7Ol8titx3BdGjpI65L1+/5gnMmVTPPb6FLVdrIfaPpZ7QO3u6a581y
D0JQu3kCx+2yppLf4ieOoEJOyo18sWxDL+6WY/O1PaLxNN9Axm75DAYMXAGDg22S
yJjfGpcPOum2NLA5KcJmQtc0zJwZ8jSwKf0TzsJ7OUclXc9O0nl8FV+kvfKbyDiz
Vx2PrI5Th8PdrGF/xPcbMP7/+eRLf3hGyfsqoLUub7gODni0NYtT+yIT0HOgIex6
uQaU+EQEMQhrhpZf4GTavn1Ni/DQN+jz4N2uVPU3U5XozNCzUGZP3YdBEecIwJyU
rozWnzVFhZz5llXsAE/B+YG3KpPp/d4FLuW8+ELXw/d4xD/IZHo0Bh5qf6brUxmo
KXz1bGZsTzHZW/bvfbdEjaM9kabQOozkPlZs2xXiCwkq6eAYMeGjkX7CS1+4u0q9
HL8grecmRyWElAE6W/ZWJNhblP9t0bkZw93eQr1xdElgPbQJVQnVvCiD/gU0rAPt
yF/UuUz/cxHVBU0P2CU7LlnGZEv3EuiE4np5f/6eRHB75z23rsuM4veY5xUgU5OY
UMqoufu4Y8dYYw70AfZ7sw6b8NHXIOK+F2AUJVAMujB90rr31ssNcPXtQn0rSbQL
iojy6bl1Jg3OrtaduTvLkikKTD1sBJpaANWhKW0iANtA8PUMK1LHkcjjif6YO9tQ
RfcrP3jZcgTIekOWHJCj4pAzvZCixZBLUsUvAmU3g0okAovamjLj+7ae79cEPEtF
URaskSOmM/m8UgGy5iYdNevuBODIKc4dYaxEhUZbfNHdSGe6auTNPHR+mOK2BeTQ
4ebCPUGtMoZGm3aNEZJE/cekjDaF9NFU0VTPbs0U2ibmTln3MTm0UTS+HYW3ua7D
EBFpikZksQY/bCzXxX33+evP1brqSjlVNmgfWWcDgUHnlOl45Te1Hc9YgGmKoqP4
T7M754AFzmxby8OAt/ZL2Th9T4bRRQN4magfV6kLpuErGa+YvnnFl1e9dMJ8r1Xz
Z2yoINii4CfEyrkXCCxntO5tLBwOZjNLAeQ7dbh6LzzB6jMgiC/X9mNq0e7aQ30r
28wELUVauq+51f48w2UPo/nkbGECSTqX/YumNclJhhd3FY11PlHXAUhoIizPSgH8
ixV/VQ39dzwow5a9Eiax7iQfUVTkwIfgApu58qNF5LnJqYwHfducIGF5LSgbiStn
IQdaGd9wAUZ8tp/8EYr3Op7fgbjNE0N7iQsUUKURA8ZKhxStMYqQaJIOAz2uCszQ
xo5xgd/qW6YCZBX7NBttGRTGuNf+n8zQ3Law16fv4QHtMyfo6sWXOnjUlBrROzeD
BPM93zR1H6Pef6P+fbgbKnMRuwSa5e3N3bpqiVUNxiCZUnPb0i6O1gE8kVmIa9/6
Iw8zdUvh/qt5WwavO2Kmc+7Fa4L9oe013pHIn+crqTh/ZPHy3YDZfpxef98wwNbi
pxYanliavQG5unnzUkDuijju46YCqc5T3MFTJvac5Tyh/Z/a1sUtnKBdH1JwlAG2
e1LlL4wwy5Y43rccOXcwWUQ7WjIjiyMfdDImD5BtVjXb7HgcojH93PRIJ3slk2DL
XACqJ3fubvTMmNvHgEAMb9bbWOZk8aNEzd1um/LNSB8/1cu9ZSj1eOoiQqM544K/
cF8YQjGFQBuNe+KHLmL4DjVgJAhskny5bsHQQfw4bH5W2I2oxZU4VgIwCE/Dp37V
Pv0ih7LnjUhA+LvRXAiC+IbyCLY+B4yRkC/roO+HAEWfKGKsZnCI9d1UoB4Oh/aw
BVVS2XJ5a5yIgI8sXbUSA7RY43GWWhzXKkc9PF7LJBeXtrK1R3TM57ro4MWBWrqt
3yor67etp/3h7U8H1kZGSSOYPUYPVjNZFTkCu/Q2v02FQZNj4HbZFbsuu0d/7ovd
vjLUjltO2Lvf3mVBNFUbLZa2rFVWQc8fMztfrhJxxhQSdwOhj6cTrCkbZlqAC7QM
RIlohSCpiawP9zeVSIL/mlYC4QToaaPMf1rUD8GwK77uGwUgJ0Jobpld7xhffPrh
boRr0l2jDqTp7ZpkRrQlKfSBOv6qK4nztbdSzWaWX4nwbBdsSm7MLsRK6rv4NF9F
8CF7vrvz7YK4D+lGzuorlWNC6drLkQW6CSzyt3tgFP1OBlgctIhwB9ruUGCkrtja
3OrXOC2YmnOshzZylPZMue6BxywHSoAid5YCIImv6vcN0RXNFIbSp/Z8GMuq5rUE
mmdZlYDgH47Y3Ds1EQD9jAuSmvUI1F6zK848bMZj4QvYxl9Txz1PumQOMm/Y0gqb
Bi3+bKIW0+KizL17jV3bEUxH5V6BIf2bl0bOcY6lB1y2RukAYvyNWHbr8g8eBp0D
DcwD8y4D0B9rFvZ4l1RCYgbPjfPwHQnUNLnYL025H9uXDED8UQHJlTOyGBvpu2l3
pPsui1jfSN5VrWd2SEgVqMXwR2sLCUu8G7EtOjTjzoONWi8tMKY/iPAFbaBg8ssV
PuVWI3I3GlSTrE+9XOBIowqmLKc+IQD81oyAEBFpnQDS9lNgHrIxUS/i10eLC85+
NqpKkn4jVi3xFQY7UTuIEGix8F607T0ElS1fROkVc2K40g3x+nZF/yzQNmg3x7f9
y5sZVQ/3ZbTGVKuFpGebHYpCGFLwjNMiUsv97LchCOWwOYlc9rjEjV0xspjn7Wzt
Hznj4tUVQgLzJbDDdHVEq3kVKciSw4ui8o3DSmSE9hAz8S/ec54Y46sk0Y+7t62T
Qv3O2Y2N2ROAXSgvQ7tJXBh69319LR84IYQQnCu6XhqwBfC3q0FTbNNDKKci663q
J+qxFMqIF1KRR5viqn1/VOFb29VgS2v+Ih00u1yUY/BfOsYWgEtJmYS1acQh/giE
na1KWnS8CqwJ09nsaYYiA4yJhljyDoteIsdiiHxBL+3b13DPU2BDP4xBvYqEyibL
6Gjn/b4gyUcp4Btu6/ExeXvfcgIZUDZ0aXjwfERV3irXiGPqXrC7kZLrJlgTqnQ6
pELgw2tBIOTc0quZSSbUwo3rtRlVzZ+TfK9wnSkn7xLTWsNtv2JV+WG31ITU34BC
s+mTO/jNh5Hxmp4VP8ghyPHKbmWiT+aauG4E/UWkscyyNCbRZaiNuQK9oW0Ujdr1
s03F+miyvnG7/LCfTZyrIg==
`protect END_PROTECTED
