`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mvhT4BRQQSn0ZgHy9sG88Sd9x0boSomoEUTjS60pGOMi7rx74akArm3oU1GVtXL2
4oq719N/AsHgphouevuWl2l/scwbB9ldDXakBZimVkf2axKnZY8XQ5/g10XzC8LV
ATmEYct2zb/QYCf1/8NbXT5DcJOqVXT7XIks7ELqUAoJKyFPmVNcGGRU1tv7p7TM
6/O/7ykqZTjOMFN1MCAUnfsJJjHVWT7JHKaSU4xccRdITrVQ2hOsYxOD2AdOtFQX
J2i62UcZoQquDJje1HEbsvgOykyHSEnJEFO7xJWJ0Avm2GPp5P7WDXgLGWVYZVR2
WlTh937cq53MQTKux680ifj3RK1h9JVZG86AFU6s74MRpHCn70hvS/zMklAzEVYQ
6pxND1bF3+0c3QhmAvBvM9E4f+LPNT++jEzOE4G2+Fsr7b9gHXeCQuhjwz9wVDGH
hOyUhtu6lT4JahISuD4jFpiO1hA9EwI5eO7klyN00a8whqOEEKFPJZohp+UkusG3
I3NZRImxjgEX7TBYgjpMC/aNyoSqxShMAPrMDgGbQHrHSj4GNoOtuTs4oysCanUK
R/LRibPAP3juz9LDZAOMLVfMfCBJnPSeUn98WjRpnuEhsU8pOW939xYucl8kSrNv
9kHo7RiD3ArBKRo+/fR60Lcd7jO4Ymr1DznJ3iYFBjhZ/OQy6I5w8qOFxpMQtX2A
Vujybsx3TfBljR1SXkF4rRnrGGRv11+5dOiNlOuo2JmF8JFUlVy8kvBsVFCxgu+q
Py4/gyRZHMCISJLs5GiQJIoFvJGePiLdz4/7Jf4yHoWJqATRM+BK9L7XbEcwXokn
uUXdcgSYZIF4fSRtstpQEfomcXtTgeWvF1BUqgRHwpHXy8VD5wNkRH09DQdSgXA3
QQhjk1aT8rWPVHE18S3DrRwM75RyrUUj64+mx4jwkcMy/6XuGzRC2itb22lWzquL
19iTWd6DderpiuQThXxC92w7oy3KBtPEsj/7Rja2OiAwgXXfcfH/Qiw+CvGPJJqk
ZXTOj/zWOCokXkHLGTnLaw==
`protect END_PROTECTED
