`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eHqC5/lGUvKVfoIEGO/vPjf6UDPZDnKtCDEH9pJSR9TRJVcIVtfynujC8QJ/SeNb
6JN7iowozRYSNI3/5WX5aMFjcKEcNjTj07PYrgbPAoOMIDKZU4CFDMWLKK6AM/Af
UmqHGq7NO3FNJ4dneuXM2y1oJrgqZTe6jn8lVBNj/7VOqfK+SKnuk7WpJX31t4PK
1YbtRg1ysphOVA4Ik6WiWQulaMDheFrnYV1JdkA5A0G/A2Auaw9SjG1L1U8zfX3o
bSMV60yEX0IqZDfqUK0Di1JiJAZ+FqCV2pI1/lPtoUsAs4t/PDApI8fUXYEj9x9p
zmK8RMkz2XNU1QWX3FDffyXEk07ZNrzW/fWXKedJIcZegQjPngVW+46ifUiZJvQE
sMcjigeQPujsrAYOtMpTWaGC8ZfySjb14+RWTK5YoHDgEjo7SzFknDO6aTsee8Dd
OT/PIOdDRivk7YwV8vOJ0/Xylo7Q5KuCXUlrRBZr11n8KCqpL9PN5nCmVJOHuR0z
/kjVGixJRFI9jOwx8auNzW9HpT3vKQsteB1N+zjXdOVm/OXtFuRiKH0N+RFI6mhG
IuIYwWEvrk4XjqUwgDOuldJl0te1njR3GiC2nt4ACZWQDPtV6ca91Q0YkBNWIUTd
csFtPlhvgJVnHYda2DN4WWuYHIdBM2w3HQNrjZC9RMhVsHZPaYeWBOg/zBn7uGaM
Fu4OkZSBNTSCQF45fK+MLQ52ziGI5zqjIjmfGJ1th58800Xq2r10JYZHdY+B8aFN
VsLm4ohoFjrF1nrkCt5fSks+yvJZsoeTUhbtGk1sOEjg7iRy8kykpIciHaOsEZ+l
ul/jXb8KiQfSPX9Q4k4mgyNcIbuifwJCqmtcu1H1EylbUrlu41V6quXHjWzuaicl
aIqVjRTKR+GWjC0BPQokmQ7q13TeZM/gHXqaZnvU5PM/Y8wAOWRnc8QDDF/QXWt2
9WgicFvkWBHy3Dso45OgwfazMPDdssLSlrZL1Qx5HCabQ7byxoBrbtXhzdUh7e+Y
rJQWJ5vDRwG8fKDvBUAoVAJvXXz1E97i8BVJ/o18/o0ISiXnqbmYvYCkecThyM2+
VbHxWllr+ahyO9dL+ReT+9Z4OYjTkUIwZpf6MIO1VP45OHXhtT8+yU91+B3rnWND
c+xgKi75NMy6e5W9/2YJuICRXvFPefma4REtibsCW+ybmYi/bEth2vUO2uTNjHut
qz7u9rrsnlXRhSKqZbiMLUc4qF51HMbQ1SO32PzaZZF+BcNQLdkBVpSQHykA7Hf7
i7Lr/YdEt4SlSUeyzc/OxJdIksDBTsCfPEbuj8fHdPzITOkBc+z4d6kuASdcIOuI
JY8AMhdNCUg74Mwp8P1uq07kkmWsq83wxGcRy3TF6L9mjuOApCJ+vB7TjpKjoNnz
fdfUeciLxDq7JGeM8lW/EKZAp20TELyLKxSasGimCvanSgiqiTr4gt9FIeEHSu1T
mlmXQTSeD2PZkkmqcepvootbQHwju2MDt1htX11y1eIKhg/2FkUZO/ZMMsAmlNkS
ff5Xr2EB7eUpATKbGlviBH/PKlX2QfftMDynUHIkpwLKyAAFN21Y6oxJ9zSdK/LZ
697GtHD6VCBj+tW+yXmHlRUqYGC4CfxY7YfukmMZDYEwZfu3ORx7zWuotFH1HYRE
qobVqWDrcoWyvOqDKnUiLCuxXlVOWe5C0JP6YAnPD+utdYxoFOFv+Z/w2FbCjcJh
UfoTrvXw8FTfixS+YzcJFt2ahGZ8wzhRVE6P1f1z005VtHcm50sgeZ7PWL6LPe41
NmPsmRxg3TfPKPyPpbFb105CdJ59CxoAiMZHqWxe5S2VDFe6hV2SefxjkP4g2/3y
wsnW1bLsbQWiI7ztSgqv8KXz9J9iFJmZgHCqfgeh7RdM0yUnEgJHlyRXRWKXmdNh
QOF9CqlgiZ7EsPJ13sP4JUya0QEeOt2jVYOvCpOZn4qoMAexaUN0JyhzXZTg1EzA
zMiOcvh54vydunmGRXzJPsfPeooqnc6PoKgEiOJj61O1iwrMgbC1av4Y3v/QZHxy
UibJjh2U8wjDXGdoAoqxLCR55rExFIO8lEs/SjSSI4jLZnTY49q0lcAS6CZsstwN
kqwaHukXCy3s70+1/aaxKLAdFNyQc3ko31xm+2AEfU3Z283QHaY/QoX5KYUvA8BL
B+shNFwl2LGVahn1gtTEk6PtVTS/aawaB6LtangheGxHPn4hQUJO41+KN2dl/CWu
N4ZSc4RVHE8UjJ68fddNfx73oOIV08w/Used1P7X/VSDXgsbUC3o7wpASJJopkUj
EFOSZqyUSbME9969MtFlp99FHI7KNYcLOpR7kqIEuWROj2u6EqQvs0ffuO4e0VDh
0pBrZGD/l8uYhhdFwdXLNLlRE9zPnycZ8VBJrPHUWv2/w4qQq178/Ml0KhGyyvf5
SpEzOTbHNW1qzFvPyf8/8fzcyp0M5mX3qio1G0qu32NmSMPX/P0+LoWipTrDjMAk
tps+OIHdEQUaBNNrlbIpYf+pShc5ieuTgI2OzJYD/NBwqnEngowF+8soNMAvhQHk
qez649O5RJumf/O59EJnRXpmhFwBmlwXXD5rYhoaEScIteCJ6aVGQmGeW8JRMo4M
3QUk3gjINBaTHR38uxZO39ztehVHr46QEZ+bxvWnNij59CUv5ySkpD5k+NHNCo2V
dAria64IYgI8UY2nfZLoG0jo2hONAQcSpDeu8IYDnM7YBMCehOGFD26ArBBL+Bus
hJVJIENDSn/+IF2YokEuX3QE6dGRBD2VqprE0gvPfvukDEEh30fYCMsEKNXaqsNw
m9/XOzToJcbQqai/nGa7rrnlx7O+3A1SXaFsOOCUiX0=
`protect END_PROTECTED
