`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OUYShp2H/41WRZZuLyj4qHiUYFoMzzHnHokoTdolF1zyhGWscTqrGtBjrdX+nI7l
DCKMHH5N/nLLvm/jtkqYqqnj3NK/UmO/gxGwfmzGJxQ2IZwZL45Q4sns2A02Om7T
eOTs2Lhs56LJ0j+RTfZa4bVCh8z+Jfvopz/wB8AQ7HEoEZUB58u4at+w/k/gSIAY
iefo2kg9OEQCoRg38kBC8rO8+AeS2fw2YsUmsmGeWRZ7a0zYyWwExLOpgzcIYX1r
g49EQnjRlSSA4Q6Nve9Q0OYuvGXLk48KVVe9B7FEk56wH7Gry0hBfhWuedQ7KPCF
+0R1eX82RmzlMFJywo2DG9KRbePAIjW8Aag/4n2j2BS8zcL0u2/BmZrS5k0FR26b
KZUHTWu6Uxl29xuPqf0qssZyCt/5D7MdpxznCjC6q0POUbUvcY/lzR+Lx7J0b+D4
CeFkU0H9OVjsRDkW5u5iIdSDhSbkxSCTzD3mRNRwQT7ntXmaCykWCuR/2/E05Ciy
uFybUqC/TDx8eGTVmAyIjqxoUS6LMrXq5kJW6qxh1TCBvOckuN10NmSasZUMbojf
5Y/xCThrtwYU/eA1GpKCFGDN6JF8ML2WFcjC6hxgovfnprUFRXSyhwfxG2HV3MU6
+zdQ3iaU2YA2os1fQj+aR8wkCdwXsAvQL3Oxr+KPuggVg3gQtxRZcuCZwQIEgPzR
HCvlY4wC9wBS/hiJIUG8TQhEeGQMLHn2kpsL1pCN1Zb68ASdm+o/L/LzeOXMNDqS
oxtUcMBdePPc56Z0osw3hCUVubH01yf5+4s5jGbDEG42RWkYHmU1N6flIjwKr1dO
Ld5zgpw9lT9wvkMngMraTLZHymxQp6yXGadAZzQpjWzLifOeLFIUOeVw1IE1NWrq
3d3Nc0gYLzHoucds80wjlXn94CwxlDZ7HoE8SXM2ZqL/E6hkfa1W/wosrG6Sdt3W
sURY8+IxX0FikNRPrjeIV/jdxZuyoMQqY1QZI394RiqQrejLagNb2aY1V7L6rA/K
iSgV2ZQDhbYhjDkqncrXARZ3HSzs+GOR8N8mlQaVu2s=
`protect END_PROTECTED
