`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iYMMcsStnRpLIQoXmIkLPadA4fiT1dXKKJRiJcufrHnaIhDg+QCqyFLkySCtU0cJ
qrf9+9nLlK//qVq5643Uv5QIomAUsLJmTsHKsK8bg2V/DyC5/vn8dVAOGvtV89Ve
vZdfKAplf/+eKN6dn94HaxKUq+YygpWTdksMBfZD9aFDC9sUfvxoFMVjFHKo6zEK
JIohkrHtXdU8ejBd3/jZ+MZbzFlWhZ49dvdF53uXZe7eftCyc3TRj+QdU9NbpS11
u1D3wZaYOiFFsfB7PcNrXN7Qdiu/cJNf/FgLZom9ZI3A3wG+0bzCRCKe6RuNKocl
cKGqx06VmsIy8hCw3wa907QHmUqZiaFIZJ8XtH5INnvzfXkhRoRz6BygUr7pFM9c
VL9YVLBaC976MYLrS5wdcFmL1U3eEwhk1TffjdChsKhH1ZPC9o2nu5UkhHF5dber
jfgTEIvrqXrTg2It+s5TAAgnYPc2y7fVQ+pEmtpOhZSPRdBjSsqbY57PRGwPR3vG
wpnxLmGEEkfOnpCLhZZlpgOgqwMKymEGy6yR3TNKSh7RbfBMYhzTYtKbxoxu3Um+
YPq+DeZH11C1tqNrK7acNnYbHQ0F/fTzbPFHKmas2w1p+sQMIdXJvp/5AXg022Ux
hF1K97JuY79plcK1CxqfXvvW0974axcPcO+m2Du6Airv09T4QTV5yoWTWc5pc6o6
RWeFvhG59eYmPheo3sl+xtDQ3oEa1n/aPs0vzfwZH2MjFfxtxRWeqGc+mjV6Skvp
9XLl0xCi8YdyBg9IC2Z4chAr/awewybNGwOYkT5FTjRyoOPTiEKEWJwtlwSHHjW1
7f60Gp6/nm2wM4umLRpwNuOSjc4UbKRh5AKZJdOgpbhn5gCwqDMhT6o2Y9LA7HhD
mqEb7lfhJZTOcb10oW09ugGzIIoTzz2zpPNTJtgelgiohOD5RGpYGsMMWVtDWWrY
5VAeegavxMm/QooHGpclKlA2sG2CEuQNHQJhQ9c2F0pbcK+i+pwcnUzuq6uIj6TF
wHni/HuugAH5ExpfHSkwEFVYl8fkgfOXw/2RgFEUhg28YlPFWqG/Fg4uywJe/PcJ
8aCstKb98MxeSBmWtVG415nNguhLvYniAHcWkaKLmGFdJqY3OuBT7LcoYu671135
0XsXg5W47gr5l//puG7P2EiAG9k5I5R/MgLYmpLxyZQ6QZUYUp9fn0tpZlFaFZrq
n0TSUwzXP4ycN41U5XTydgiBcICszs4swTMNbl5V4olDGgNWwR9a09G/R3G/cG62
m5p85c5G9lWDhOcR+UtOAjmX02l+w2ZplWJtjKoBtQKicY6crEoMi8n/85FyDyxi
uDV05/Rrt7aPnrXvdyo3V4OjWENClnMvO+zaFU3hSA+oaKillgvM8UgS5kQXBIHr
wSFAUbwgg/NzMs0Xep6IQYbdTF+ZyqBewzDz3HAojjRc9AouhilJSlQ0wCWnhBdV
uREJaCmeSknF+Zofj5c21UVO6k/92V1JBORVjoH2beEHi8eI351GnGwR/CNP2DFa
Vfa0A9ucD7bGF9TvqGcp4jg+QlRUgaU/pikjWiFfDesYeqfuAfQcxnDHBY0TLAuU
0modE285MdO7RiaNMPjgjDZoxRaUB7s+8S3+HudpSg63dQQ7sbL6L3f9RdDry5/l
R0pT7FzMHapMu2WkMhVsP39ffg3e4U6jhAjDBlnIW40lgTSq6+QO8Ul3yYfRxc+j
WwRYT9Rg83xzNS0S7xtANhZBAbPjvaYhIPkEvo1FAvRVEcRnQ96Yl26VC8KABG41
hABZcJtajR3sCdIfnnwCJuVlGCooPFTm33KxPzzK+HvO8jSRA2eM/LU1V6Pwita8
K0g2CTUhMQ7/89UvLXpYVcj4WCCihnefGc7mhae47lzKxlVWq6hsCm6uPkt0mGXV
muSfxKFgSgr+cS+cqASGYz8B8N8zvohEtTM13h7bznbM+PGxRgfkEbQDTPxqOsvK
5ncj4bbIAYkj0Varp0jWiZ4QtaykilQJb4n7RhEWjAIzGZOKxnc0odvABXxpR5mN
x1x020UHbH7r9rAozTzFtfwV23Q6gxriacIRIBNmTebxtuN9I/h2ebbXE8MZbX0g
I5r7d3dX3D+FR3CKM2W01f319MwO2EUTsbfJtauvpyNDhUXNMNoCODXvbwEvu4ws
lc8q6ZBm8/Rc5DTiJ4VHA13HjnDhawxjHgn+1KJRQ1aGRFMuLWb4BEZV7nbTTtIq
X9GDyXJZbssJB3nYXpA6q+fb0FG8C/QMURq4xCah4ncd703r6tWJaFSyD6TnhuwJ
cWdWAj9VSntcLarboGawRsPslXHpPfJkqOfzhejrwH26YD31GvhxqJTtOy5V/4CM
CCIY11p/i4BI9ViWBtfFex/7yeD84lYK3BoOIZ9a9CQjGvPQRaXMo/KobS5TGVyp
1seDfJdC20twmkQvwuh1WGsd7I8F6oxoo/bK9iRt/LdkE66/PsJM7Bq73OSRaCn3
+jvNLgWdlllFTdO5AMevrGQZinLqHTfbe/2xO2XselQ=
`protect END_PROTECTED
