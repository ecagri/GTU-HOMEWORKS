`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PLPbhf5jEZpz+JViAQ+A/HcaEfrbVJpM0kzsRGqZrTc0P8hO5RDfigAxMbmJjEKt
g26boQLuG+fAFbVBGXN0ouV9m8XgLULalkRrnR8P+4nwOynMugF446wKVNl7CX9T
L4U/TzexMWw5z5er3Y1D/Rd+/9zyxMy5LEIxxyX5NO55GoK5ld1ioyChciqSOEKw
VlEPqG96pUP3wSxiKSdqC4KUv+++o5dZcPG78Rwndsg8VNcaZJW3I9E8LS3n9Cbb
NI3X1I41FXd83EFFSx5uW1t6BxMz0tbNpGcFnS1MpvyLltccCw86vvdsFNsZb9tf
2vizo8AR0dh93yHMitMfA9bQMWa6PGVgetUFM/rP2KLEZDoI6+vam1AODZZH7zFo
594yDmfkJfNBXymdbXX36BD11IuwXchz3x8RH7Ek6K+02paY/wM+w7cNBdWLEDJB
xqkaFG8jy0Tny7WVRt2l+2K4F+b9eIAOejSBkUOogP9QCJ5S2Bf61vPepjLWDLMr
AKP0rCpe5bL4fPOe8RpIH/YxOG8rSbJl3jszt++KD3uGPU4ew/SA7rJ0o4rP61Hd
w/cXasuHcyxvXRFyEsJSXuMC8GEw8NztUuAyuNNL22jCwccJ8CFZAyHZqYlU2HKj
0YWVcugGLPV/6U8I6JGZRE8afFfFTjr/3OB+FbczQIs97mizFx78SLd9bK8/Fc5e
cnJIVWC4mnVzJpxYE1lOFkcdgsV64GB0QqjGPeVmRtlnl2rrjfdMhCUCmLuetbz3
2Ovi2RNnhHulcGm27iALvCxNFiNLyJQ4+CoCj0BLET6Hfmv7ph3JkDEs744krnra
Gei3KfxvTouiUXVtj6KMncbJIBVwhom6yDqSDouB5K9NjqFqiUD4Oqpq0qDt2jtt
oSRh38UjvM/Nfaqs5dwh5PvX8A4gwDLvwJce9Pv5vpTAhfXZ/njV22OdquGFfDht
BITUtPrbO3b5x1CcdIzMc3Xa89cpxmDUGeIjXwnrA2YLBEyL64QBD0TsMQeVNX6F
6R/PClkgXmhH3cpmeoAdutpV7MXyvZRu2eLzFpeTItUchTn2k/9ttnxXd6FX7M9C
R89LpZCWnXjXqgRQdJnE6Rmvq7Z0cw57pOUMI/67mn59EVws1SHCSExuQE1Uf+pG
5vxB4gujyTbj8XJqNxkKPrKIj5dnh6n4/2vQxoebWxfAYz2xcYKCCXkwOBr8gR2H
HtbvkLCpkjKMeMg35+To4b4Szc0Dbu0kCm1q1acCEC2f5zg4v6lwxcgEScdZ+jDc
iB8gX7GpCpPtOTXs50lj8uDA5SzqGMl2/P/WNwTU9MU8zejvEAB5TxSVQ3BZNFku
vuwC31xPopVVnu+qIWuw8RIdzQ7vxR7g4avW+eADhfTS6H9G1NtPyGAYCYa1lFJZ
VjTwgUcOvhw0LCxtlsH1kXhR8zXXyTTYycLfSS7CKib/Ji7Yffnr+St+ZOIwoAVe
N8miLtyCt5kxvLwip65VfFG92g5ZvgxG/jI0DE++D4rzcCzF+nykCOZKbOEfKzlP
CegAeL3JqZRXYAr7eM4Ig5EpKMUKq0+65UgyKieNBtcUnTOJtf4JXxYaXfanGEoR
TrnxnzYkEP7iqc3iXERzuO2ndDqHwFlm5DHXDHk7MrVLyh1XykPhgSMiDNc7OVxW
maKdW0UpSymeS++wMn3+fa5Urypm1bx2CklCRSXs9MLboC7312tLvMmwHHjWtiM3
fYGRcPzwVEYLWYkBLmMRTjGFQwFoC5xxNX67NUjUZrscExY0v8lPZjnDGmY9JpTZ
8TcZO02yMxtsOn7U+Bm/8GDdJi9eCLqb/2qSXWt0pmlLGnaaOF2lO9lP8Rualf6Q
ST20QqSKKc50DyndtZrbGQne1Z4LPJFsLorEmr0eKnvvJDessenelcLKaWaDIhoh
2GCZjzisug420XrtDLntxuZ3QIP6y87S1TtAbj8W/ogrNEH4R6JovWolyj/aX1VZ
uD5NPW9kGc0af02bHPt4E76KUmbyIkH0pQCFSOfFvV2QbS+oCSTRuSu3ffV27hsQ
ipC0t9hhap+MYTHrMQZ8cUk6iW/Va/1KHF8btDlvb2m/o82oMt6A8Fe+LMCO2hMN
gUm3rraJuhxuqsq/RXGFdtlzfF7xOdScBqC1oyLDGFS8ApAsQzLz4FRnr995plaQ
3qNdiiTPJqfiqE3Khjcjpt7TgP6YVECcCtwIW3ttNLI3RLCDUA9AE3KDK5hozuo+
dDQFrkbzUhhjLgPSrvCey071cEX9rYP5yKdutNygz67LwYANZxsrRNjZy+QpgCsW
OFsjPG6Jv81zApdbFyRaT73xSpDOauE6ZJcdA6H6b5j/HpS9Yw8JpTbLcatAHOw8
NWTdnMMvyagmzr92zW0QrCmzlEGignsvCctNRIN8dp73SBS0ZndsxJS8c/GtuJEX
RL7QhG3OJ4JrE4C/zK4zhdmUGdVMt36fv3bIE7szVJuJzlCLzG94i4gYK4n0shBq
Cc7G34V4KuyHROzCPGXUDaI1WOEQh+4e8GkA3/JxACOj+jBgdfVeuqFcRG8+GHxn
DV9JdX4U4THBoQjIH6Spz1weS/cuWv3IcMOjN7ogUcHwPmI0H04UEwfes9jEC8fg
CTmbifbEN+Iat9aWUwW0BxyW9V0HxLbTG0mvDLK2pDOgu6Onx8b9lPk2x/3Rdsy+
FxskkAHGqpy3ua7lD6K/SOxEC8gu9GgUVDR9KM3mquBijw1g2j1aiITnKLNQm2c+
4diTcVCabiGttm9gIzwODGg659iJHmWa6h6WALUKLHPgDTSCUISqO8C0rVg/564r
RPuk8I1C8qJYp7K+NtEGybWbNQnHdCVxANp6C2Cg1iqy3fQ+kWrQTQ3qI1dv3gN1
3qFVlHPpVsqG3Y4hfWMqZ1MkGNSmR6VBqHE8kbKpuwPx55OFQUXETnJq/5gKnOYs
GmgHm9gAKz56Wdx+9w3groq4c+xAT7UHv2H7PMaLxVupSDypPhw9rKT+xvFYmgJk
Hwn0eXoiU7gt4uE82GveWus9i90+orVFBlLYYagK/X5Rs0/yc+msVN4F2+4lG3QU
GNJbeT5DU0Fbrgr6yYybvvkbWxhAtVT5mnZ7+bxIHrYPveRTMwjSYPb3+kQY1XdD
Q4daoeUtubE2gSEHf1V7kik35JLRsHc8Xsv5gYFKn8VsdkKSkifvoAiYDZl1nIgw
siDmgJZZ2XW93TDTiEHfLFLgeBzU1FBRvhqnRzn7L/+5FcBuxCFAN3X/PHdpYiaB
sstgYhjoE7KKioW96BC0KJoNhOeeuxQliBc762+IYnlQ4Ip5cPx4jpN771rG0Cpu
qKUzwhzwHSjnGCKRyY2/qAobFIQchkSYMpgiqmw8nCou20SvDIBtmdTYg7oMB68D
+CI4AqwT6L9I2cjw3bjN0kDj8Y07gmdCZfJ6Wqnny7HuGNqPKRsuOG6wfOSoLfkO
Z+m0OVCKxqhLU8Grp+fC8gTNhh+Vnius+qSzBbAbnko=
`protect END_PROTECTED
