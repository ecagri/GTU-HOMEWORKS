`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9l/5uf9whs7ovw177rktkHgQ4qJ96Msv7Y/44TjKLRfLgM9mNcSAT3XP6BGXme0D
XndkadvR30sZa+LcgtGCcmt8SAofh87b530qSVnH1cfsKka8H/cXc+YeX3MWRXv1
wlRe1koXITBXOj2UsWCWf/L9r8APgRBIRkRC/tFqi7zhETzQiZkjUKcTgwVvgBYo
CZZY7XpruIXJso+Hvn5ERNy7qNaHpZMh18fyr36SOVy3JDnHLzdG6W24N2ProqbV
6Fwk4Bugk+/+VArDjuooumExUFNys3shr7zBYoBdQ8C4Id0TzKoEbKtYQnmfdL6i
EaiiYX5r4jxuRWWAaBmRFP3htTOKrH94Ml/XLzujniE5HqaMpnXU1GGaU0wgCbaZ
/CfpO/Cb15cX5hJDO/ysCx0V2XkzGTvPWrcpltRmQopWeISppKyK+UtTNheZ994b
uoiPF6WVjicNPP3frGs2RIQIKzoBNnghfpuR5BaELnORePwBR5K0syO/gNirl0oM
iTK9kBOqKxOdHWjYjbcNQTTNQQE3pzcmSO/P8UhhYJ8OWU3vaTog2Kc9f/tMwEuy
795+jKcx5nbsLCATHv+0Fko6DV8hj9pGhLi/F79+DfGZrK6IdzMEploNDorUxsFh
DG00qni1QpeLJFhbQGjI6eS/vRryx+hFbY6vCr8uLtcG8Hp71/8azPe7uNEUathp
rU1yKihl6qsL+nvQ3GyhzQOKJNgJKVlt8FCE/QAlckCHgYz2W7BhPspIcKb+xePi
zfCDjRyX1QIgmazYKG7ohOzxYYaJCobOpOw5kpJbAwzOZ7C8QO5CBbEVH7CNe+A7
igUWDzA8xByd4x9EMqlBODZS17aOgrlE7K6Eo1svG6m8KA08k7m+ZH0MKrIv+VN4
rjIMWYwaPpUA348iWo0v+VjOOCW0J6DozbDzHbfIvSJgmWKcWG6NmC+bwsltgxyH
jtjc2TTb6aoVqXuNp224bQnojCxnzgb0PRQg6g+b7Fc2dRKzcCsXLdKQMN0l2IsF
co4ScI1ndhHL8tFCrwDV126KZMZAtNRwGrpWlNA9nXtzCkefAoJJjCCWSmgbCB+L
cUQqbs77KPZVfvKmuoObGez0gCuu60bWdxua+LZLHyk=
`protect END_PROTECTED
