`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ho2L4pc0oAbyTEmFnb7JPQBvkxFTaErfIDMEksO8DfTYdMe8bWXLleVtRhdrqwV9
PAoHUeKbrqk97DrluWHwNr9m2LElwqkvAi/ulubpKd1qzgsytwSWVa4mjLzu9PXc
cptfXUkOZVxgfzsUfNfzT1d6Q1l8+0cbX8sUZJTEW17v3mKkkLcjlV/Y7afgWnHq
GkjvD+nH9/Amr7rTXg6Axto8rA13BAyLIPlAYDvbBwR3pFAfbsf8M9DHD2SiHAEm
zLxlHsV5w0BxbTTPvV/q19UlqL6TaKiy9ZphTSI/28Af/Roe2458Jmj8P0qdwGLs
8r1aDvMZCfn26+r6qR8mmS7TROlL8GRyKffalPUhWsYOZBkByEgO272h9epOrwtM
JvZneFRL9pg85HFJNWxCpMWQObx7jgU76L+JsXltye4Dj00i61TdcE+oH5gQestS
hHIg7QyKRdDqwxLoEjTTxPlMRT3RyR/T2lqPIcCgWA8VapO3q/zf78pIyMMKFoVg
xJuMM7bZ8UDCx5OKmbK5x+8/p/oN1lkC77pqtGgWfhlu7N5Sb+9Ek4CAQf/Fca5e
dPVUGyZbBA9gRxafv6gaoK/JK3tQ8g/dDRscqFsP5t1/TNx1y9Tq1ZwiWLLrzoly
U3gb28Tl4XZCYbZQvmJXnUshLGLm9T86s+uRFLm5Z/BcaOqdtbD1cRTG/0axKAQ5
dpxD/62suDYb+BglC0OxfA6J+c1Kjqcoqo3w8EogtCh6YCDaVvhW5IdP5i6Uj+6W
paaqHUQPFpkf/4lDDvm9R5mbtLANVih4zUvsyCFoIu4/5P3BRBtW7FaJM7V16azk
JXtlpr3FeRprLTpie3o91rNrIQ7RxaNGGvX5DesC/xT+6qaR1uBm0W6siaD4pKik
iyQsyFsxrYysFwdXlL0GHQCHflTIBL1pBeBekk5XBxXUC+O1E7pHpmawPnco5Q+a
FPP/ovqW0WWDm0tjuAfd4rr38dr7Cj/3odNg1cJ0tGu7j56j/+zF93kbxuVUQGkn
2mZCo6JDdhYjhCSFdSvCTVr6tGAzJVxNasytXsrUCkDqFTLbBHG7b7mq17xqjzwD
TFbY6tMSvW4M2j/jY9ni+Gm3f1aRvsXf/3QHpMIH9XxfXLOS3aZ1dwC3Z8xbuCji
ibvCSOPQ6HhBgB4f8TDm+kZHgec1AND00698Z2V/2hHrMMsQkrg4C8H3MrN6K3Om
fnL/ppewceC3dWckK+AanI3gDi/E7BvValV751t1ixgU2Uk7wjgPCw5UeKE7xfHD
i1XSKbFfNYPLI8KoDWB1ojAg81+AIaK0bEpSl+6ZeVr9V4cVf3z5HE+nyIBJi3nx
t/N5UxFRz78MYgpb0crrp57aml2gsNdLXj1ZDUEodBk5Qb5WKGd0dqdNuBoIeakB
54GLV3DUPLD2tuXcBUxGnsTZaYa5Awapf2vDzGTvh2mjTZXUy7GzmxyyIM0jIWsA
`protect END_PROTECTED
