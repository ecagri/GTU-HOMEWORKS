`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SmwKLAGX5BYBxJNeXvEp8jBbt4wspGGZ8U2AX5v5tz14oaIGHaaEf8or5GUE4+09
N8p7qqpUI6Cj4PPxEpnuv8qf09wOziCtW1dH7sV1Fw+WbXNrAOaFlay8jLZC6dBU
IOP1HgTYRiEQ8/DxYHBAAhsy6cS71d8QnytIi7B50YiFaZlXDbLMUuCCQ9CLeGgm
pIrwMNilwFSPYHWbnHjfH5/+VuEpfa4rcJilJdXZVBWCoCs7+BM4R1whCFBjiTqG
UdxheycCiS+AzTrhKv5+xKTJfoaSyt3yNXFSSNq5wRqROErfNhu15HTL6nvqVYwG
ajvtO6cEpwq4w8NRRba43wvSYYM11aj9xHzX/X2Af/C2cwPuS0f5ctqu6Z3lOltP
1EYEQfuMSx27leZ3m8UFvOOhgZRmUDHGt6oMosTfWjWWlnZrRG2d1qTzwkvz+Ebn
OQNzE8KDalYTVlrLaxcV1Cc2CtM4ulfdeZFxqNqyLL4o+kkyhhe3UfcR0O0fcaYW
x4bIzzLMwdHsmptt/F8J8NUfdw5aRalXhnUiEI8pb71O9l2vSDVL0u9SKVf95pe1
AD7PgLcTpKs4XiAwFuKSMaIIQZbGcAPs2mziihNU+RkzJILR7zBvsyId3X6KRB70
GN5a5cR+rF61JLEEo+kOwzmu+SbxKsdoZRVpHlsixcltBTwg3Nr4qPjVbLVWyAOG
sGA1/Sj4+wGOhO/9ZI71/Q8eQkUXqnrVvNwlS3Lxuv8JLwmrWPv1OlJrn6VNgsRt
3ZR4ohdwWmmCueEciDCEqDhnzid4TasDyZOPBOhLiwaL9Js1u8iG4MN1w1kv8MWJ
KZlCjA4bi9H2b5huLy+bZD9BnXKpUOnOgMiBSsYXJDDkukE1k3Mf3txogxTKxnKF
WkBvreJev9k5HTRHOHB+YyKZ/5CJLrRUKsY0nNhFj2g=
`protect END_PROTECTED
