`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f9jWInFoVLpJZeBTK9DGqbLYxNMfiauPQKSBhIbvts2dCjw9sEb1KlvAW/cymD7Q
Uaf19QYTaCOQrBobwCkW4P0ps4sCG9d7orldhvIrn89ZOtBN11ZVP5+yb5n67dEx
yS6mUQtCLpZ5VURsmw/MpYX1OwvEKKHykyHY+iKJU5u3xLYjAVD30eO2MIne7PfH
1Wm5s97ZETnXt/cw+tBNmBU0UCV6su5Ot8kkBPZxm9SOyFHevnWhs4FIDyXfbxHx
qNAkKmNX2szIRrexWQP5gPzF6XPxuHrMB515uytAnOpE7HhuvKm0QeOApyVYf4yu
fmj90k/vqmRjJA+utzdGDyfLbL4tTMV65lByrmBBZU00B23RiVnEZCE4TMh6GNK5
OND8qwHrihxuBnW54ZECGeH9cezn1pp9UeTpdHp5lw25dfUy7/YjDFHxm5OI/3Kf
drHrbxLrrAuQJlMJRXuzsK8dk6imnbY+gXbMpedFm71vGbd4jk7m++vq2Etci/4E
6Qlz5RnCjGFqg1yp+GHjbLvyaYjKPlM+nfT5uiDMTsg6yEXYDcl3H1SIpRbvtylV
/Ij173d2f50ugHDfiFRFaumOc7MG0T8NzO17jcUWrlLXUP3owJJ1h3Qu6HJhWFVQ
CbQodNgj/B3A47avBe7fn5G7vKPY0xEfMT6bAQYTzyXRbReSrcEMrUZVjF5ztGGj
8ob7eLkbFJJzeh2aoBeUJFSf8nVJVP/dqh8LNoIKGBDkNCcjoNOVQ8+HcVbJBaKY
3I5wtBmAcRCoC7g788Yc3CzsADOEYz0hmTtw0dh5nNHQk1Pq8mEqxpRtwg6auK4y
jSYweKQPwzEkXAUhkIu4zl4uQ2ZsQLo5F/PW2kZQ+DCe3N5zKQ4UlzIIMfcMbqSA
`protect END_PROTECTED
