`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IvhogK2sjCWIF8NDYKSGVGcNeLSLN7+hut14GAQE77e6LXNpXnZTh0B4qlalB2nt
SylOQHWwpYoIw5tXfKHFAXvqKJHX1g8983K/thHGo4AdAlZi3riH0BvYhzrgMdyR
8W9UCyV1Wfe5YgAFhNz9vsuW9tX53zoJhLwha0BCotzVAQ1ZJl3eF/nv3W4qXAt8
T0V9ndXmNKpT58tlg0AUU7wtnS9OmabtypMeCJrj7UDbUzvUxAtLcbnscKQp2Qfh
FNiEJq7H/2hQ2g4OglHwJK0PzdaRhKM6hLi/jXn+RU8P7C4TL69n33TNgUUYxoIP
UGGC53ha2nQh1wY7U8x/0Ve32TSo5/SaNsJ4cLy/b3HIRuz5LBu2zKd4h6DK+G0b
aBz1Ll3+IJZCxVn729TD5eyMQTlWUP0v7gF7kNwuSb5ylW08LsLE6KwMZby81Lui
vXFGdUj9Uat77Pz6QJet+E7tyXf0DFXz3iGnc/ALqTy3eQyQKobQU99OXrgVY0HQ
K4oMbIpzcvvaMCw4L92Rfp+OD1OREV0IkRA/up6P3QWbQjse/ogrEO+1TtqnYoBm
N5Q+4fhnhjnQqQcY12gJr8aiX70cHGmJBUuPq5IhT0dlOc55VabHJjNqXEcAH5J2
YZbOvScaxtPPfSzj7JmHVfq98gijsRbBFJe84yTxCk04PjoyHh8+VOS/1JZxrE8e
UeqbgKtdVdkNMq5O8FLB/ILqh9IcjYrOcwbFmWKX8b6/LY/z7N6kq60asBqSdjrb
2uzXJr6c1apjFlZbXIwGfPNggahacVzriBi7BMl19ZkCgNYC4zPkBdcOHA37IVZe
G8iA6IgtxqY4lx0QdKGofUpaZG/eUq7b/cYmARCt85CA2NXxbJYd5f4XUadyIVBD
p7diSttKV2IPbMOLkfY5LTBtSVOD4/m8Qba2g2LF/S3xc5ii9JHg13Uh5Bmk//hA
`protect END_PROTECTED
