`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jSk653J3PGUp2cG0RyuQg8b6DLVTUTawhejAs0X4xrrz5c3Qj7+JX+QsqVmx7Umu
fx19R7LWteDdzahNF5aDab5VNytvCYaNGsDHI7R8RCn586qe7JmK2/W6YxnKbt2i
TX7N+QvIjHChrmTI9MnQMqSYw4Cjttkvgykg4xsf23kFPI+6XjdbcDCWnY565kCf
aN1VjHyw/3uEpdVOqSbWKM+HhR63KMWsT+0DgNaTz02TNL9RimTR5m/y3ZAk4iJ7
HPtw6qHZuMweArgX84b6pxOhw1CSukLr5Lx4lJwvqDD4ZmnHR2T31PXymJf/vIHK
JovG3WS1jaIojIB6DKfsd3amFt1CBvAjKG7YllDOnR+WhawevqT84Br/rfjIuyee
FKLOt0HCJrH9ooOw4HvYebKr7hovFv/uPdCuPZIpIDdZtwGtZgTLFgEuNOlgnau9
bVgZtSICZkg1FKvMkVWxmlQeweBY/SZwjEbjAW3mxhWPU0erss5kW/qQr2i+QI2m
LeEXb0E889pJ5EONXzDEq57YXp0kdoE+HViV+JBq1AQwh+HMUwqDJhEHfjcWDU/l
pgmy31o+XOcL1/W2HesVzhZte7SEqfggRP1JggQwidaFHGOT/R+kADqxiWS4pNUm
PYBpbqNvUZk8dkgtQNRzHoecCByBdRMFITpscdyICoxPB6cjnQ13k2ZQYHyTkL91
hj52kMkjCnKFuqBcX0t/E4FLstNBbetqx/17uUQFtZ3f5x6unVdWE1A9eKQ90jCo
ecCawefuHY7hv2kKuAZ0aMeP5Sto11JrXNrvMHj3xdhnki+ZzCii0ZQBRFcVAJcz
njpt0x4A1bjxL8rzRSWaPD3sTHkQl+lBPrnW+kxj05AJiYz6oh91JEA2Jm265TUH
WLkDOymv700oVOu7NOOibGNskLiKUS+YyQs/mfEsOJuSkTFceRDB1A+N9TUT5s5R
Ryb/82AjIgToey1lI/9r8dAJPnR0+/PlWPq9EMjpVvXHaEcsLpdjgju9CaCMIeqU
wr0suFEiKUkt2frxgc/LMPPxTgNCYRqd0+T48i2VXLo+zaMS1ttKq+XgOlpPZHfy
dZIYm2THgzuSMzC76zeKnI3vXeTZ8lREnFpkMItBWZfdzHrMEKKW6mVva8f3dF/U
xHBRQBkADCoxO2EALsndtID8XYiE7kDosXrtPPkoGcF1yYPlpDQkVn+NkQ9xOG85
AcdCzzDqcsnDIthpjggJUNjNygJ7aXGuSGZhlhA5n+oibhf21jIDkxdJpcmHo+3V
xT5Mae1hK/4TT9i9uAcDtaV+nKkjZIHPaAnJTdSeNN4qDAL49Al6qfXEsOV/s3rA
9iqISVudN4Vc4ZwcmiA30RH6pAXO1yyX5wig03owO3QdG27RwkGmzTBnae3crfYe
dSgQvpoyAd3eRVFxplW31HtI4rWXHGgCLcrG3wvcn9vH6bEvwiDNayQzKFf2wW78
k134cGHSqj6xRkOeYRL+Pba/2hsVzhHoSh+g2qZC5u2jmoz+7zxEQeGvocvLtmJa
WeZLytvAs2RmiRHhJvCY3joc0hx7D4uaYZF30fjoKFHUkSUndW+iPFbiQ0s9s4Zs
pjvnz7QGk3cMLXSEGLk5eH/VVFSRI8AvEqOIcgV8OIGQjgY3Mu4BhLX+qmim2sBA
Zw8WoP/2VropVgBLlj2A/Xg0h/TElVh1pV3J6AWh3UOhs3qsIQhF8UgWBewexO7G
1cbUQuAARypYvLSxIeSaXFUF7xS2/6kVjO/QSVZD6yZDwepawHMWxBrgYUSOELXb
umKuMY75o0o+9dVUTOLYvkedy3xCILO7MyIrseh849fYdOOctDAnZLMu30RVLWwP
cgSsEteFF9j6rbGpY1pFfpC3I9G5FG3UMPSJk7qGeVAM7qyevrXtnZjQRl6vaXmK
o/cB45BcP5gbwzx4iibLhJCzFYjDTtwGJvoSpx1QQkoPq2KUgzDjKIMSnmKePpCX
Y7O2ad1FIEjU6Pg6eEf0ccL/byOjyR1vKbNj+Wuyu/GKBhqC4OUQS3KR/IbnKGSh
bl0gMMEXHfCRAfMVniuzTpdXvh4XVmdWBiszO+nU6UdryAnrrvnSVOO0RSis5PVi
eSYdHieMK/4jtUpgdUCh9UMtTFaHco0X5JJNnO3LKMU3y+OSROx1CcSYLU3853MT
Mq3P7TQb3720MWSa16JHoO2VWeOsSVFAOmh6MZQsr/mka4vuWEDUuXZ1vZjgBnko
S+b4ERYG2zuEP7vuOtiBkSiz4/S5nVuzAFeWS2XRsAsvq+oogQsPY15L1Cn1jz07
OwMcnouDfN8ZUC3pv8Y6fTPip5V6TdWU5zOmuPtaEm5CW3DK95AuKS3Wxx/2A2fP
xSlv85RoqhOtk1LPaGsNyf0pntpj5PRAbqHAfM+cjFfAX3N4psolVSK5IJkLBMRW
tL1h4lY6z3AvMdu5/ua5fSqe1rdZY3m2dNAkeFwLgbZAvv/Mg6NiYF1FKB89EzSo
i9LFSoXrK5dN/5ZzcIX+THkBUd0B7FbE1HcHmuyHSkE2u2RzIaVdiIUt5gIeWr3B
iI/qNUkJ9UuCXH/dH+B/OjVlM9YC2qCQmzQX/1xon0FsWU8DuEXth/JAoaqNJLpV
u4tHecPRmz0yc+bWYZAUXb7c9cKbBS/WxdQptUSMcsFxeF1sKBdCELHLZzf4XlNZ
1jX06vP6aR5UFYWfr8oNROIUPdXPYl8spn2EcWc+4DRNfBQoMO+vWRgSdIp5DAMB
bfMLhi5q1mkW8ley30ZvJ2wINZ8ZHizw3F2aj+Us3CO/vhaYs/ESCPoeZ1Sbh73u
GH7+nsSWymFphCBA2UBEI9WARfSPSN8cFxW0qsiT/N5/xtG7pHCc7rxj0jZJknic
7fh2yCLrGPJ6/Lr2f0D+qx/4UDkNnyC4NLhRFWnXWZSnmnBMiLKbj9rAjX54q9Sd
BUdECBxlJqHkkLi/n7F0bsxgOD0AiyzEANAbgom3MPrZZaJC8JOsjawGVaR84plH
o1uKz2nrwy/yESqkh9Es4y/aqh/cmP9SuWCFppUc6StkjCtYYpvBAB2+0EB/lUvo
2wWFotfO4SVMJ1DMUxR/CODabTmJZIEtK+7L/7VlFMTTSIv5ZBoqIMJFu+8VENCF
/g8nmWamoIO6m4wawUWovz9T2E/3OWOpRB4UUUH5JlPifwsWtBHaP7Xxfpw5HQj6
bwe1Ej0idBpEAiu15j0Q6SCcMf2vTp1kBD0XvsGbZbC9ds3eA3UXRLngcaLbOBM+
aY26ySMiaPjRUv7Fc7vHXfd++IqNXjGGl9l2kCpNQUdtf+nUNwTqZwTkzKDjD5pb
kU3eeQnGdX72ppBVdWjI6rsaZyCQjqE9JZb1sJord3Slu1jdhHPbctH0F6Sv8YKr
X1+sQf6wZu1kC++TurtrGSykQLKAMfnsYgDPuDK1dwA=
`protect END_PROTECTED
