`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kluO66Bq8tgwQMpbM6kVfLy+1/bPiQ62QPEQ/BOI6oGPFbggEEvtVyms1SxKS2Sg
BzTdlhlh3at+KequdbUyQV64VmrF3KMF7easOtNKmwTGqOe7wwJRBPW444O5VPRo
wMIiMXeqUL5zA/NliiD8Kq+95/eYilMciXd1nxdD2TOVz1j0bhM75XdJsAcU8hlH
cuxu3f7kqqkHeqzV9KSvEZQeJ+U//FtUoyz4KeyRQlrJ5cwlXFKPCOj7LlFq7NTa
zyFl2tezL2/0ZRtQ7KzkZ7c77HphHHKExoUS/8KFLlSrGnAar9hvosw3JrI2EtkT
7BG/TehCgHmF4muJZ+bwuCvWNZ+IkAwYS1O7k9Xd9K49667LDksyfuJ+Fm7AENHh
JxewrpYOXZbLne9uwgcrGS9VGCO0OtlPO+dK+xjXI+IH8cPkaEd2m5Ea4wykvMEo
km9PVq46f9hXU0jlMbvxag7fzxUEJOyj0DJ0rAKJNTQSdXsvCVSOLw59v04RE1Zs
8oSNPfFAshXg+qdKzYJb7YK9Sl4Y1OMBw5jhymOsCXg4VlQoXyQp5sf2eA1UuPKr
nSUSbVjKfRqNQkUq3iLmBrqrxxEtHukYmg5Z+73zuAm8lcURhEd0uuSDOK37t/MJ
`protect END_PROTECTED
