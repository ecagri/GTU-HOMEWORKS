`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
65vIgaDdt0dc/ih6eqCgk/0ZfyT+ejTc6ti5KETVXbi00AaHVatW8iZx+H2ujBlO
ItFQMVNITGr3i+Vb31DGugdyPUCAWM4LkyTG/XJo6rw2kGo73Hr21EFG+SktVbFc
llNBYoxkebVxLUgtkYW46ZngpcNkL5VQO5u8H1H9sZcUDNzULMl83jjmMD/zXz+S
eKY38f5ZwvBtyrTZdaV4UtZSYpu0HaeLYkAXRHtmj06W/w/6oWLPhpEe1Ai5ze36
TD8DXVMg0XPSKLNaKgG9hHdI4QcNQ12zhU8xrfJ87rjsa6pY17mF8KeAR/Hu3Rfq
7C/0i7u9e1UIoVKuSB8BXQ==
`protect END_PROTECTED
