`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+xqiZaANmt2Ga6an/IqmZjootwClDX5JM4NNrnOQNRm6eBdksOX1rkp4NUgDLR8W
mdrd1bzPmpRAmsiOK94hokaO89p3Vq5Q+h54bopBF/81R9tOpb4Np6npyQz4PHmv
ic9FnyWSsM6nuyjT4JdhRVXtrVBfOfy4jCcfGrrx6egWcInxTuKchzBraVS7Lbog
LUiGgJyA0mdV+UtXeuIsyqdMI2G4SCt/ApqYdRO8R4jPY4Zjddn+2Z3ChrSEOeYN
FOg3KYyzHGdu3fCraoaJJgT8UBjD29QYHN+kiJENY3RGdFWhXJg+4RtZdX/nOgFg
yCw9u/6Ig8Y7DiugZN1Lm0DUz25fZH7iUdqkDNjOfEKl8DuOTl42TqJLO/oM9G7r
OGQB5bPzLCMKqr6wlnHtX/SxdF4yJsmAIdE+Cd5RmwYHWpiTzRUeC95Oa+rIs/C1
hksF6xK+Dc2wV7kU5U0NPdVsyD3Y27mHZMgTwxOYTHCXhak4m0D82XSP6mMECiY1
rJOEJdwTFuBEiFoAxtOpavj2kbl/WHgmlQJn/iGiu02hXIyjc3jkZzXGlGuuDVRH
KNDGXsTtox/dAHdhmRwnAKSVpoM1s1TZKyvmfiCTxUC2MSeA2/vxohCnq4Mi+vgP
KtuUQ2uu1g16qZsj/NO+CufNunxRoVZCcU/mkCzVLx+1Eu4IJtkYFZ5t6rf37z1T
fFZSDVRrEwxtN6e5DMRsnZtIOCeBf3K33JWkL5IjGokHd0/91O3ITojIsr58PZpL
vgR/p4MBy2+U7XGnW5FwVUZeHy79ivE5bN3TMTAQJGt0QJ8munX5fzgEe3TQxR6i
qvEM34mLFjHvCw/RtAcpYu9qfQGJatSyjvSSJnCD4TTKBJtRY7zyQIW14jws57vA
lZPcyWzI/4LVXBpgrQqFfLVprRQzxOPMLj6s4Xceoh7D5dMc8fs79ZlwBYGU/g7c
cXLC4DY2z6IApV/PtleWxNZQmMsgNV6faRPE08HxwA0FPQKLH6GeVD1aKR5RlRTE
TVklF/aKovYpl5YEnZ1j3phjHwBHcHLNSSdsPTr9/1CoGF/nlRPXhhRvzFv2yu0X
nSgr4A2AhUHZuUw0knGWhfjDMW7ISRSnSiM1yEZK6Wg/jLXPbGzK7w5/pCTTlXwj
wznSJoOc7p6irl2vWI5UtHhDGnWZu1g20/7WNYnHwJmYjzgIcYDDzw3DJRHTXDjC
bWgBekclZN9lwTaGKbp9ysypQ7KpFV/LrHd6I0LEnNn4h3qOL/i262aFUKQjGlA0
lyGwS+FvkyKjxppCm3PaWawhM2ZmqQ1/ruVqMXSN8aSKqJytI/Fwy3FpD2bAWacv
PzlGdYAsbAHCiVjU6UeBeiGvUvEsV/ntePm8zF6Q7JA=
`protect END_PROTECTED
