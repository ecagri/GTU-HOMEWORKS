`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hewa/E95xVkOpBZHX1b0/OS3hMnsdEC6T0OzgzwIDJ/tP4i+yC596vrma9qy4JMt
RNWhPipiqKqxjV+i42Brt+Q1hi0BzOjAwUhUq/t2+PY+dXF3PJYK6EkUegKPwpQ6
m6jlr4tN04SIojL3vmkzzXvkt0VD/mcnp22z/kpV1EqI1DVDcY2Cy+rMbQ0LJ4nZ
qZ9mgCdGWYN2DSNjNE99XhkSi/IKNbu28plRTDGVv2PUoTPkS/LUgyCRi9YI/JHp
ZstNlajG89c7PuPbPACRMi2cqJvtGstJ831ma0ceIAA1KyX4mWZATyfyxjdZe7sN
xTdY3o1UI6m2VQpcPsj92jW7SkZOBamUe2fHCfXfZHE0rEAqTfGTvqMEGzJhObo2
B+BiaFTPYhC4zk58IaEq25XCOsGzenXhK5C2FAQkMTEq4lBkn9Ae85whTI7vMfZ9
5vuwwJAysKlXWmIKk+Ziq7vNGvZademZlBhxZDdjKy3LZSObwam8xfuzlA2+X1Dz
ahNhVpu9ak/pvBRdEPzFf4IdmkfHs/DQA9tbWx+eMI+74JAvGHrx59Z/tj/aAV8g
QiYLRnO2sf1wo5keGFnTWdYkE/OqFmcB88loKiVW+HmwVQ2Yxg6Xt8DdQT+C9rKT
2D3gjB3oYL10TQahWknLfXRKRzRIQgIPcQB31wcJiYm92yMXA+k5aba1x3C1W7vb
HqxK1dB1rvbW/SCP88xMPitVDO07MWKFCZ3nYHpHL3PjtsGOU6YMm5aeb4TR48oo
LWPPtKDBT+EoGWNB4DZgWMU0AZ2+bpmmOlfs3V+TD34sifJArWbzslVVo3C7wuc7
FfMYrOCBf1nrnCz8B8xJJYSi50W0u3T/iWH0HZ8zdWvnMe0yhRMWqKv6NdDemZTN
YsjHHFsrZNsbAwotTMNppExcBEQpOCwWMwjbiNs+9s0wLW2xpl31laGRH8rqdUtt
5Z3pIZUQq1DvQ9PUmAoaFJXp+ydzrrLPpJxrZWjQe3SH7wMCjIP0N7KEslWJlkbn
Rs8dH1JilR0w8ARFnjHSV3iyOs0JGPRMtqjxRegAvZ4xbNcwHrdblSn+bP8Jl2cS
pvKhgwHZlKjHiauVU9fZozcKTPwMJeEyNH+mLHZD853kQQ+Bc6ePZ8xIqj1rlsCl
XpCuaACjs2y7GVssF+BY/zjZmzPRz6cPFH86xGgDGA9x4B2oYRqLRkRkwe2TnGpD
trzR+JWUyh8EQ9bgLO4toUmzBk4EMDjguvkjuIKnOl6Pt4BePJXPxRFj/fu3MTpC
9l+2q+qnYzfP+Gxi2ibFnydy/rhGeySNPIJk3GFnlPouh8g14IYrZgIYiWWXiBCb
eyscf3orDMQBJrQB9mnnACWG9ih+17QvQZHJIFl6KkLNx6Oa5I95qHg75wDcOXiq
My4EuWAcMvJZErTXUx0EEMeFCEzITLvYWEGNAvvgh78jhLUX6r+9Ve8aNkWnoJe7
nMGvVNt7+BnayrQLLK74w7gtRHEGrTSe72vC6ZSYm5I=
`protect END_PROTECTED
