`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
znMn9JKlWHwKA9VFBC6Eu2dYfagFq80j5uR4A1dfMuNV0BPJ+8A1MkEHHi741l4+
D4S2vjbqTwcvIdFWPDl2wTuwUOeuCfDPsI5IfZtGq3S1xC+eBl/34VqQot8cLvv7
Zcj1LIwMIDDJAt56isghb0TIGZ+lblhGCAWQQwQ8HCGsBuv2vyNzALpOCf1IrMwD
zrIZW1KA5cL9vs5CtQFGn2scbLgHklpw0mymnYqDxxiFVT2vhRJ2YfXuPHznaDXb
QECwlPeVSYUWsj0I3u2ebppPwCmZgkuttPPnOEgymlFZ/BuB0tXwNRSXKtWAwOG5
Hy5tDosXzior4AZiPVAalX7R08BaJ0XnTnV+eM4k+d2N4y5WD6gMs5iwWl9/JQR8
GhywYefxOhuw+FwIZwOjwvGj2NE7SF4buUQcf87iCPb4e9G8EWJ+4Yr/U3utvFRH
yi+JGG6KBkh2IoPQ2Dn8lNOZzd1uBVOTqL1Xi2Msou9gRs5pKgINVB2c3bKbAlW5
mEh16/mAev5fDI9TJIk0Bvdb1gDUI5aRkOV46qJfgHZtUQ+f3azBa+Sjc713wivb
93nvbpadO9fgIgSWA9QcYXlLBImOjtVntt8HpWrMIWIuEHj6MnlwWYQ71e/l1SGL
i3TC21y4dg4MRV0z6l+j2mUzux0xXJeyrX2tXEEfNv8apqfd2UIYItOQFLlxd4M5
Wal5O6I59mS/1AERX+vxnBV0mnQ8G9P4UWs1EGwhXYfVbvsWC1Gxg2gZ4yzkqLKz
IPNv9wdyOohcIai1jabAmSyP/RFoEX9b6GKVl7EfDC72O+u2CU/18tYx49Mtw9V3
mu5ldEAxm93C46oWRbyKYYOEbpBpO0lVAxzWKFzp9SQ=
`protect END_PROTECTED
