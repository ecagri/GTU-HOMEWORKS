`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6ONH2D80IFcaeE1c99OB8jGHJSGmtCeCo+IWrKTRMJByL6HCvWPetUt+5kh5Kmdm
WKqQ6uezUu54SNj0kySXf8cOu+cyDrt6M0O3I8jF8suLeAyA+HFGT292gQACoxEb
Hn+/SLVBPHz9V4CFLIy+SB1Ux6+rKwSMR0H8QfdYiIpJ6DlCWeAVnaOKOfKl38ZA
JMgQEmpLwsAyLblyTTM45l3gk3Bpix4tRyiO6NJjc33mfYJYPnIfMKK1h64Ec2uc
tALgx+3zC2diFXuYp+16qKknQOgkj+H3uFTPThz+ftvLPmlpUPmNPHyc/NsVYdjP
8acdKaZziH9mHbWqDglRpVChrNW7AjzJq1PSxCjiPhalBYPuuYJxst2+8hMXCV9a
gPDC2ZH6mRNGHks0BcCLRxeGQyN0KY2NwRiQWyYUFAQm2x5v66Ar/2GdRynAc01v
S2uw3vMP5Kp5EjwgnWW5hjbQ8lGVSiuWuWiSPziWJKKY0GNnFLv+ElFwjcOgq5yn
umiLd4Y4AmsgHaIoDaOdmWwl5fJ95LwAJQNv4uCOI0vtre9U22UFN0jixddG/oHC
WRZKXKZ6sNJaQS+Id7wm3NsirXWHoDNyiLh/BtcKEpo=
`protect END_PROTECTED
