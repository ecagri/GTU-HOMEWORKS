`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QMpS6Fhotqn2E7jSCIDMcP6IyfqryFKEheBxl8XBHBSIGnOW84j6yZRganbZzUkX
e+YHZ8ONoESs88rZnKKovpMXzZoslR/upjNJSslh4jYkgUI5xNVcg3L4pnbDewgV
wjOH6Yj097idiDUxCM5u2mhaV9n5yJr36YkYyioSW+ikuOLY0SFNHq/A4C4rPGvA
CcJl2Q855Bi4ZDusIFGPUiU2oJqKmAzTpeLlq4fZHKHqv/gFaJ5TPc+2gXy8YeRT
Aw66V2u8S6HtlZcE1J0NAgBf2DZvyfph5CVAjH2neJjZsfdgTyylSc9H2sPChDIa
02EiUtwuZmJSnM2S3MNbTxZJ75w1fURy9czVKjdvsl1yc/ur4eMJbT+jUpDpT9Q/
RFo9ZpDBDye2t51pWWIdkLFpGI2g3tzbPu/ZLJ0sGlRUySwSs6R83LW3rKhnzwHp
s4JJLL4afhquUVFLKt5sNiDFwjZ+sLIxxBL0ZasaLE34/5SPViNh/xSEJzg02zwL
IadQNA5lnagCT6uOw8my9uCwuV9RhcuKiCiaB/hWvZD9mqNfq4W1DGWYm7s5Rk+Q
h3X16JR/MXWlIxtN6HN5yLAYnYjTfeUZdai8sscIAbA341BXGQdV2WhbY+BKiLDK
rC3qIJDkiIKn8PLQIL1vo8/tqFdsarOCVEAf7aHfC1jOZXFRRFNX/Tz9+SO0+f9q
1tUKtvlquJWzgKO33nU0iy46p/MHeifQvPgB6vDmKmJ+ALWfs8HqRM+ic1nPCK/Y
BTe2QIjx8ODbCgmu2NbMtojXoebOBSiKdigHbktCdUaU1VTNG89Sg7faW+dX/oEz
R7VQU4PZuua85t3W8YqWPwiI+qxEjzMYkMtrWSDTNEWPIyFDm5Lzfrey4ieKExrQ
NqW/fKsD/Cst9UCTDixefL8+KRloSGMl9wHGhthyABe12Qjh8tf6E9r1gUOJGAV2
C/yCrMfNdU8WoNADxGGsntkHdsiSnkQFJI110COZVrrYiQ5dZITrhYnZAt5FOYUu
DyWghNH70yGHtHdhgiAYtvwyu+E4BRopEBjiVKhBUfpAgg2KQDrxu67RxevxvIwO
GpoQEUUulKcv9x8mxOxl2g==
`protect END_PROTECTED
