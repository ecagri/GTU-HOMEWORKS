`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8q+hpmbPMUZll7qn+c5uvsvrgr6hEeSgvWBMAAAJRUKMzhHa+cYsELBHlZVN4JD8
0xA+HJ0G+lk+2k4lMSAxVCkuJV2+C766QCpNHPeV4O0xCDwfZcDoGPIYnxLVdYUi
oxKASHiPv63xSgVfQa34fMSJSDChWtkubyzfNak5v6djtRCC3NkDJgLnrk91VwCH
ogNdvyYwXlAvMeQVqTfQRcSdLfZ2XQLGr/GlMcMPs4BfbhMQbuukqjTonWmSIc+W
LKSlKbefxwuksCp2nquzvmcaTNvLRDrkO6TKv4I+Ndg1CfmNfiV0SvKvv/J1L2cr
XC7Um2uDJz+0nzWg/iV5cr3+hyN5L3FS6S1+7wLWFHcSAwcBnEikBbtkvZ1y1S2l
qDb2XgP7y57ackpoWBofqo+XNFIYzLMiG27KONM+2mtugluFOBhz1kxlp/AAzLSD
JYixZeJVl4MMaE1TVDEj5yc+bzjaAgqCSvbekKVLQKGXn2R7WzOmGZKYHsLZXg5U
k/vCTzfjHdI7f/te3X65rfxdkhxOzDe4n5vM8S44RCp0TWgN7mhOAJpBxcTVMiaR
GlbCuR2p2PgbvEgKDRcsFJBWEc9lN4CHttICOuu7lzdFvcTnHtzSeG974jHGjvoq
ryl34Zoczizk+zsVGizzwfjH32zL4BfOmxUmdwRzvM7fA1nBbPjAGXUJ2jzLk1WE
gIo0FNEECMAGr1dlV49INpKRvKY03N1YP8IHLBVH/Y8p1GqYxjPX7eGABh4+yM9J
m9WfJca2IKqywTML0e93AFKcmhx4SamZv+lyqFoMScsoDFG19bga97p/mNo2mW/Y
rgNTATEtbtaeaRfH7k01/cg646RyuoXP5xtwrI/uBmGyJrEEBcgzzJEGYSSt5j8j
DFIP+uio4mw+e4CWrmRvLhUJmdxo7VjpHyAChq3AYNAeqw5QQsz3M8K+qeLm8zlX
8T1ygMlrO8pyLKdDiBcBw02kVb0vgH7nUts63W/28dyqaJceOrnP+Dms3Mi3lopZ
qaAJ1peq+pgtV6C8ROASEY2dBuC+ei8b5JqAMMZenz4SP7WR43QLrXRyqnxX02M7
fNUll2AmLQ8ZGDbOE9MPsyS99mXQOFasXrJjDrV5vjMKYp9iuOzSvNiSlrSxSMCn
kGBwwbBmbyGLrigqoA/Z4lTMDvbVyCz6Uy0BYo6AArjwwpkgahjQO2rf2+iUhS3X
bflJGeqZw9QjWZbCHFQTO+i77HE9KfSXZpd8Bk7b1auROpcv7fwY1vNRm2Of/XhD
H6KzSn7iRss++WjRtVtgvVl4q5gZONXAO2Z1wA60cJBDWFPEsNpDXmtiJTmBizK3
dAbS2J/Drgiv4fkvUwntJF0+Vr0kEAMuRUUq+IYMuDY94XDQ8jdaRMZW93Yb2dxR
YRqNw34hXpZztfibNy+tV2c14w5S15lwubGIBm3zjGJb2x2HsTfbuR1L0pcwO4n0
MuBw3DnNLRat9AVihpzPoSZEGg4xkJ2s3I7yv9x25963M+7x9s61w+YNmx63ibGb
MUXEE55tprPf7UwW5FVgA4uACdxfXevVIz/P9nhPLfvbsBxtwmD+eEKjfzQC4TGE
0k2ujF/fvRbpiaYjAFZaN1ezoYVwRXX5Z21Td/wo4t5aRXYJWp2CjUnR5I0Ibro8
5edEE/5Z6asqachlLbitnzqZIFk9y5gRzQT3zyA4+Z/jTLAVd6Xi9VeObc6l4toD
9oUUhmxpkEdb6v7JZ6Owc0n6RPAnLrvf7i5+6XdSuVr7Nc96AgNPvBoVVEzPQs6w
ffKWpLqD3DE7yfxR13PogYp19EOfAyelq+j+/P5AIFBovxmE1KKtIKL6G2tfQF4+
vB16EZH0gMUoexX8aE6nbE4bg/njz0n/Ic6pyaq8P8hz2HZZgsiPqt77Lvjt7B3a
xk37GMgHa1kJyEdcDf3zReFJqnHXHxuN18P2Nf4C6DRrxLNuADh39wSxqeho6Ubb
Au6qj5DWCYZ3OGztuQAQvgq6rlB7S33a9VyEmis+5vtmI9cVDJ32UgXsH2zD1Mh4
VLwTh4ozr9+yg79GOzr09f2qYKzS6TIrp4wa27sybIJLzsYLtt/PE8N9C71HqR5Z
8+49jC3BwHCSLDam5eEKssAhK237EAHo2TCYloxDjNQoGzJzHXTrg9+vh0NT9QW/
1IhSQC+DFPKMLNqlbNBWH6RnNp6USWD+i3uWTSAwQeXBDW/Q8SrPVkchInyrO11a
XGML3CCw2bbeaFrrykjGI/kzDCSFpgtOLiX2xuPftwR5Zc/Ffq/iNyKCMwq8Vvzy
35ITARKCiBK0SSi/IanSZZMmlrrh9Wph+iWRLnoqyyEzHxbUXRNIzWU2ai97pE0e
Pu719+pEgtf/OqReGyUSZjAOHfXi3CmA6QTwwJ+WjeEN4MTHDwVnX6w7isZZ4AkH
NRZ0v8Ud0a0LRTVf41tKpKrNSKKGXuhcq6p2eDvXvwkBUHpfU26FnS+QjCmvUoP1
9AvvoPwmI7eUMtZ0ffKuDcCJ0QoPMl2F+QN0DZaYcmMpKrgOFGHfZiY8znO3tVtU
19npf6X6wUHVQc/LkNEJQaEI5T26Fq+AzA3Sb6GEZHwLfMKDCGqq26iroWcjyelO
KBak8brzEeObWqWX2o2q8v9psy7jATxeXm/+JcPHMqoS1jpEMhZfWMjLRK7GW9JZ
QGkVqIYmmBwvBSlzoH3zJI+XhIhgSLI8Kcns/t7IZp0i4RFTPD3r32sbkVZrgUXf
vmY384vj1rzHOwzo49ljelT6S9GfT8KtZ8179SXqZ0tOUIFClB9dgqIWDvmgmfJ4
2h/xAxOB+0zLMIr/qi6hiIOB7npPPP+cJQ+jBivUhgsc1v8B0/NCmb55MuGjTx90
g/FCfYvZE+hw0JvKXfysbP7fyvoc38B61alTxhoIB9QqMqPJHU//VH1HNAwpBcXU
7zOKwYe7Vqs6rW8d2Ce23W1VSm4O2DwktJQ4qaeRirNqIPHx1ONlDkvzLnLb6pWI
HDwK6LaH9Q5ldO+2TsYacOzfaY+QAIzaH5EQ4YkkGS5UE+aOur8i+lPkLwgo1d3h
H6LnB57r517t2+8ynm+SoB6xMdbBfBaJa+4XdKiw/93jTHOWb1PSMjo2CZk2uS0h
Ni9k6kmSg43/RKm9Hg2FIJswvCraj3HLJzNc/Vpe/DSzKG+4829soLjtpaYul56E
CfCPDl4FHGdXrC134ptOVahup5vs7Z6QujrUwgcwK+s+DAyz32U975MqBj8zv+ns
2j7A2ESCyMkjq2Y7friGSzzIZcWP8NuIZTHmeOhC+R7g9CBwzFEmy2bYvTenlMH2
hxNueuq15Ao3olmBPSE89OE4j4g9q9yuTSuzJVQOdRskGIyiS2phoPDY00OozTyQ
5pJnFNvqZHo65nEBExzgAKCW2kU/d84sxjAOE1/csM7+ML48X9QUYG0X/Lxp7AaX
F1idHTrRF+I+A/XJiqT5H3Hom8oFHovYtnNhH0cBsTw4HJYcTZ3MpQGRk2Ne8utw
Ip1V+Xs+LUSfZoVsRa9jd6jcv2x3f+M7JDFTB2+keakC6WyjLP7O/l0Ly2PXZ5Ap
X9SkGAr5JzzA4B4yjQzcsQtoGGB0i+kvjWUNkfcbtjhHaPhB337uUz9x9UYWygWB
QH0+P7ikmBU48AV+lNganeUczOMa2zJuo8uvvPXD3SaZiEXaQvRzpUz1+Bl9gbzh
cxt/qP1dmShH+83glVEtveEmfLBlaNJ3sVPYxR2PygmLggnmmGKz/aNc3MG/ZtFK
U3I+wq+7vPkPS1adIZ8eGx3l/Dpt62d1+W1Tu2UGBAhxjDou5wt0waBi9xwGJE50
ROliLN5FJB7DD5YC3/KpcQ==
`protect END_PROTECTED
