`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mNv4Ng38gEEUjkNmMtSOZ19jo2lvdkjD16Ln3vgsd7NzidR7U8VV7bouN7NcJfiz
863HjZuVa5pe66RAzitZNkQrGYdSpA2PlMV4+ij8KVUhmM9bksP0w1QIIAX99+4h
j4Ix0RvbxWynvnBUJ7YioqsbDAR+XukCmbpYoWOEWzRv7kXsRATl8nLI8FSFY10C
n7b6P9ZwPpdd+nQZelxruQKcOXuVOrjrl6HVDfKWk8nc9JNyrW3+qElvEmk9HdR3
xdBBI4+/1e6LJf6ueMukxQHna6YYZQjtDx56rBaoGM6mIXwZv/qfmIc8PfEltMhA
lIkGAeoNtPTmg8OgM7qeWxy6B6bbKnfQx6nl1ER6C+GkZ+QLVabHmQtzS4bTZ2b5
/TsZ6OOBCdXsIQKl0ZTyB4G7Ysb3SqzAgTMAgwn6YnzvqGktWG6NyPdLThbgPMGg
oKhmEpmgHqaX4ZiTs59M38B1dhvM0LtI6GVp1az8qUrJNztCGUqov8RFdjlxd4C5
iAMxgN2bEhVCBaucTDEh8kOVg4Cx9vRn3NXIAkse1reR1PyaGffqj42Dq7UzsQMx
i5gYcuinPGc8gGGPPA9DfHPD6o87Tjef2rQ18aNO8Ak7XYdd144jNFN96QmFyBTR
0GbcbCGS3L3u14YL6Er+xlJk/1cxiz7WDamhoXaA+WgVq5MojxTaII6R8UzGoovf
Ixe0zMKC6uc13dXdvrIBWKngeYrIRZ2quXp5Ljq6Mk9GtUEWSefPlFkW1Jxn6esl
/GDcGPc6Y6kloWbHVJj7ur5nbDR28v6FUzJufIpQdDXcgrECJ4GP4LbpDCfQKgmv
cIhLUfJCxoi4hhhzGwLLRYiUEJ7DK2V2yXzqFay8L7NTKkeFWEKdI4rva9NtfNv1
rKxRBzGDqHQF8TnwCxNsNbzdEX3HIpbG09/ViWfa/XNJcLxhtBZPQYIvEL1nZ56r
3bJCAvPNHubLLyxZsLAxfyeqJ05cXALxRwbjw7M9i0GFdwgCf7hLF/KqGPvSnNTm
ShfBp9GSJTexV77dZ4FoxYmKhfbAe3cBCAxvuetbTNiXtiv1oGgFOQqyxKQgO4mS
rBBFcZzwORDXBk27Q4Gqn63xij+5NJ7zibnqSBBeumOiGeDeDI39V9oNzro382ql
r7M0QNwy9B2id//xtAP79dcBaUS4craJDxamMj0gO9ErZUw5cHifN0ZYy54SIr/G
GQnOA2b3uF0ZbKamJlDeccxJ7LXlXrQCmi20TlYQ11KyILJK5SfmMVHfaCZ6LBkR
CAIXgCRVo8BQyDAO8SkM/ZBSia/5SQ4qqt+8MNMoC/ooy7YbdOeSl4U3mNmPTmgy
hOQ0EvGEqorIpaLRPXhyJOnTgwqnDPYE8blDXoykIADgO8IQXF6e8rzlSpa/TmR7
WQdwyZApOc4V+cdmc2wDxCVlmzmgZ+Nkplq0FD2nOrjtDlttPScwChvi5nolpjms
0Z4AQA7Ve6rc2owDMfWsQS2UCAylDfNQX6ScW6dciJbQN9BUcspFNdagy5Dob5no
DB5AQWwv5e7Ybs0VkRWXeHOUqqs2D4O6m5tG7wqIHaZ/I0PZH6MrOjg4XMUuBD9J
t8WAooxo/WbGI1jpE/kRcFLBKPvrcmoota4FamUsfG4q5FEjg2azuKGnJcbrkWe5
f1iJNrgWB8yZ3mDjge/v5cFI61j1+9cLOzi3+6yiN+urLUhZXGszONT8AoKu0Zj8
GQ62+LmaCneJIRZT2TRGBFNpxT3l191v+LiavSQo1Uk=
`protect END_PROTECTED
