`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lnSBNy8Z8G8lv4lLwDl8Xqvs0x82Jg/0kE1uZNHfz233gqZnKazU68sIm2MKcfGk
TP9q3ujSzXDX3i2n2ulLFIoGh8XR4feTeeXnB5A3BLi2KL6wCjZdre+CwSB+7Hbg
ORdyh1cX6ieksKKsLS2uZc85ZeiHioNFXlZXsJTLCHgw3WZZBjofN3Pl+XFDezzu
kih3Qi/9zsjyQt94E2oBTfikYPwy2lZ0nibpKwc5mk7WOwEvRxsbx3kcdeqmutHd
s+2VzKZO+mvSCUebaZ+T9pbtpLIULpOCLvIBW3j4npUqMZV1jx3/ynSAjHeOQZrx
9VlBJ5vmd+tBOBg3lg97JeO01gELi1ZUg30bAkmusiihez1h+tpg8uNnuzsjhD7Y
SwilxefSVeqgcyaep9vyboGlAuoCr/jxUqHII9Tw/F+2Ikakuz7VXqBRDuqyiMyx
`protect END_PROTECTED
