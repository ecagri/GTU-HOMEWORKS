`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PO8+SaL4fKF2B3A4/9YKhBD7C3BDxl7aYIF0M7rmx7jr5QXniBA7bUEnlj5dom1C
VYGKiO3RSV97US2kPPY9eNsxIno3JD8wK3OUrkmuLEyx+LA7Bfj1y2BLONklez6H
6cMYloI4/2KWRtrm6q3IqO3KKFIjXWDuyTSN2pj4FxtwKnuqZHogw1KZr8abIa0C
jANWLBiryEiw65DNVLWWeEBXnFhnXtn56ABSwPFSKc6X6BQfo2HkawZAVig/yFrQ
XeaSS6Q5SjlpV69OFC5UbmGSaTBVB97dl8lINokriDTeAUuJfKv2UrA2beCnqdbZ
YEoX+TFRIvLXBr0yaDyKhIoM403jjUqfMfh412S6rXP5zhNMCPHWMzjPWMqRaSA1
uVr6NElY8RBrE/DqCGunni2ZN4W84cZMo/5YtbPUFRTu8FFYUTZzyUAqiO0GpeFp
SinPxwBtBGifNr9x8TNDBu/RHNQqo3epxmBQRc7ZxfAqFphj2NSP+u+CjYtx3NSa
`protect END_PROTECTED
