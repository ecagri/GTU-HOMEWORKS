`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5SAZByM1wmeHjaP00a5LWj5s0FfNF9dnKkEbbBAAcxmaLvtl/eniGqb8m7TyYZvL
OPqzwj5hoeAwkbkr++wr9E7nt7QXlMbBkN99gKSW0Qb/oqlcfGpbW/XldZvFh6Tr
PIVWUiJk/1xB3nSt5uoK0wHT7NCpzW/Mlzan7eZ3ll7thxxBNdnz+V8YX3csuJfd
N9532FLZb0HpE1BKZP9/9R57shuIE41G8cKZfb1rz/9D/nC/+36tmPj7tjvZFQgR
NMigePatzAxml3/CSYpyS3uHtDWISgZJYKfIh49UptI2Za/Sc5/Fg45GpltIT91c
nuhJlWuXXNtrACnD5KBf4hD03R4H9vUz2IWye6bZMTwXX84GFVHTXHPUcBUPPGy+
zPYb1Wg0R+rD1zCBIfEmlhGmIubKKDHGRBhPDkCNR/LbZ6zjByyqlndLZGsnIgH4
jvtkejI9LyWoGLyNuqCslUVTEIH659dtsAgAZQTF6637HFB/tlx+Jp1KJP3e/TTH
yz2l8UG/91wpy9JY0X3WdCZ2TnSVhMNLyNO/DMBUdAqb40qnSi8UnyKGcJDhn+SY
9qijr7fNpR585M3Fv61LqZtaMYM+A0mWceL3ePsux6lsGVaR7KghBaZ2MPXJDz3E
3ph7/97Q6zk1bNXm3AFhMLccFQW0iqHBA2In+GJyt05hSHpVaYWxq8ym7YdCR02M
uyMSdva0VztACraXswnQFPQNOG679mRKwSzrjpMf471fZQIsVkaUBPevghFQvGRc
BCX8JLEGqx8VaeCTWMIg4RteZKrpt5+hPhn6vKB5O6ArdfDceKuRsJ7mNZWPbhee
cjBmO5mgQTez+05FFpXRsf3QlTEDo3a0hwttHcFb8Llut8yw+jby+W3OXgVprDTH
QyfgY/oV4RlDTCFvHnxyREcdEj0KSZhNIMXiGSHTpozON5iDLQi6lsSMZB35Fsvp
zfcLSfwuO0S3m54MvX2ftby2HsIym6AGX31CW9800x0OISoIk3i+6O9bmQs8csQB
LSUcDuqKbFZ/dfForcd0N3pvAziq+WzMOyoIL2L22LlBG40FqdUEpEfXZelVjzY9
qJDgOkosst5i1x8gF6xYKwM7KuVBUA6xjnSM4yfgongDB8MpBvdPTA3zO/Nc8+Rv
Rh/QYC2bTw68HW7TZa/meQP4p+h++vBBGGFWWUgsj7pk3/BqEqzzCh4s98jgM3pF
GZMORj2pOHjw08xmdltugWUmRjzHYMVllvI3hj3etFWH6NJFmXeaKo/7KRFmklnP
5S5coWI1ZvXBoR+n4RCPS7Wx4O23g+KeLeeM6C6Y0DGnjcISZuqAAZLAGmvxVgo0
RwL7y2aqBYcx7Du//EBYTNVbz+kj7xgxj6+y5OR2G8tcSe66jMEuASYLmDvDy+e2
dmHJNrgzHFrX+KqwVzBvHoxwf81QU0/RWp1VS8TQBPKc3BArR4Tx/u6fLOWZafzO
YgwAYpDTYdH1Z399jTIzW1IRBhDt8vb0RyUCaUX4mAQ5oiDP31KW5yx2dQNWK6nH
LBHj+u/VZ2SRXmi0GT1BJIYBY/6fwHAFi636XHsJY8U3UyCA9DzOtxuvag7t/H/C
a/zacYVF1Z6H/DIlMWQfbbu7z6AOR2N2BSIbnfYsXqA7kW+mfBTBNlKUfX9NP3Sn
AXeOYduDQK97CtJSBVKiKhAXmYdcCp8HCMFOVYKb5BrofMCWjXp2PQ312JznkF49
1iH+uy8sX+PVGjGWP0oybZr/HNCDVWIKMxclyud0+HVJ6KORtiS+iEEpoAkAOElP
AjyaHDpx0EU+LNXcbBVEtFMSbPCvgHuwwlElTfPqKVrvsyBreAh5HErCaVXDgHHU
df11YdUszN5AM/qgkEt5PyAkbHbyC6eWTCKSewvtvJvdbCCKKGo85PNcUR6A8RUf
BPM4KrmMxxxXQ14ojC25VZQqi36hH99heMr7csV8NA25APbvPKWxa9QAdHx8oSEn
REPvRU1sSWzKg2PuSZJH6wBmdMO2I/0QxZJw92zCGxg=
`protect END_PROTECTED
