`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0rEptMfCOre0tI7sa8C+QFsdCk8DHtd6kz+OtXTGeZeKyAtfKN83A2AD1T2oCe8y
ik6BR6eMsUSlbpvTDtD1Gl1tPv1OsGlC00VLey0ueDJNbasrtp7bRkEHoHvXhauK
6FbYQWelGvEYSQadlgpjyIvE4tCOCvDmrHWwIJsw4cLiM9dsh3KErYo8201uXgam
H5nZzLpjLjWQC2J878OjDdPu8QLCcwsvg5AWntlyAqzkdmziyohpHNLKeswtvFJm
WjG1qpHX9FZMYWS68A6koBUGk79CrO1wUU5VauswoHV9OZzxipRb1pGn+wpPvqqr
arf6h+1G9OLd740gXuOfjFJxVE0a+7Af5n4FpAGQfyTAXNC5GHmj+C+gxpWbwMnj
6QlijZuVF/NMuY+C2uUfdioaSbnbe1PXsa9DTIHY4lsxvjoW34r5kd//9yYiz3sZ
8JSqnHSAWgrMbRLaEuwdzxC8ICHjnf1zASEirHic1BrfCuMDkW9s6wVFs9xdK8oV
jMKZquNDBfTthnOqVm/eUw==
`protect END_PROTECTED
