`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e1mA/dVPOfN3jW3OR8ifAzNLsCflJXLVr2xogrq4H8Q4F3IGE3qQV+upTzYaVtso
rGmUZmHJWr4/AHBipURSB6KL7U5N4/seVIkuSQbV1+sLTJRVvc15FB8F+tldJaFz
KQdDAtnGB2IQ8BqUxYbKRczp3Ke2LqvMV45+LrB7/va19zpuMSJHUNLpR5X8uOg2
j/VEdNItBMgUsagJGItiHDNTzDhHEDSwfqv9c85/2SpHsypwI/yQzc4SAJIfAXHf
OBWdSSoMlDBl5r30gruACEqPmPRum/7XyRLnx+voZhGbIAGNXMb17Si0YRai29+s
dM5PpL2Pt4X9kBsQM/9Hy6W6oUn7QkSIklhXTvS6/X3o7MLSusS9mi7mk29QevuK
ezQhYtuXEPNAabdHBYNcK6Du3+S9+5bG6v+MZWG/l8UIx3tBPwogToU5EzONUxYC
XcCuhossc1XQQqKBn0oVaBWUpNVbnIYO8UG0v27YE2vzGN9FW/Mq87Tp68V7OpPZ
Q0V4BH/m8KZaRB0MIdo3MS2YNj3WFXie+g7ytLJxpRen/FAJgzRJHXD8FUIFNg4U
vRTllTKSzQy8ThpV3zeigDwdOXorBTd6jQHhq18JWpIEt32YSAUa/pT+ubpKld0a
+p9dv3WPCdl1Ce2Smc/Qz6Fx4C/W9CKdE0jG86ttyllmAWyYMxmuE7naRzXIM5PS
mo+lHRylYvsaRpMSGDmjfCbazCAQ3X3A6/piy15HFTmxkWcZdyifZoyhVjpYUdtV
vGG/+MjQHLjGsEYorpMw2gvyAwzant7uhiS9py2cbpL4d6e8p5ifizsAaO2pT2Fn
Tmrio2+W5SBeD2k6knBDCFw9S2X86Wy+mXRiS8Vm3CQt+ZRpurzMbuuAAo7hxVw4
XMtxP29IDp35e21e4mT+3hNY+A6tf+g8LePnJ7OByLVhC7MX+19rE+mX8MvOSwYp
dGakDP6dyc4mGVi4ysViaV0EFaZF7XUKF5k0JJveWnVLfvOCJngYP2XxSXddniO/
7dmPZeWIybBg9LPL9fJtYjWJ/E25GGlZesMQGtO60N3vlGaa3CFTwop8G/iKusVd
ChIH4MsF/nODzOnUJNMqoSSNWzLRICg+rZfCKZjRV5LyLfxvkW/YUK0sohIkpbGb
YZUmIqvE+OU25HEBJRRoIrbGuehhjEOaBOLhZgjIOdDRs5bdcfx2QL1AUKoa3uwS
4OmiFSbGV32nI42u5sfUQrcUJqGB1S9cNfOVncZNsODQ/XzR2Ebt4fc4Tx/2eEbw
Rbf2qjhiNTiT3rs5W7Tuf8EL3YRbqfkcPUsx5gVkCN3F3fl8kDhlXCKs18g+vErp
Pi0XUuiqVCizQzhS2kRsy3VLEbUXP14G4YdWTxywW3GEunVBShw1UrDOQ81jmhUn
4RUTFZfd2zRIwao8DuMJnOHoSA0Lw9h6Cllu76+1/XCom9M6GvRKg7nMOBkYPqLQ
pzijERTb5242CAWREJcFR4/Vx35SBfZ5FqlMebt6yqBecDOIkn3tqFL8AiJgfbY7
DCIqw5YvvYOt444xRL1t0Oes2bmuqxqk3AKiqSK0emeppNy+on22NBhVUCG0Jnnn
fm2bKVV9O7eMY4CmZhIpVXsEi5GN/Tcy9OZNBzb+rZR/3yRDIpw2XHok+uxJpj/Z
yg9kTU/OooutB3JqLyx+RtHAbh2Tbl9JaN2xNeBNbrVFspq244yphh8U7bpPwn9c
X6briHXILNj4C9LfHN9zvGmLfGdVInmIemWUaStumzOjGg5VeH3UZeBggmjMtiUf
5WPB2ZDCps2dHgwjFPGVQjMSUvDLNJXpynGCUF+GFjE8Sq9Ynk/+CavqBM//qhoi
4O6JCdqB+xLSePBvJF3coNcjsCXtRSaJchJK27UqKInybczsYZv0RldBAsHYRJ7V
EDFB1ESm46YWIIYXa5MnVdLb7CU+tLjWOwIG8o5h008=
`protect END_PROTECTED
