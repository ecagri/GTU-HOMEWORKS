`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ry2PSYdji5IatbRqQSMD4XJrAEv+8iQ/mpOkoPmi+NmV0t+7RxstDoU0hHj6nLWK
B+6t20t63Nx7lheU8ndjVomIucNWMx4Hzwuu5TjMqnpOGjoESJBopULx6O1BsgmQ
2frBLhGuwzNc4GoTklOkYIuGQ4qFWFV765jFQnUh85DIpjqp5+m9y1DNg1kap6/s
+4QQqMvZRb/TDU9DRLWM1JKX8Fk5NAJPegAe79nsW7+fLT1a2zZ5gJ/n248j9NsE
SO8JROgj83reYTsvxL/XjIf9zWNyI+heQIoOAMmRoD+xv33pVHBJDLkXwhhHxq0/
u9O96/5FnkFgxxFN+E4Yzt05lg9tvp+jmsEVMax08+rIM0j8B0QtcsBm3+FUb+lz
mLbGmz/W8Ft2ZQSzhuHmZ8+JmuwwRGK354pgbPVu6De0bY25yjfNnpL4PrfOVUhZ
BR7DiOJCt91H7uVgW1MTXl2sdhXL/sKPCrT6mLI0TzccIySOebKgzyMe6FBuCYqi
kZ3n76UQ82Y0ZxOksuKAu87KYybqei7yCh8/ysFbYfbDUvsYhJ9ck8sM7UxV9d3J
YK7Tn8hgZUhliGta3hdfQyGmaTg9OznckRqkZeFl7XO+dvrOvExDj08QGnc+3Ivn
p0xo1eD4n39Ykit3H7PKwHC+2f3c4kgrVs3+Q31jo82WRuYvQfFwjnkhbePYTIMW
kXixkEOLoSF8p/qrA9/s+RRCARSN0FClDBm4yf765ydXUxpdR8EhmSA/5Aly2eOl
T6zJu1Pd3bgKhLah5jT9+iB3CCnSsjY74EGgGvzeytIzQhfjdOOAuqck6iZ1z3c0
lV7vZslEqZk63W+3HNkMV6dyVRUKq0Ni8t7EeIOad+gS319ir5g9jH2CcbSiu2Vy
R2VbuY9ihWKT426BpnR7i72qqJ8h+ZwBRAGOQee45hW+uAIZ0S3dK9VTbRl2e2fd
ND/ApBrMvMAdL+BGJnVLjS3XGPWY/U/oNyRSx4f7LDAWsU6v3uRJyQEO2pUFzfRf
uCkESr2PMQSTNm4Ki4bIXYDtO0jMztYZtrSiOSRMXbv9jk3lAFUYXhB2XeQmmtNq
NGuDPlfrq6hIFD1cBv0eEZRmjh+5SD9Pg58gho7xeHAg5RvSJBEGQKkr4CftI0l1
DoAUGD0H3GMco9LQXyY9hHBDQNOMhJ6zTH7E7IUiJaJWe8uJ5/aOxVZl4+O/0b/M
/cd7cqvJUyPs6cEAKo52SGqdO2T96MbA1xdPHoUvhxDF9EUNK6lIDnjtiHI2x9Q0
/Dsx/DY6QY39ieHSslqUE6q50u8hbNn9UcOPuRABvxFpE6bfxKKVUUPCFcgDFZHx
JyVHC2tj727MKFvVd1yBL2EWeZ/M/DnfjL7cj33OOXnKz2V2kXA6aUDi4fNIxxsX
DTKr2Pn5ZKu6/N5dHZHCMiBKvcfk9mOfhWx45G6oRVYZqiIeEYM6jZPW5BvxM+9H
V5lW8JL+dM0Ok3lH9NLJ6SgJI1LO+MPeEmi1qPPlcasYnb0nPJYYSFPL76rdWZMZ
sMzrv3Qcr9Xp4628LRG3rkSJl1o9CIIUC11RBYVcHSWDFChH90Z9Mhb54uZlEnO7
LVseWaXkfeEetypQmskonHpQDVVc2ZYfmYGJseYeNCFLOS0jsMnx9vpw7T5HzU4Y
5jVRa4CINy4CyXivH65qNY76C87EbvyutO+t9SyVL6pIsftR09q3y9uSxyDqH1z9
l1W6kUtpciwfoGWptSV1Tdsg1yhnqhvmNaBFrdQsl7dZ5vxrH1pCUSJPmvUZH+Po
h/64s5bHOwDMGsZhrmCElWGtIOLEkfVVTs632SfkQMZTrY718HxfokDWk2oLu706
xyrEG5ZKTplfzDvFHfGpwupotzdpxeb3BL33r4JfIrAh0tZottgbN1TFw2/aRcvC
0N++HMOT0GXSIkamNNgYodkiftzAKDzS6guTgNGCe8IWr11Sd6EhoO2UoCKe9/is
rAz7iE4Z95LSICO/uNecQChCVHKhfLeh4twlFm9tUJsGlFqDpKE3a9tuKuuuePY9
fFksSvzFzOtjVyf0TSzi3tBk4WQdtsctSrgKK2LYQbpQqSXC378FM7npF3lBIhKH
ipVmqKpSRuKtf4wS7580Q3lrCTMAK2pyBD5RiRC0xFMReq6Moik6nj5Sr/x7pXZf
F2r83aq+Aa3iCPHtcNxQ1lHahsK2JuTbyfGN3vh0+kuWsF/W++UCq4HYaPx+cUfI
TOze0KP9IPb/x1VUJ3s3x0gMgHYVH9vhRDyRqGtNGjBv4oAc7hfTFNDX/rhPddbY
ErdMyrUukyzvVGxKsKUmCCMhF0T0aReQ0JRnXG7Wnsv+zXW9X89bHp0lyI2tWtMt
iGmkG9+z0NbvsS1m0fql2D3g+ZknVNXdHate6tdoDs2V/m3WAjkthkOaqwq5UJim
T0ly54VdEPtZkPMdYGCsRwukBkcByd5awr+Zc8pYUMnYxlRZt+5gNKf97RhAmzgX
3taLXvwWCSWku3Pa3l4IS0pvMwdyHOC9tVvazJoSAvGgJC6OW0sai2ZqUnuik93i
/GF1fQMem+30ZkGodZ4LL/hZK/Uzr229k7X83vdYNM3/8yrbUakCg4jrf+aHxW6L
gUOyaNpJptDUBZKNjoZ6+wOGAiJn3ww5Ft7f0VTmPUN3FRcM5jRlINkXv/aReNML
8oOxzTJjKw0Y2Nc10JSohrFx5yNK470EbfCblzDn+FVhh/NxigtoWK1nGU3oX+Wo
0zlaGiV/Yq6oABdALqMWUOptgXrS4Y9lBtbkZsMb4hn9Kx0CVkepe2dUEjY2cIv+
7je0FCsxcgOPlI9p7KtbVG4NiyytKovAdmA8HmJd31UeCJvHxHvlmSzuEeaG7pF9
Ixvmp5k6EVg4IrpZrC2qTe7AKmAqaZlpj8Fl72YgyrwvwFaNf6nWG0X2pcaa7j3F
Tmu8u5X7Tz0p1OmeyD8Dj+aLcngNve3Jh+u14glO0ErvDm8TDBcEZoNMHwrO0VGJ
sHYdt8WXluRwaHevhoIuyAbxEDfJ4ZMB0jDJ9AIKowWquPNT0gHQ32sQhLpsk5TR
jpJVHGEfg6axh8iq/wfv+pGOva3gIeGfyVvppnl1rYCSMH4zmO2R92gH2NLDRgvh
t/N+nCbxtOjT55ST5a0bgq4axR2vpS2+AZEAPNGKSZ1dTbcUj2u/H57pKBI+xrVw
JI666YWwf+KWImqdCTzPyDEPTej5iOTxbVn3HwUPAAxbW4nWnW9KuJCCWk/AOHew
r1xV2nv/uaTprqZ0ivlqpbXPoq3J+nQmZqUQvbmWxQP0QmZ6nmYxCfI6PTvCTWdR
IfmmB9AaEHhgYPrEnvZTf7LlCRhLyEelTaRPa7AfXnNOwZI7bKdG1U8aZFAW/qRr
OvxJFxIMFKReFWALrFdtouXEoO2vq7KP+q+fLdIOiNW3GQ8tiXheBKcxfU5qh37x
7ivhkR5xzt+0Wvbir0MEw5utrDIK7iJ5xMijcOHgv2v6U1y/7VwBKRAIzxZ9RZeY
TP9Qehe+9yQ2WdQSGKRfYF0g+vE5yXaXwH/pqDUtio2aaKS9fJwY5G6VZUDuqUzC
eJz0WhIkh4/iZSMy5VhBtKtGNsPdmBzmuRCTCWzZOW69U1k1zeis6XMivRWOGx9v
p4A7ds3zzEG0UsjSvKGNJ/yvvsXzYAMoWXTDhWZK41xIdUDM5vzcNCa/dACljRgZ
VZBwcjZdrkIERUGw+kg+9VywkdLoc7Sq+J7NexCZ7sEYBokCglG4VITt/GX/ZnFY
cb1hweEJhT0YjUXi2Zldyg==
`protect END_PROTECTED
