`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b+eCBSVbY34dodVi0socbCA+knZiYQFfPJ29RqUX7G3BL6m5qf5X7l2wFLAGXpoY
987j85UFpWVQx2u8tcSkc5gKTeumdhNJCqnTYkP0D0Rki9T3q3exh4jWCJxRe5e3
LNW+LsTMFBH1ol5Md1N85sqyl/9nMZ/VqXA1Th5r7vuxuxgGpvIUaGQcYhtTXq5c
hfq7x+WT9UrdhrtGOTc0P4T2VyGDybM+pUIb8hBFeXtIMRlo5xSAuGXSTz1ZJ14E
KgHg2XpoxsqImDHomUga2S7jXM2wbDDv4DQGiybMEGSG1fOWNU6pyIRyLW9UOZlD
0BcsQY/5VtCJ8xcsLBdNzoy6p2mpvI9aitkxdDDJCXj4ZA78XyMj5hw0yQ604aHc
19Y2nus5+gtgxEtd5eG3Tqp/H1XOJJrYDiDINwr3CyaosADcaXMk0Fud/ApPkpyK
vfndjBMmA9P9WbAY//+p8Dvfscyi+Z8wHvCRDExCMcU+fbmP+gVwVzOM2y0mtWaQ
qvzi0QX8bFDD/F+D/uZj9qUZ76bZBjx/dI90X/T8HmY1G6p1cnPywzoQ91qWkLLR
aXKQ3CF69vLIRMyZ8nxkRKEpMi6CV21jS29vwv8kmIDZBVh7UQHVfKBn4pBzc3C1
PeKLadTjVMRO6W4W10hKBbgwI6PWzzT+D1wGTh54kuulFA0IGlQLYR6IbKhvk/fl
4uMFZyUoiynjJE5bYVUAZAnCb/2ZbiNu/dbYNePF6pR698AwXNg7aeAcfn67OgHq
0lA/fNQfbVFtCvpIfHb4R5cwOnTvFJhqO9uPd7u2uLDFUwKPojJmc5wNiIJwqCn1
X/HCNRaYAU44ADpdykMr6h+PtoqntxZPfnnrmNJYPXawt8sS81bbzR7yx+X4LwIR
B77/et964u0CGpKPknnSTH4ZqGJKz3aImJzP+57y+6jLsnjtd9TRBdF6nadEFy+z
61DIJaPMD0tn60PZtADkcwpeuImdDlt+cpoCYp0Vl3NmKcNGoO1iRn2wfv8dXCuW
NXazF6Gjpfxh3juWyGyZH1s8gkmajV+3P5w3eeNycpbOaesCKAX3biikzsWbpR4m
/9qMFByeyLi7JR/LiuHNd4oR0pgShRkIfFRmNcqoR6dxheHphiSTG62wbzNDGsDS
D5sudLZBFN5fbcd3C5oa6wMegKDhyCu+pIKaNc3PA1VKadpDHi88vxcXveeaew+2
X2S30rqn1T8o0q8O5Sk8Vk3HMwYL195W5hc5A2FrgaxiBqyra/h+4l9LZCmw0dzf
lUJY+WBrjhTmzv4MnWuk6P50wxn59IG5ve74eIwVsUHwNM3e9Aowjfei4WzPrO0e
h24zQySBgrPvEOJ3x9qVBy2mKPtoHJ13DdUB5UFYstbW+vjz+2U5ELJlEMBJWg+K
0IQ+8+L4a1Q8ZyWRMJ1Ud8pT6x1ut4ie/kU20cWJuLNXXXasGe9E61Yu9GwrXOdy
Jt7XHB0BYqNh7f1agt8hLGaE7JNtPvu0pHPav6Gak+TlE0YkZFa2AIYYrnTWnzex
QIdcSsIAZeNZ81uiwqnXciMkSpuuMyvtzfazflsC7QzqLuguT7sKEAyJ36Yger1O
Svp2D8/KExwIUe8Mrjvh6MZTw75rfOoDOxCNoPZB3is/pz256ZShnqPRFQ+pDph2
r9FpoQl6q9afiyPUrq+scUxw5lnLe6DZDz04qdJeesNU+uB8JjptDrPYm09WFnsK
ogseQOZOpLggwo8NZTuiajYZFb7sGQYpdBvuM6tKksPPg6r21jHHOdN4PtpmoB1J
VyuVWaN/2QIY9pN+cakqXfg8tivNWeNo6leeEEZ5XowyNdzILKivpuDpR4GynDBB
xs9/WiL0OSRslNK3THupZksxIrLm+jfFGJdKmtmssULcY5KLwp7weZ05fzQt7JB2
kIc11T5ig4MQoJwgrN13U4YvEuf4zs1RiNkdmKXmzVat1RhtA+c039KPBBNYsi4z
9ENyn7ii31/kNHiwKwAq2nZ7ZHiimj0d6bWk6YJFcejGtPX2gYzWy45Tl/Q+ZqoV
KjG+PwAiDh84fvmr7/XC+v1O+D3HLycwrDEJ35U42/hQQDNlzQpiX47hULC/8oyb
KUwehjt7Pxb2Q++eyL6sRffe4Kc5g1nF/cCfacOgQ0ckf5OhUuiwFpcRsZQESa0f
8zAtnnznVqmLnLhaORMW0/ddhzGTT6vsrCVO/fCkNObBtFcoQRxDqfuhH4qD7v/j
UPi0un5ibzMIz80uJw8C0qdPs325gWgeeV+kVolOwOWYT+eZVeivKKuFglWWjITQ
aty0laNO84QBcs9rirVwhJ5fIx56KkEEg39f+h/IGFuODoutQUXfO6HeS7KKc9m0
M1rHtRrSJG4O/zFZ/8h8gkqgI3E/4LZXY2PwHeyrnfA8SNNreRxL/wIYTsZij6GW
ACGtcKmpEi4nFIIuRPfVkrEhBI0s8Tnqj0h03OEOHxhZixL7lg5EqHLLLhkCMqzM
5ikZG0R06Z6Z6zeAiAB/Z0vYHdMEFJvUkoQkrA/WJZbs97gOYWtLRMiAl4be1XfD
2qfaBv+ptlj+YXzP3Gpv/dPwR0Natn2PtK6i6dI/aYBh7O+++ZpXoP8qgASvb/9a
S1L/RtrDStYaV5gvyV7kVJGohZ1uL3iT0J3rnyRvwco=
`protect END_PROTECTED
