`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KNWSAK+OiuLzhGtIH5J74Wi8JHDJ+UnZU/wG5JE2k9PjXzYYorV/e5b1udxs8V3s
8xtsx4XIx4ve5yYwoelMdsK7dZns/UC0/+8+Eyupeic0gpUYyP05Aj7hXsA30baC
/CcqB+/YulDsI8i+IQpjNBgtCXeUtzlSCtkK1CMliE1BAb0BDyXo79+RH0Wl7k5A
AN5oiPtqbuEXtraEQeqonply+6K85dfYtlUoahZrIYW4yQ6HnQqvL8qyb7ZyWkFw
ZAMG4Wk72pDVIowLDx9GGlaC/ZmTTpmmGDfMIjUHS8QyWz+w5FO5+hHJiV1Bd6Z4
R2bkVEnMXTD4/3kMaqV3YF/n10Bp2pcK+29YgaGuQ567y51BxRIiMB6/Z3qMxHK/
0pYpqXbp5WoRQnBDTCXqLElLZODrmO8mBMyVkhg4kX4N0KbjigiC5PAygkjVNfZp
vGGGr46bG9ksidsTOi2wEc2H9xWBVTDAOsqeh2/m0e2fexB6n7X48/Iw5vqGKaVU
U+T/qCNtHny+w+Wda0lBFh7RBwbiWm/y5fVR5wFqNK/K8j0p7zg4jbwzfyD8cM+G
/3XrhyT7kENPezZBiCJXsIrouEBpqcLlSX5ZykqAst23lZROSSF72XSoJrUd0KKU
N6hZw3jwpAaPi1d4kgFVnP+6Pf6n+rsmBZN2VEOpd1yBOhjz1/LGSmmUiTzdZcHZ
5Oc0MlMn7pbB4A23TuYEwta/xnaI8Tobo3n2JVQv4U4AVt3skOiNMP3NyIm0u/Rp
LnoXv0ZZL3S9HQ5ROFlwD9NG8Kbs6LV9cCnQzgBzK00+tv/sStAt0Qy0eThF/ybg
GrLSl84GILdZXA9bFe5bMrsRvT5m+lUoyozQekon/q0MaWdv1lCTk8D7EMvHnsYv
26J0+dqOKZZaqqh5igBQaST9XEh5qdONtHKvqAwtgT3euFP/l0kAzN6U40Hp12D1
zyqwBGi99AGIXqbnSYkskMxenQNAO74qKAHxmxoaTbUokr0rTuPP4Qmcb8MF/jj9
in0ZtJt4TEs3miCg0J36/gAdxfftyhvPgZY3PgNdcPF0e+51L3rJsrmk8qyunurc
DBje8m7Rqcl1/aqGwUgHnCiI9VLX4l0LBC0VQUW300VnRcLRBqLhw8Rm0nGqXvJL
qiNhxYKXqtVXyU3HmjNLs8k/UmogYgJO4tNb+PDzbouKX5rVDotP5e7qFB/vdWqN
hRdenYdTwNz61lQf7+T1eBYMJW/+GRJIhiW2uhyD0XzIwY66gXL2F5ZC1SNm7zgt
IxXPkTI8uUnDO9yL9cw/DQbKBns6AyYmmEe0cOPhfqIQdAzF6OeH2sa5pn5SlCC/
ndWszdpbCSaqLT9F8DNM56Tpd1QoxkSRChLAXy/3wSFXJ65ntTtmaZP592NfyGv0
3TgSl9R2qU1HsaGJ/zZjhf3LGpwcuX+eOrkkaGi7Vt1jbPfEcBD8iwoUWQ/mv99J
KFDT5RSsecWAT0YgIEOq5qDcHURsmjZimacqCVGn7Cz+Ivzrzwqo6p1KqHErkcIi
noOZrP9ZFImqJ0RyyIilAK86DcjDaXnEKoICUtn3d+gKkedRbdPGLjeljDV5ufPj
GYErgLmj3moBqQMva1xxEhh/n8sf8E/GNLN0cQ7ggnAB2GU5oSmqolfejs3hgzSP
xTxEkSXxViF8QE0xxiutdEdAzLWSoe5GnUqTYb1jjnLcrX6o3X8nDO/arx0BXaqI
mP8cxlkyS/VBdu7lzGXnJQV8NQxBk1kHTs01CM4vptud8+VWQx2JRVW1CcaJcSIh
i8ID+PToafq9FE+047u6YH+YuyQI/jy7hbrwauaFg8WzLVeYk1gcUZhdVihKMxqA
iThi5OZJWNWC/BQ35y4pWOan8+PgllUcNkG6SbHQoTfADW+uSE65g81GPfCkuC/R
u7QxW6qz5WASVZlIQ+zGBEgQ/qj8m73hTCpNvEwiRoCIAvZxRWuwfdQZbjHxKy0H
96a6Qv1Uh8QvzsSP5Womc/A7FOCmkCulJDklaFWwoxxZ/qWKBjuBx9MsYaj/avOH
F1E9E1liRCKbA3B3aCFzahbyNfHLq2Nd0CHVhmvI0dKEJNWIn4szbSl0robRO4SF
5s+VZ1VhH1bK2mJvBRsZ0cdVJ2hnIN4cqfo1vgbZvB0JGWyfyHegjIB7h4IBq64E
kCIQd0/QBbcrfOoBnbwuCbTbMTtBoaG7Y8zK7XMymLzGAOMOey9E7Ojc6W3Z+Z9b
yk2IPGuVQjdrK6L+8WOSdmFAsJD6XpGm9GxD26oqgNAFShtXP9vUJNCxZ6pIeHJ5
GDwk109y1Y4fiDqwMixtGp7LGiLDjiPVOrS/799EGbft6eJpxKZ0/crj51ykJwUg
55msDWTivrIixJlL6+j1RMYWvNYMhBgCUhHQNvdlklEOutl95yMf61Jgg3OfY2Nk
HUwZRgtkM1vMzeQjjJnPNZ+/Gd69ahGpBQTRuZ30KppPSGup9L3PKi7Y8LowffFs
tm1PU6lePiTKWcHaylfz23tH93qbRCRk7QgTIBacG6HA4qMMf7wTLA/QWUHUJmhe
Kd3bNrejuAs7AE7Qtd8274HXa7Lpk46RyVZBA/kcyp01InOrZKYTmzJtP10sKdkz
kRmCIjuTlbfo7/YqpvYIYvlp7I0vDlzRW8jOIlknqdR2UZVQ0Rs2e6gERHnyeW2S
HwSEwo8/LdlTopPceF1+ftf1Gmdje5dJvh5SDlyILd/dTqr+YaVfyi6uQWVLHxPv
wrRK0RSl+pjXv0dpB8OiXN/ZPEwzQYlhF8IdM728exx84wlVU2K5o3OAjoxsmj76
qC3bJH/w4k+GqGwWgYABXCXjzVRv5FAFChqfQf2oiZ1nFz9rp//pBZEybFMMNvR1
qON4TV5IdlUYSMt6NIm5sqz9jExTarY6RZvqMOa32cPFrViff2+9v4B6AgsCHgd0
sLcRS0s6QspH2LTzDYb+Wc3BUKNQvtAGaClOiMRBpbAlzv0KpRH3SEkN3T7eEXWN
Bu1vzaX/9kB8/9yITWFfwwpjmuQDfkxewLmvbRUUrTBOdu2lg8OIoE7047V0uzyg
ITMykrUxwsixCUNKramynLrkL86LGuDZJC/OcGWw73npyMwGGnMsSScFf4W7sTsi
PWv42Zr/vsCPh6vBXckrlF8REbQQAsxzBMYhrjYIvcugDEzIlzR3J5iDY70FOhjr
KTgNE6azdEJ5L9JAV3cpn6cqVaPQ9IGnOW30fgk0k1HcX6mgLAKNEE/fxtmjxSzM
0S7n4LwFJEqSamoH3f6Utwmby/ZLIJzPTu0hOEEbwmjQqrKR5hSsoigdrjiGhXpK
YELJjiwy/FQF4wtEUmS+SWmqU9zGCtrzjJXMEt881dN7vZs3yFvPXRFkviYtEIbb
LoDPeJcONL3b+2usuN2ZM7QrIh8IyC0O9Mmwj1/36IuI7F7gRkd4bp5TqyGhUEyP
`protect END_PROTECTED
