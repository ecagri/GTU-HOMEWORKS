`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oRmGygVEFTHrCRKx5bN/9UK5D/dbTbKQqptNoYagD228ln2+OU9rWQIiFa1Oep1K
OhWVOJSWvM32oHQSZ2ZKgERfmwWpYeWNPqWyV0OAbgX8MWrCNgwWBp106RZdipql
Uad09q2+OORV+jbCsrwHmzqC5j7+x6mO1JI7VMVpl5r2H0mCO7kf3gliO+xszJ+a
lolorkcHja7FJRJy2sSD8SmoQv8URIFJtxEzn83OJMrMrLG2Ejk2m8tGUMtWm6J9
R6zp5GD/nuJGW/ITs4ZzWwt5jIog47L1eSEzR4vQKnX8758Wh98BiJhD/mgOiTNe
Me2pk3hrqgguKsXOojQSivqzHj0GhkkQ9A+Q3WyFyFI1YLuIg5QCrchjgFUBsW6Q
dg2Vsgb0/8wbZyCf5husVXhiuNVM10BgnOoFk9A3l50+MNT2FyXNmlhcBzN6ZhZ8
nS9Tzw5aS9EKmCTdzrDZN3VfuBMcKJxmXKKTqZhesKUwdfqmTHMd9vj/bGnMCzXd
lBLu31j1273E15edqngl44c+HwK8znV0DMJgIACqQ/GZM8OfB3gOPxEtR4Xau0Ec
RcIUSE4fh+T9dyYESJvBxtaafAmnoI+94iZ0J6tsPXERKIJGtdXkUvrEBW/nkiI0
EMGJRc7V2ufEPXpA/sVmRV3YYjdisydny9mKXpGbTEFCGJD/vXmMPOIHgnUIniek
o53cM7ExrXQwE8ll5amlK5yOcvLsSJ97Vnl4MoYg6IU=
`protect END_PROTECTED
