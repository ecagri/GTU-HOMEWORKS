`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4fvmCvhLMHyG6385UmPfxC76tZBfHrQzwK1zuK4jPLOE4R0aD6SYKHbcT2So1y8W
TqTKWvH0spBQrA82jKPCBfqiOXqaL9+VEBJuoTa0Et2KFEbHPcdR6LVvmimO1a9t
bcaXRa7OV50X/dgE2dxa3q4XTY58jKToUfSD0V7yutt6igdGJrVsvlVNVtJFOWXl
/CWNcL4AjMFpMFo9yaMNq8wBwS/imMh7PfwLJvyuLFyIC2LoykX9QgrhfTfkGYtn
TVdib3h5RltAq+CjYU7bszslcCb3yiXAmJTAvKvakbIKhfoyyDBO4inKBxc0TZlo
u3bkrvDXJEdOuj7+aLobBDb4OaLU81hT+sNwYVuTJxvtvLpFjyCz72Yb7dr7OId+
UzaHLlqOi7G9jd91r5++8FH3/+Z9RvXeFB/ns2iE0W8jmg+w5Yjz/MbBbrbT3LUe
a+bMMXOHXDVUDo6GM8YXUNjVTVwPyrq8RAbE/0Qgs43AI/s7/Y4by2aTbS4B1lg6
/RTGoHMtNYmmwqj8IxMJbbSYsP1rL8BeMW34Y+yI3Pnc+u4QyU+JuFahZhsrisqH
TqRt9g84swgpAdXwyRRTtGzHrp5gmgkyrD8OzjMM1ExVx0PTdR94wx617uGMp0eR
IjNMGMNjlvvBWKzG2eK9B07YMRR9q0bUeZL/4Ph+utVAn062SfdBZ54tDrYMxgJv
JGEY2M1ga6JC/dy5pcYcTdNwhnq94Ai8ffIRDAxbnuF7pQm6gopZcz1XRBqv/V1C
rlAMFVImYAY2pmE/YYTlz43oDJ5vNzkn49udIStnAAsM0cOiRXuYWb2DyhC2VMqV
HTxvjOgJWdrNAk5I/8vjqoUjzHuojADpxZYUOXlUPqtD4+chDwKOikav/HYwpDBY
T+xf9XNmmHhDPs9+epghBh2KIPY3nHE0SMJD/dkD7dhr6JDsA+gWf12J82GpWgP2
JYpLZRB5ofwWix6f967Nd71lFQKH+QuTwzl4hWpPyaF6tX6eZULD8Fh3dm+ZZUHw
xjo1rIUe+53+nLpox95rZHNylB5RGZd7FvUtXKgvs6T+O9401rkEpTt5MzMm2yvk
If8r7/DM4y4sfKKZ2DqQrDCuzPM84LILFTlnTWycGavH1k3TqMHS/OuYAydvv7F/
z4wltQhjQ2Y6jmm6IL5R1wdVZ3ELRoBlhNR/7pJJob3lpgjohbgugYH4M2Ic2+RM
f5a0BGLBozbHra+E+s0DqZ1yw+zLdN/eTeRkKS/PHb21RiLyJmh+Ihlgq98rS1//
5TzgIqr9ZPXD1Q0lGGyz0wzIS2vxwn+dKUz5A4Yxdhst6hnZCEXr5hK2rt7/XSHV
7j2zbPSHysxYFbONG9gmRIE0vTTN0WZ96M2WfA3KoDk=
`protect END_PROTECTED
