`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4T+VNT1ng8NPO2cW+FKuXQVK6ZJegCrNz4Jy+6phql30OXMeSpzfhQRNWdWtp0v0
h25UWX7n3y+/qfUNhaxNY7wuj+T1XvSr/gOVVQy5KjYyVkrl+jhvFMACwqBF5WTV
++izcGkUs5p874pOSbDaVxKqIB2Kp8AkSyf1s6bJKQp4nGkKsjqfRPyEQutS3a6G
8K7NVcNcgpAGr8P/Fp4s3W7tb3VXeQ2yRDYCUP/osbNy8II2BCvTSHRSfG2MTNGq
pBtjIFmmjl/r2ez9j6dXPVu2wrUT5CIpP4Zq01H6Zj6Y8jpIVlIpY42prmUMsq+k
pXD5SnYqAwz+OdyCqKNalsipaFY39rvH97RtG9umoOdn8zPOX4DDBgzGpDfVxZ6X
rkTyAuTCWB4adOak4oSEXoO0V6jzOCv8HIPalPpyThWeDH1BJu7OR8dRA2YfkD0p
KhkLhqeXqS9TUw7umCDS+8EJ5IVehdSJGl2CyIx+O0aGIMhKY9WgwKjWkymB66x+
jjnkapJdXVnkcnwrXBLmxyHSmA+QlV0PPEcsw7wdE2UpL+ofewHpLBfF2g6XXKtg
QdGjvmftQoBlJsAP+/0fgKndrErxy5AD4aBul1A0Vz2+FbUS6DQJ4tRfRIZGGh+E
vw1Nm9KrM8wWvnVVTwPs9a4aE2G4Tu92Z90SUJ/43244C5chlQiFtvRa925dOJZs
MtzNUnopLJLeDc7qs5hPbU1L3bD3TZ4uFpQRc746jUxhYqm0zxFUI8Pbal2PbxGm
B9NdI0Y2HAwVx7F09p0W4sHqFuP0k4Vtq4XcSPhy4t+8g8L1NmLqjJWvKv5Fm1w5
NyHPClxgyExqpAKRQ72KrTZO2zcumdLs6QvAjGYlAOZq6yNjjWHNFTb2nzo7Z21l
fKrlKJjibRc35c+deWcKkCK7OdZcSeU7IRGRA2cbcBRTT/HxfgeVsGg7E12dxibV
q85Xh4eoo1fBdxZQRTHDxsmrOTSu5Lae35qQQ21qDc0PdYs9za3nZl2Pg7AxgdRK
/FS6QxJIxeNbrL+XNkStbRDkVkWA8MG7D59Ai5IfytRCOVUDnqsnpLtpkv0eeY9y
gjdqDAyrDG3nmpPdbWjGdxfgLT4kp5k5DngQlvtgXALZSS83gMf8DJM6YeyVZnjT
Jydi1HQjHJe1tm3UPsFd9Z1PC+POxruov0QMTKVR6MFTXdUVYShSEVpA4pjdW+Yy
axH1rYOaSoG+BMijXIYKJ+H+uf8SgezuI8SCabn8o6FcmVwS5vvXaVwgoDkLQPOO
SWXHFqhMLaqfU88Q8KII3edgiITG9hZzXGSCZYD9vBL+toAxhFxpNc8Dr2hAqViQ
7vlL+Qq+aknURiUqa7FaNiLmHWx8BrbGQj8F/UdK+DVAPAYoTVIMrecrWrIA51z0
2SRVrUZNJVaxqWBLHh7Fs9PAQy3Bj+kFnw/A5LB0es5vpOWZB5kDKN81Rlufprix
bnD+UAuIA3MKtzivYz14yyFfm72NerCxHw/d3fLuRN7gJvZc9OpDIxS2s29SKlXg
JxA3P6efSu6dJK0Cpujh5+VMn3oA54r5dazPHmZu497AagOyrvrYZbmX17XXS/od
fRNxoyVA8DwXL4R1e9KEj6qrRHkoBsMJgj8fYfaMFoziygddNE2gZrXiUmkToMTH
9bxWem7eEhs31BdyM/3bFajXuwK7L3kHEEDV9a+lU84lr0+mJNuQ7/RjY67tllNO
7Nwl/bZmQmgjxrA+wDabE2O6fdpFuKjkZLogoVfL+Idn9j/rt0S5jegzTprMBkGE
aZJUbKSeiyDHPZFj5abMOmBwLlAecVbP0GcPfgA+8sic6EynNUZJYcjGiddOJg/j
emtCHrRwjAqdkdFlNxI8MTv+WcwfFwruel1U2IPhln2i1J1Aog77ISCLrUye4cni
ghf6Hgq2ylsRNMGbgM+4Ui+pqAWWb3n+DQHNX1y74G/MGw6A10p9/NjdkUeqN6wZ
6iYNwtaVR5ORIs1ocH3mhY+/OZsZxUxLNYIunLOk3UHOcGEve5RTzcgjyjBPyrkc
VO9mm5f7QQK94+HUAK/fTgcrn+6ToIataxQ7zH4zZWh1w7daQt3be3CLvUmpYpxp
16NPuVMwg7en8zKrwGuuN8ofY6QSG1mJFh8qYnfI8SOoH6BjIQB3h1K80dENqkMD
de/zoOvvI+Vr3ZlQ74LGI+xRipxqcJQAd09OdfDluZlcMp59EJyQcqHzXLa26O/a
CTKOYsn9Fw2ljWrFuVAs0U5puNfgmduHcY6JooLSkyFXdtkW4fu4Ls5iFSPNcjTn
PaCh0NXwfGsWL1OGnH2Ab4xjdqpS12xIVxhfijekWNL4wrH3imMvrCripYu1GuAA
tSnf46rPopugXBtnF7xTVlIM7xprKjSiDi8UjvIVpeEyEShGl6jHM3FdhBVTKoBy
+YKse9pBvN48fg7vz/m+tIAVvInE0c4cBuEAe4E84yRs8oy2GuLxiM/t5wlCR65t
XiY38wnYUcYrD9q16XTFBzCYsCVDlke7Jj5liDPjOiNEl+BbySkH8JOhWOG1ezYg
psqpmMt3fR0bOEjGc+0WrcJamZ78vwtwK1+YPAz2GzvarSAM/SvR5uM4Wde8nPgF
olnLhivBGiReoFCtVJ0s+osPiSqMVWvgOZR7zP1kAtmVBt6kHhg/NApmGEQQg3Cu
UQSVXn0tIATCYY6upcs4imqf1iGpKGfDDGtxrUtYnBtzffGpcf6dn75U4tNATwlo
4Hgj+a/XBYDQY2lI0WNiRRutmiMLguI9e11KgsjOBKs2XQs6mG55DfHA5mSxdtlz
n5Kx/1wJKIiIcTzEocRfv2hAAYdC1d3/hEDiS1BTkSAizNSpMlrNrfIiU5XA8fAf
Rdn9RWEPYUWlJreEYtQgMkz+deAdpkN98WzwoIh7Knrw70FmcpH3OJetl0GSikYC
0Sm96GOPjOmCCTvagHTEMFx0FxsOfr9ZBzJXEHPpyR7OzuXp/81K5+polXLMFEMS
pAUI8XaiyITExgHGY/LFAdXf7CcEiQUS06LEwg8estcurrBPWLmLqNDoPqXF2Uhv
0rDRq+whZDSW+9MjuOX3ykGyz6uWnjXKc6v/hWQ9Pgt7xIa6kjWWjP/wcz1G0weJ
hAZ9z6rnA8LeihnlxVAhV6pqTl5900r0SR0LkII8KhoywSXbhEYyrWlyEbZBCELF
Ae1CaUpd8P/2QRz67l0/zDhTyIBTSxRn78h/reZMTxnwxFuaHIZk3ES0qrYkxQAg
6OMj4uhKEPgBpIy6DjeBsRSLhP1JcKyl9UIc83HfklWinla1iqXatvzw+4Ehdu9I
2vJxUFfxC9UUekqT+3rB37rsyMLzVFcntaBnroKunHNhJXL+kp3ulfZmbgYoL575
`protect END_PROTECTED
