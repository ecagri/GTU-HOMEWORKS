`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
scrzN3OnYYhREYmr1rp+y5EJ/4o1d8uEZBFXbUIl4wXIDBmNJEeKyK+goFPWdBwZ
+QPIbLa86ZnqM9eivO2XtvaPHpUo12/T/f8lKKrqxLBX+QaNKTAdCKsXfyuQp2Pm
de1TRsGNAoT7cvmiL9bINXvUmdIMaLnRsLMgiQUSdDLSb0DkiKCDrRZcoY+QE9Cn
jdjnfdCGfSfmFhGwl2PaRUnOgf69hevZr2rsFjAPs0K6dz2+yNy5w+jVVlLilkhp
93jeOFOy8kLNZ2+Pg8umA3uUO1Os7Rtr5BzqEby1pV4o0XXPZWptEt7CGRjLd8YR
emidurcVoM2U23pB4p3CG3er4++xh8u8ZXMGPVYKgcWZGUA1mIQ4LVctPv+0hja9
AAr++963B6mTumrMe2fznawVUZiZOS2Z3XR4dmshCoUVt0esx8bWHGtsDPhqcl1a
GPHEOmohLAYS3XX0cLmN79xwuDtV+GN0QmN79wvu2kMW6DH7CKTIBe4Q3dHV3yez
`protect END_PROTECTED
