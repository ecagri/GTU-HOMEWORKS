`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CEx5FnaOW3aTcfqqI+h+Ckrkc85vWbk1Do+FoScewA+WGxhXjcNNRP/fad4VQiAk
4qj7PKCBZQhWhw8H3RGQ2RF9dJs2mZQWhjQVNisvscRomwAu26HN1d47Ug8KFPoA
8Lfbhn5wMJbjzmni8F27ecNmkhq8ls/TBhLeaaU0dj9pOCtED2CFk/d399ZRTNlJ
im7WCI9yRTy5cEyZ6vrzSsTEmNREzHpHlVUxZmSZ0yDPMvaVUqYbJL9sA5xdHPUu
HUE6Msf+tiUonFp8oiRvBx4yRalIF42Wj1FVZObsHYRoX9BxCZ7dFMVfaRExK1yB
gLH5dq3kaBEosDt3zGLjvya5RxUCJ9rO/PVXold2I586MHnggCwqyhCY3aBYPyvI
uT1dE/0uHQJrzSDHtRD4v6vYCILpmFV232iu6MAVlRB6fU6U5KO4zydIcCTNpDrM
uNOSUb8MzC5KBug19u/ZdVRgQ4aPbypdMMG2TEuFpSsm2g1cbfO4TBok0Itimdx5
nw4XF6tveKwcN4gYKZ0pZuBHGYvYWkV03dvgumJuW7ILz5FKGw8phaCC+jDgJHqc
owfVO9+OwnNYolfkoXUYSJ0y6NR2FdoJh8HOse/SP86ByWp3oYV4OBvPJXdu8I4p
z2apksw+aKCJRauQmgsfh4CUEcfBzgVWGBmUsYc9LfgHPaiRTNwz9Er4rQmsMw5L
TnLmUa+fL8NNxkdfVOUuo/qYRyh7UVrgD1yTBXOVDCDzNzORbTeMTO1FETBsN1xz
Lywxn2CHTenbwKZ0HtMPNpLzJ4ozQq0xMV+wqUfDmCpcnXJI9kwL/fSfWHItR9eJ
P3NwXJZPVVqnF0OIJ9O/J3TChs0+H6y377rdvcemrPW4Zr2q0MZvx8XASHzZum7D
mJzPyR0T6Jd2qkc5JBXGudWQUKf0cfQZC7lqhPsH2rXWaUgnVqu8ZY6wcdy66A9L
tysu5ylbLXUuZhfSq46YGApFrMmRVPsYqAIG6zQ2Bf+XiCc2WhPFOFXRlZ+8ZvI2
kw73RHLfufgWzwaBs/T+ipRVsSk/u0V4WACOEfigJXYbiiGO5qKl9W/PNvZ0UAkA
+wFkDnrEsmlsdiu32hiQkrie427nwtigCcrZsR927HzgREJkw4IMO05hpFTY0D5h
LkMRziZiOe/nPwj+7sInxsbr/jKYq8tZtqQWScG5fokrgu2W3vPS154yS3zBEndf
xgkAsyms1MLL2l4Tni5kZdfoThyDJxiQxuia1WK3z72vp4opuKVAJzKhhgrp5uEQ
M6ssL3Emn8pDTfaAMv2+3YKeb/2p+DcwSwzvzJ7MByNVY8GKtKgyTRf/Ozf7J5yt
7WawbCvLyTbhoyiOo7PlbXapt9yCILc3arZ/YG7xwqnNB1b4ZuNw4Na4ShiZ+Jwz
dmznVRGszdfUqVQ5lYVf8GS+N5AvtGnQUpdx2xLt9Zq+18MQyf3ahvYFItnkEN2U
n9T33ikkg8RNdVS7DqkgX0KaX8OTzehGtOA0IXwPp70SrixPXBbbBgBxZLfgGcBy
rC9CYpRcpgOGom/t+rhErg==
`protect END_PROTECTED
