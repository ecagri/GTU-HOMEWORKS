`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MyC1A0yGVKJhbOX4AN9VrXR1zSK8txFTXZnAAqoRXscjkGFolpWgo7QDZptwQvf5
BXHOyeKb/E/jbxHl3aDq3T9P3V/t8DaKipKp905L/7QDdPupzfwjJJMGlm3BJyxW
XS94D4CBA/JvM5h2Gy0X6YbDZNSExMwkOd0Wyxqt+G4BfBo80Thc37IgpP1Xuhg3
4+jQFDyulmrcrjcgT7H2uSZuMnjiz3Wp4CtNlfxENt353ADMcij8hsHnAra8MmOd
gMO8HohHy44WoPVxYe61Zdcfoo7LinG1bg9qE9AuQNiUn7dJOIE3q9NRGe268IVw
UG1bXESCdhZRXRDSUu2ej/AAVZ7qTfoh9AWGmb8DFfxS6nE5NlKJQYGJcq2paCcH
3MudsSBq3yZPWuYxqyJ6Hd8gj8mRJH/1n+9jk0MPBB2o5NDe3l5ma0Vu1hNky/Js
dCgKQsIsldbhUfjRXlJvPGsZKMwU2w3Lcg7PFW04u4yldaHSlBjCnKIB1cVsdCxo
eaakjJMBHFsSnv9+gWbyf1nCirWLI07d08dgfZqxJTTio02tPZILOK+orzm9dO9W
eASApQD6GO17Df7/LJyNEo/blqWe5xQkOy/54n+uK9NJF4CMsogFhuEQvT1UZb+O
hd5lb/NB6zekt23E0q3smh7IGG9pMVxiOSehx9LoWNEKM2t7tway4ZCRmbGCoBNd
Y3jpAxkrDdQW8xDusNc0s7z6rKsiNv72JeuFKyBGjPRJda4Yf50USlPWZsaoC20k
IFkKQq2qRJcnLQpO9Lq6ZfFczMFKM45VNTNAI21/47c4ErObuwWii4Btl5339DIW
rUME6X+niLMcOgUr5LXNhm0dsEpKwQdirN6Fy04Q7HuJD9KSExX+7tdh7iHgb8DI
FEGnMaUY9Fl3NK06hG+0Rueb+qzaboFjG2NnS9QvCF2PBr2UVHqdQ29UvN/YGp9X
fG5ywiydjbjFTgLPiW4A8vH4MmPC5ogPfBayYfVq1Xd8J/JGS7u07oAFGGZk7TyE
s55wlPfixxmNUgXfHBzKY2epka8F74IPMHe4rfhUxo7GhgIFXJnBZA00Dp32tvcy
moIMpnawVyDWQigDBt2cW8SZmhOCeQb3NQX73xpEsJ2LCajyVxyokCmke9TrDUho
OP1u5v47PSiO0qIt0P1Nao6lsYWn6XKYLd6oOjhtq3u4NKbkYWbTMwu+CK85cTBm
lvUeYjp2EO+/9vxvd+UEAcHc/OdAwDuejLXoOATSSQujTNBN9NqVHVY+3IuucQv6
7cIpO/zawa9hL5gls9xleSXbZLrXdRA6rPnfuNTPw8JOOhJdmuas0T2ns3vZtZO+
8+PHMGycJhJz4oTpvradYYhT7U8vAhzZFUT1dMuBEHoFlnzt+9hgHjD49hzIX2xY
pL1YrJgF0M7BAf2DecgX1g==
`protect END_PROTECTED
