`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kPvzRwIqrmXYvfpAwTA+cLd6dnKjCzaU86AMVsRj3CImKCA+u5MawKufPJKS2G5d
s5KPpQI7iUlPkF/c/eJRjkoRlQP0SSaa6BtqHPDS+95/Xly3/5w+1QMrWewqcVv7
ZmIyz07+hYIiHfZQvQa1CTFUkBAz/sW+1vM5NAmDrwO38Ap1WojBlZu+YGv13Nuv
/TZ3T3C1nkWXdyykPbNX+AVf+P4nauY7Silio/Nz5FFpaYHJYKjtpDCesMrtubWZ
QUxfZeYifQsZyz8ySTqyEOEcwByC9nN18514aWS+yzA1+h7qTWLxvYNxe+aIfW45
kY6WB0DytegEC4zV3p5E+1kdDsMORn/UbCDM4NsYN/6nidYbjR7nx84NbeXl5Li7
ThQoss0UJC1Mi95UTvseTWa8OmnDiZf9zYwBEKG6SdjZyyy3X5NWZ6B3Mug9wbwf
Girsbat+aMWiCJ2uXTVCzS08ZFENSxA71wfQnU3+E//VUgFUe4kvFm0mAW2xikXX
GBcu3q5BqZCtoTJ0uHrvBBsy2WQOWlM9o7UCZsoZlPbriwHRlnuPIcsxDBTfsi4D
7mgVI72LQyqho/PokRpN2iDZd3Sv4kimPUxOMNFe7ersLKh54gyRzyIgDO5juf9M
fmautsg7qNiPqrc1Wt+wIFJmXgximi3xIObuJ7NPKG6X8O76H/AcfU9f1rRwP9no
NihXTV6zm1+Enr2ub3RrqxWLrOFmaVnsofkjImhNvW/WP49RU07OYqyYF4/HJy0l
GeLKJuug4jAB+l9W2bvsxqAWgpd0JlcfjX4+MsT0oHnNy4Io2KGvJBwyS8mti+cp
eoL79KpPOPn7cFmnA0YCPdOZUkGyNZcM4BxYRCwyxrpnRmYfj9/Gn1lQtPq1eJye
`protect END_PROTECTED
