`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lGqSaTjybP6umzuq/+LvQnhqydw4h4uzt6daJdeIKXxcnv4+tOrlsLgbG6/7bnEC
f4/3RCFYXLDYP/OGuot/FXddLWv30z9iasWbSkHLozNQLdcwW6fzMMmCIXKG8DOF
P0m+Gdq3Vvlmb/pJdh/JDdUM+YQzsOHbVESbzYhhCuVQETy/TSnYyPq9py2OkVLB
kJuI/5Kv/rYP0xdM1U5qCXwS7llQ9F28eZ85AAIyfvk8sP37IHJbbHTTJXGhXQQs
+wY5eqZS+c869V4xW9WKJ/oi0p/jm6XFtmXqJyDBwYVznaO139MVTQbO4fXmHEpP
rbDLMsetmiDwZuWza9J7tCBIB0KlT1Y/fzWJGgpkXM8=
`protect END_PROTECTED
