`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1L28Iyai7svawBSDy0FyN5loHM5Kfq4+HUalTg2pNXe7+BjHsS8msZsea3CBVc5o
WCbUhvwPBvi1XcHJTKUPcRPYiDfPVB4/eDQZTCkXRfO6wTGM+PYyllCNVMDhwW49
xcVfzAV7mmvLUL3vX/zGPDCPvOVUiV7OSPNXj4mwSgcalz2jHvXmHV8M+u9XFVyu
fErjcR4dR2MJzCAYy6CoP9MaMjDBw8VsoZDCQuhTKPRHS2e1EVh9cXPhS+B4DZyo
M+oZLH/PHkvOuM20wPV4Pre937IfavmHMJR9OXRTKPT0KiHgvQBdhi73GVCqMYUT
K2XIxmAujI0xpakzxcCA8epb7udiRdcXkTvvy59Ve3VFMbiQGjV2beqmRvtJlroX
Ju5mT7Gc+x0wvUqF2kfoliPSrg4YofEpubdJfdJxdN1Om4bbnvQw0n0a0AJdG98g
Vs2iDN1jfZoMj6qlgWX1vgXNaRiNPZRpJEwQ4/AnAQdXwiGlB/rvga/BLhUaAt3w
uT9SMB572IdjIi18VwMG0nZ4p9laZNuBSq+bQ8hH3U0t90hYEtJn4wVyXmzTNT8u
bklchm9pMvmVNQRq5PCGOR1Pva94wIG89boQq8aVVVHeTg0y/KIIIwZcGNBfjsAU
YF5PXudLL4bdcgptok9LZ9/lvI6Y+X3SMHfStkHM70ictjaG/d7ZLAbqxy9NBpgC
IXwqROsFYS1weXRDA6H5knD23tCe5+3W4NEE4C3EcdjA1HjOaawzsthRILsApaJP
emM0LRPZ/bMpTACXsbjRctVVy3UJYWMBMprozehuvJiVBRzoetAMPny5ts2Q1V/d
r0LR2K5yI+YbcQDSZShVq+U8Uqul6uwXZ7Sd9XAPSnHvBfPEdC/VdowdtQCNUT3d
5mrBIIOUiBgxC8VGIufiSW6QLIuvJyxs75VSvTc/uoZD6knQGxoiUHM0R1DRKQwB
B9LJ3/xGxN+g/UlbTViVV9TATFyAt2f02UkpQuIwnnJ1DbMg84FbTwnP5EdX7V7Q
42VRsbrK1mpCEDO+CsEB+s8RxTAF8QF63IDf5OY8LZfj1372S5a55RnyK/ZfFVSx
OLrsvhIh8NXw/7WFmQted3/KpTs0CucmdSQmD0s5WGC5ETisqJjhsadA+la5TE9m
JULY1IUEZNLdp4mr8QW/1oZNxXBqRBT0ehYzBX7VnjL0ToRsUeb4i/SVb+9MyMrY
qjYwm2uQbA/UARKm9j4uKCM29FYwdlubZNUpx8s/8uunXddpQpUHPvXLCuOhZ8wV
fb5ucMXu8GEvfuu5YXI678rgwR9Q7Ay29ywLZlDoz63AKj7/3mUm/eW3/1rg3195
vOS+7DjxiwwDyB9UTp1mn/Z2GUuXhNiIDknObhG41z5tpqOt0U1fVLq+bvCU5/nv
9rG8v5qPSnfivVfW0oQCQIvutyNiD3q7NitQ58Af2bCJWcIYlPhW5R0nDzfWvfBh
Qr4IpuMHLoCu8Ir6xtgJavSNGB2lrRJUbyQzp9SUxWxXnhkSQmVfdbqkfK3LYE75
515FEYUSbs647GVuhiSyLSrbZjc1mQ6SSJ7SOCA99r802hF6XlslmhZJ1/sEQs4T
II3TGr8fXAnH4Sij/pICyEmF5lKkW4Qe4seTua0S7wGasIFrIW8g9OypWVTaEy3Q
nV0zE3r6ShH+c4UBM5V1pOzoXGaTCHtuUW8gsIkTeyk0fHZTCj7D4gmFY9uM3/Yb
0xi5pUUDcaXYAcafL5qKyQ==
`protect END_PROTECTED
