`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E9ovI9/irTP/Vse0TNgXYfaFXTNvbaznBTwlRHhSZzQsk5FR3S5CHaBPxCn/J/4U
txzpUwsPmzJMHr8LKJsOXu6MsIhf78llczZRmmHdFi9oWTSMdE+/aQtmnCog5UC5
WotBBfAz9Cr56cZYKbndgSLyoA2EjfLiklZribTYvaPgyNvsoY+q/RbKoz2Bn7L4
GfRFuwPOygzB0UJUDBYIzbTCNsQkRqCy5vZR0GNbhh80Yt2s5cpFEuWelMr3qy4z
zmp3x3QDilS+0+po3JONW4sFidniE8GM7oSreuWM3TnLMjLlyN5iimNGGUZQgA+7
+t6QII5JMaE0UJr9exxBUD06XHCppY4O3Yj4CfF14b46fQpP9xD7Fy7H9kPttapY
iC/DLCeFk15wnW1WWIHov4NBKWKndjxsMwU9FXpUvKyE3Dw0bJFfzYl5fhcOepA2
lkGY7zf23vaEOIA/YBTAhBoQR13BkdAAypAeC+KDCmtF5jAUFbrAvL38QTT+7Ccd
mJa1Tpe/Q8V9Dvbbhj8opDRbSgg5NtNA33zSGIZYFimrP1k2sEjozW5ncalaZNOO
/18uS+2LCEGxcCO7F67iZzsSfVPbUmzuBeyt/4CMChuzuv2yH6TgIIEq9MtllvTY
vu3mlN7CspOS8bp0NyfqeXxxINlZhvtJ5yNPsrGfhMEx9hYVriEVUzazB9xwOr9p
2cfQDTUiyEFK4NC8a18MJ4l2l7t651f0ZjmUBs4e4fiOxz7nezTpaGPonLB7Dll0
XQYcWuYsHhqZ2sOmj6Yv0ayexJnm7IjTBVNF/aOsNVcmqxeml7Oek/ow5+M9dLu1
nkgtBJxzqxoetAgTD8R4F+d/lRVbZ5dRuhjmQDBYhlpw77iRSNjuoZYdZxDdQi2j
wPdGQHiwBLyWtXoBlww+EDBZCYU7mfQeDY04urJWEJ9nePgUTF5o3j2zF9bdQj+Z
dWqbzL0qhAVj1irmWk1F9WpEJtxYXZc9XHpIVFVsCXiDOqMdEuZ9d1OaLBmDYY4q
YiTSKL0m0zU0ZHf+1pFdL54eGU3MQMMUhsBPjnL3WaXKQKehBO1JPDy55Nt2h3yo
Q8KdLwReFEP+Jfh9WI8gSswuki/VHylGPxnzB49HIikT1IBgdYZPWv/e6ku6WBSp
EC+j5jUVUCVDaYbPFWif8ON+EPXpz6dNbg4Jk33GVkEPu0DKpaDHi1s/kmsX0nJn
I0XtMpCkQBErmDDK58X8jXsy95Ady2jjVDdoZkXSo5jAigGTCb2tOpsfWI+2D0vn
JjYXdRFpq+Dxgwrmw+d0zXUFZTprdHIT2sE/YtBEHtNUtAslS183sC+6+DVYT/c1
R+Onf7Kcb1PKVq6FEqYGebNtVpntQQSB2Af3w6apj1L9u+bBunqNDk4QGLAXeHJ4
uAbGY3j5XuRHoc4d4pzNWhODLiMgwh2a1r+meUVNk1fQ/lDYTy6AxdtCOlSuQlKk
CQ/WVSQA7xcyRjQJnl5LQi0aMJHWy3vGXgoTD4MVc6mYJSXoPPg4pmQQqpuzR1Zu
uU0E0R3DGTeFPl3tWf3ZxdnKMw0B9IrT/0thMSzpPb2v7PStrGbDQbbSjWBizJ1O
XIhln8veMQXcVebuwOe46ZXV6N63UnhkhaOrcLG0B17MfP9y4r3S3i2XqEdvTLi+
ZHcFXpW56Drpjke3pBY0EybghoStKTxpSr50tnYDW2HkwhS5KLyM0einypY23LiU
oYrRgHzSamVmjKbg2JKeNCM69ReV3bt9EhoJ9qFyLMavMPLSA0i8eo+cQ/P6cgNC
zxkZYc0h5f/po+nM2EwFI5EXSjbXuEm3v1+AK8FvB0laZVdB5NYmXnYMZHL91AMc
BOI9Pw4Q6xLIQjl1P/VHI0szYwukGQUS0bE/O9P+aqnE5psd0qod5hg4/cHzRsO1
LzQxBmuu8/R6IjeL9NhADOVxJg8KmyBa7WhS0Hfz2QIQaQhKj1dvO7YnfOW/4ICU
7aUrhFWZf/zRWo1cXbiWe4ZCBhPhhBwu4HXmRbMYuWu0f8krXwjg2AI4PL4vlpKk
kRWSKpTUYYmUAZk8eO8F6b1fqVEcKdOeXOgKhjqWh3DtoZZKt4I/cUtnIYtzCFd3
xjvQQ9++068V+D5J2ZJ+SVpFwK1nrUpSO5XoMkvm+UzLoTF9jfSlK4KeEgAQyB8S
RPiV/rMBAsk8G0toplo97fsseetp62VJryOAsTMgoj87/5cZ03aS59LuXc+l7XB/
ofg/qA+yTcXxLQ32sEkx8J+V+YvIiX6eAkJEuD06KTGZAzGg0VQKBO8+n1hIvxKY
PGTh5hHqRPJx8yIPN+xBQMlnI+85jFnL3vyPE/0tJFVUymgX37YLozexwFyKTq8W
ioTnr1kieMyQH3zeEQzXOCJkoEqOouviEwNdZ7KNVSgc3LQDdOyJ8y2BDOdZxlYr
di26aT8EuFBzARyc4mD8yVFQj2Oht0ahlipUW7MAP3k3kAGdNreyDaCPQP9jiMW7
3eBlEpfNY9MjqINRTo0r4tS6hbsphHCZ5fF8T63Rkv4RSGThT0dja5pIziSq/iVX
OkJ77ursI1957LNLlrS7C8mCnFRns67AkjJlSch80/XDWxeM1eoQ0DKVRRLk3ah7
l8RPZqA+HzG1n4LMkKyBqjn9VJBk+ScPPC4MIO13NfekE5MF7BIBGVSYAaNhlUW4
TW8lgkSRfgI2V/yODrZRwLXUYmljSx19o1/KtQN62O2sYQhioT1HyyQtmUX+6K6G
phiJPn/WbuaAL2jN2/UxEDwNCuiXObPMJU0Sy978BjDcegjhvuzr8Ld2Evqwx2Jr
6Umnm7JiwQl9j1bs8PVrVCXHzunmQozScBUh6zhSwWK6bO6qPtenaswZO0u+gJnb
hNxJ8Drw/GOptdLi0PEoIV1Wsd++Z56BqMz2YiwluqAReI6BXDWAcLVe/HaGyTUH
vuaHZ7EXO0ld7CG1aANVq5pjN+/ZGH4GehmLENcuC1qNcL/803ZmIULyaIw9l770
SsCyLfjHSeOameeFMyenw3EEQbQR2mZvj9jjLiiKcn0iR/AOegENE1uFKrc/rd/y
EiW9de45p+QNqXbTO+sMceAMauS2Q1d6cAAgAWxTTE5DvjZewyCKtC3E/WCTPVri
RohzJd0t88K1NvsF4HYh/2nAlf9PJ2zlEeUFjz/ASblC15LtB88f5w9PKhR7wZi0
gyLNKtQy79rHA6iomlcxzQcDI+vm1Uh7saVP9I4ZStQBk42zFDFIgoS8X/lbcaxh
urzmAfKhM8U/xJDtPuW70QnJsIpJmteVneEmZJPMzpR+v3SkBzFGRhkgWAE5hWiM
EbV1v9Ea8igdMXnhNS1xfVLR0bkbCSFKImoXSpYyKNwEr/TAljEd8tJobTu5YU6C
+9F5yaGcEk3kkfbaWaSSi+7znSmr/TvJq6C+S+3y40vWR9LpYAtKljzEI1rZAYEN
`protect END_PROTECTED
