`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aDTqpzrU7p+wambnzaMBWd6Zf1v9S0VwYdAM0zmwAjRQI5hHP9YsrQkddvyYd9SS
krVXI6jNgQWF7DPEiPdRX0X/GKlIukBqQID3jtNgAL274LVk+oJHoq31gCEZx1rt
rBncxABD81lNrvJ2nbIVejQvv9DRXsyY7ahLxuAmEjnwEtAkQ3kpbizD3YFJDdIg
kmCNTBEvV9djdUvRNg6bAV89sxIqdGlrO9bCjAqOui0325QsjyAD7nri7pWDO+Ue
9JVB01HAsmeLKA/Xn4A/juBYcqFy2Luj62oi051RwB3Y6uEeTQRsj53eY3Nn6CKa
GXT54inW83q/eup+jNUFIgGeipIMok2We7/s3+wI7dvKdLaAm3r8/ZsKVIYcSFWz
gdas1V43sIXWrkPhRRk/wZCpCP2eRFsHiuJgCiL6S2Ih3tZo55/f0lofSdC4C3jj
IBvTAEVDMTY6MWOYxCVbrK+SI8K1B3CBTKvYTtLU84MxROIRkyk0STFRGvg8dcLK
yYJfkfJTe8qA7IsoXUYbMXoG9/Uflwh5e1Bm0Ex4l8gbPMGc4XWDwNTAMBium7jl
4RkaPUHn3A6Dbnxkh3yn/5w6CRsPAviz1oKTCiaDktNY3aB12U/2IZhGRcBcBn0E
FwQ00FA87FaD4Q/4WxOIe1lVjt9BOBbM+OD3rm8LeBn6EoN+lsO8U+A3BFOaWKi5
jLf+TxrbR2UvBXdcDiOG0LrvoVly5uKf3FvprDh0YQjx+yvtHqv9LmBbZhUDfl1k
UW18zn5Nwyijkgzh3MeAr29MVAKMNZr2lEVJcQZ16GLdbqP4/aCL4rCxmh2XNPe4
qVcV7ehddRmhkCQYQ4hiekDq4wPrCv8uqfVqO8eG6eXCjYWfCQa1d2EKGuIlaeGG
ICw3CtsEs/H3JIbFdeR/IMmbCh8e9XQSqG4uW74V1xxa+8DMyCamr1wqUpE69bsz
8F/oezk+EB0ZCruKioFufeaWiU8E0Q8NaDzS81LpV1U3FxCZW5eGNmqojZKUFO6r
T7vNgedDZ3BKQ1Ky1BLWTEt+C1hETvByKKKXt7/1dVLOJXzad6/moYh+dmbtkUyu
djzhpD/1v50PwSrNMEhCBYAMIWyADeHV/NtF9o65J7+B5zVow3XysH1gQYqu8FdE
W9xPDi2SP8Q+A5AGy4pqt3ld4BPsNo56TanSgpV4fHyW0Q0guyGRCLNfv8dYdwg2
CuaWfGW8d6SKLMFOItl+zTHhh/YKWbBDUDMkhw2gDrYC9YoqGzsxVXk6bP2JS7fK
QR4svVIxx4/4FAI9lZSLD+mCNS3nO7iWH2esrDC1u1V2eCKImkTfUKnHziLGuIsE
mFHbiUomT0vq1WSDTCg8bGb4Ora2O1ikv771iXQ7MvKbPiO8/xLvvvGdtZ58LBKV
On8eu0ahWdgzeE9Qj/hqVt8n+/jdUuXy4g7AoWHVv2zcuee8b5s/McFYQA99vGW3
UUgKQ3/+aY3pzn7u5j6aZmUJE0K8ok1q+6SfciN7W6XzbXDvxJGsg/JsVKcF8LFN
fbYjM/a3biW0YJ3GdFQ8MPBIegUz2Yclpy5ykvmIqZhrSd4VN6/OG8jeUp8HnFMW
M0OlOJO88dyTIRKBQtcjU+jvzdF7eLpyxe5fQjIIGYVFBF6dqJuCUbdb73YIFXyg
sBVbhwvEpSQJ8dJ4oBfHm6+VlPVBUiWxpKaN4gl4SGAQ9RIgod13HV9C2CTYYWMO
eqL7o/p7dQbVVNhykUWg8wSHnu4j5pfYwFBdQh5XkZYoMVZRbN0O+42wEFVl/Ja+
YAnLmTYuaLpiSbgGCAEAQ/quMbb338rGYgagrqUhevXtClKmPP175Vdl3/pdMHJq
G2ucB1IMaZbvsIPO/wZ2WSvR8XF3rUi6GEgIJvLar+Axc9OvT92YSWBbqI410noI
i/qE8v2bM6xNLaxAxhEhXw2THtqqAzggx5W/FhLdheeskByJBHiJ4mlpXYgyEEuX
AUO4tr5clNVM/Y9N6NXuFOUx8xfFtvkm8XItB3AqirgvfAXwUrvmqQPtfOT5+eB5
N4Szv3Tj4lol3BPY8bpEt1MCP5UkTmVb7PevoD3jTzdhnrfaVevpM0dVqh3BS4V/
8IuSr/3MjUkRWm4TgKQn17fAKY+a9EKnn9zJDlXIPyY=
`protect END_PROTECTED
