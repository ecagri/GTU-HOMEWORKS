`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TrUbts5BdCkFizGYDgqVUdGan4wSXi+vfPfpI6d/9gWyP1F/MIcmIGPlup4RtzVk
Q4BNteNQyqNviADu6G5JCbRKRVUH2zVLxtt24mAZIJKOlgALiarmbh5f29qZfX6V
xpkGYyY6rGr3JYzPUPNJvYsoT9dnbtGgf44FX4ulAiRGyDmNwUodJtPktqoEWQPE
tdyQIDEc5282u5bq/OQmPu1NVCqezYFEFqvoZSuOXJuEMBwyonixcutabXKehAHP
hkkyC+9hfubwc+ZnM1hxsML742VM4qmqlqzgTWKQ8LU/VGqGjSRQq8kwYabWH28x
+vKKN4u+b4INpZyoYfZZaPQI6R92Y1ggFiWKBBbqiLS+EaUmQx1nOS1uXoACz5aK
GjlsaJM7EWBg1qSv6eEM2EFuTrhoXSptzdfkO3YaCPpQxjQ4kvvxqorJdOeWXPFh
NEy4OaQTOPhv9DiWPy51E0UPanUM9D4L9LN57WYciZC9c7vYR8O10PStp4ivNjHa
4g72ub5A1D/LfWqExra7e4ZyPnvletVbqZv83KIgmwQw5NlZbsYnkQQKubZe2OSg
PUI2TPWJVN3r9Ssn7xJ5j7qOepaHNgVA/1OQlV4B/XpUvjb//fy1Edtbqv9HXuP1
+hkJI3PHlKjqOJDCKEIDX4vfjRIGmh/M2pFs34v/+owzssUnpKvCOaayGB3VJnpd
9SUJC91GKYgm30uEUN/1ZOSM9nEhJeHCL727XjRew++MD2srnr2SVzQcIUFMbE8v
2QJfquovKG4e+PpMWQHO0vYWXi6VEfhMhSjmIS6nq9tvLQwA2wHqn5Gmc/PAufkc
HmmNxM0/yOx0prq5D2+GSsSTwppp+UxhECxgAfVPCeVbIVyl0PNFffJ1EZ1byRqe
WODis1D5L0O1Lo1Op+4K9tlNZHIJTPsZZ2wpaQVfe6mSKTgg2WlgGXR5LyXQ+/jB
8Sm0sf2HjJFyOSdDJ8OGfZbTzq23yXAIkm6CvWsRB+uiRzhKmVlPaVUmhzagi2jA
+htJK+7zcKRLLPThe7a8Yd1ZyAfkRKWf9gaqwYHo/zKN17Z/pDqm1gomUv2miFS+
BsEIK1OQPzfiPsu+5kHjDetnzpgQwVvuGDseZwLDTsrPzn+X8b5a+tIaXHPdy/SU
P0A5t06GWQohsy24Ynb0crcK9Hyl/MGn+sIQhDc+sB+jmkrPpnNuWtUcBng4yXs8
GMQ6Br+tTjfagnb28fYrt2rdKn9M4yQyyuh1d7JLcGH4mo9tANULHm+ZXWm0oj6P
1oYjASZ1lBX0CAoBai0n41Ykv4dF9gvEx5KY/yl96oP0bn0JmLmRwS2kg0GlsUNT
Elt0rk1uRdc5XxVBn2NdX0QhKH74o9vVCWq6c+wzzbiiqYHxPSh/Gw/wfUsmnPUY
m2ZspyffJFECGwZdKGxYkyQbXsJ7EJXM21peGIdYHGz0Pdp0IamHMe2ieBtx/XqN
5ALtbTCm+ZaCiCcztGEW86o4ZKkeicenugxxC801F+9BM0/AA7sm4OFeWi7r+QkI
9p1cKK7fB1VcJwlnyX1ZMajj99w7Yug7Q/QOVFZ3x1t29mv8zVEc3i5acqH/37rB
ZS0kf/zw4qWfi5j6vIDNLFYstkrPTr7C6YSLC14MlPxymlIkwnG8DMDgAA6Q2eOX
/87MOAnW2WwWZPWQduTIR+2Bof8SdhQvHV3pUlmn9dmhwlYAVlF76NY9WNHQNX6x
mevbpVLuJdL04e94Xg073Z54hwTWXilkDmglRv/6QJwEaYWkoJ0LbrNJbPDI+JfQ
mV5P2n2YBVeo3Jps5lq4IQbAEqBTGTy6repd40NTJfmAnti/nCMKytbaXPEYPwWM
cEMUAS0Eh7Qv1DD9FQvZ+IywoWcAp0WsTXFHi4ic+jh8Y5ccMsQjuM058grZkNwq
5sD5eYa1rGSVnymkkoGQ3IRNzq6QtyXX+Xt6ur99eLVXVXIlI4EzlaSZ1a94TRaP
6UG5EvjF1Fnl8BXkUpyvN2o4V9FslJKrBXfDaOC1l2RoXS/sQpJD7XhB6aYXTAWQ
Ogq4w4xaNTGCTY3y0GKOTY6i6toU0TcFcjNZmqg0WR4Y3YHrtCDKqsfEBCkP61n+
q4Q6wl+OEz2DZ/eANEBOMkiEk/9b7EbsZhM72TdErSMUPuaOTLLV4ka++uU7k8oK
6jmCtC20akBVSar8f1BgXMBHdpsz8JOXsaxVDLpIBS99bAMOdIW4PMjSJVum6qgi
U52mX2vDIa5hiIk0inhfPoveFfsSEZXVdy+o5fUNpO7EK+zcNBf56Hb36mOKkIF4
tdZrmZwyo4LvupKwdSKIPM2vr8+icoJ9FvsKGg1RGOsemJFHvZLSgysfV6/5WaFX
8VIB6/BWGlrgZK11W9138u+4Hf8BNoDm0PRhyB93ie+4gvBlrJYNWPeiuweKGsRe
/UkSAiOapBUipi95JcPJ3kYrS/2is+Q+ykDmcwJWuIOrn18ZXCQXkb/Smj+e9nY4
4lCJ+JVS6ehuBIjp/KGK8yw7reto4+fj6TkqBGMwrVSmRIQhuHG/7JYYKa+Kefsc
DprApBEyq2vDrFNXRROeFdTsnrZ3fzI37VNBsPUdCUtH5IWiWdiWQPm+zP2ktoSj
w+PDvbKZzS9MkPjoZp4+osAZ0gWVKQfnds6JggQsz23ojaqqRV0NNZIbEC8k0Rep
A6FQ9OyBLjlmVGzyr/4R0H4vPJFg6H8yMl/eMmoRXQa1qQz1gEYlM6ntJVMcmaP+
wiu1nLYUNqsFYDfjG6DMTpKopR0BJsO2rvxUJtwvuvLh7Lf+5eQKZwNCKkaUB+1o
rrm+tMMiCzFr1t7qpUC39AWDJ7zqnWv6NaxWb6v/OrzZcLMn59N4gCgMfI+drK0S
g4/qE9mSJzaQvPqds3D3PQ00TbQpWYuzRcNuWRI3dL+Aat4bZeOqz0xVfVnLrn/p
0OqBFbpdfXsTceyISb2GvaVv7G0kfpN1qt2XBubn3/+p2KrhKgbMCQ5H2RBiHIW4
lYC2zsanO7YtsaInT4qcfcNwYaVJbD77T97C1uLvbFdwyNjsmDx6fwJZWKLhJB0J
Sd8MDR1imG4yd+rcAzB0PMM3ksnk+7Q9aqUVBOb+5otQoUScSEK+oOG1bpJWur9Q
SXraVXcmS0IJbvmugV6FY13eCRf+0TfKP6wBRveOaKNpPpWQUR19hDtoaVepO1iN
+Kfvs+ruoX3iiwptvl6fVuT45nEQRpq4J9jKLHmOwBE9uf5bZYeSUKmV7NFjBQAY
o0kgof6e8VBpPFCW9gW3XgfWdRdRr+VyHoBUq9FO/MbuWkz1vvkEzpQvJmRX0epj
qy1OYUR+9O/R/thIWbUJzjfBtCWIE02Ip9PixCgJXeqnv77L8VNvKR+aRC+S2vBl
KCs+EB3J6r87ZzqQUQA6upsNlRSNutibPNRwXv+s/GcwPIa41Kl66FXeejOTkio8
sd9jW+puDqYEekpnVCLJKj+ROz5jcxxSMK6ZyBVTzxW69dDn0DXexMhxbR39sxWH
270xP4KumnaURUWCCK41csM1F5FHJ+Zpr18JhuH2aO+Bw03CCQPBtXAONsnFjC1D
63fLMsk+zw+00TGCsx1+3EoRTJM1ceJH9pKPYn3Uc6r6Qc4m6lv5IPuy8t8tlA52
vzQviiWEVy3U++ntqM+++1C8vidqYVzYmX0dtVSjUQ08BMXaqPoRItntfvLZxep2
gx6AVTMpHs93PqBS/BgKnfxPgcUaK3ufkAiyZHBLeDAbQKCnKYkpECnJdyDNFLLc
5FLaShGJIIZoIq6+ADXxBiMsGlYBgHHQXKnnqYiC81fBhJh7roRGE6Ios27Nb9TN
W0f9qUpC7irxXE5vg55QAR2VpER1eqsRrzDKUdyAPbfBQ/F/i78UZeDaYsc1zWqp
m1TxQAXoVNR6dvgY+bRO8neT+B6kHxACWmJUgtApU5MR6a6dgGuVaGdAYEKOpVNL
TPpfHCN6OwQn4Qc2DCMnRbcuOsmOdGNcIhgjdQ93PJTx6M5/dSLJ+v9gz249fW+3
qK1VZAASye06qUjuZ8JVY0ntFb/xy8kFoiRVOWYOELiadvTaqCsdTbehjindFvXl
cb4szm32pQJ+SKCmnhAN+ZikWLQalVF0AEizRsR2NZfgoVtjekuU02x6h5AAvXU5
nVLhszrBtdtA9wh8nCUSh+KpIjjUMVndQl06pEb7EfFYkmXQ36tBevyJjn0pjgxm
ZISvbM0wSKcU5I+YD3U7bGHqbVzlI0wL3vPEknyMMvI5ugkYi6e+1uNXDYFQlM8h
fJTkQA/dM6aa8yekUdVcWwpy2PpcXrN1ehi19lQW6ju85ewDcaTVLkcEHqnuqC1s
Je90osUrrttoMTtJ3YxKkbVLpOeE+maqIWYYvSd638wwuzGnzxHVj67kdSDSKZup
ojycLyz78bT5xmYcPhX11pTh8hTTFMGHDYxHaqW8EPpS5A8owX0Afns1emGm+RfS
sQ17APOKHmKEJ1frEfEJeEtgiIDA98JOhjMJL+hyCGyE1QwjjA/xEgjDxJFIm0DS
WXAyWwP7V3umYu1JR+3xjy9yfIkLhl/9G6IrgJg1aOsNACBR+O/v9e+nmxl+q9eO
Zbql4/CjrCS1tsRSLZ1KtA1AAXEVcWY5j7EKJ/vHWrIgr2HrPSYKCRtOh4hVaO18
h8HZMq4qGOo/sOVNutUYppmt4VkDyjD+n9PCAklLRv2inxot1P+yPO5wui+oqUdb
T04YJw1pR/6Hr/j9SmG0clieF7Bxqiu16H5Ei9BFFjWaI7F5V3hO1DtYbtZyimy7
fxXNAiw2nQh69PIDDNszd4uP5iHLbyvtcV0lbpWRM0gQAjCotQLlGsoo0VYzXg1r
C0n0RLjBd9Ff9z/yVD7GWjnyY3H+r500d1f2leX79YhLVorzHQe/F9f0eX0mF2Fv
4UYaTIDTOB5gMSI2OIDHuM/Mxh1Ok8ym4VPgGAEQJPxn4HSLGzBJFs2hXmHh2ddq
383wiT+Ud89hkymKP3hK4qmFHvlXDub8xD0l4C8YtEIYtdIxMWgGmHFXW0L6gnff
cPkEK4D0KONZItz9Ro+xcuNJf/u2Vrd0aQx17LXN1YSNRdr0hOhVZtA5BWXsu7Dd
zEebLCRuEqy22ZFzKugqCvUWukwEcUC+G08d4ElrdLBwZZ/68prqaIfG+Y4CNqzM
wp1WNE75prqWsKXkMYch0FV8I0P5wijYjYH4W34PZw6ck7nF6Gxli9Xk2UEyRhAR
2jtVpjp2Opm2puJucwRE+F391rZ80ptE8VXJ17xi9purmf4xPWZLNvM/onUpb0D2
pkSi730FVXllJwEOYIgs6+DFYocTh80IymXxNypsnlnPXolkp9EWusaAT1mGgPSw
SNCHUsUntGOjYRC5zjhxj2uraKaY6RpJfs4Q++u0zdIBB3asny4DqZQrcstz7VHN
9EVrKZA04EzAmL5aPStWhNLqAwTtayhp0WIyEYyCDYaNj37kwtp6eyzPHFbp9dNT
r1Va1X7bYlepmppQBavkG8lhwgTtg4yG03lfE7VdkaC/XspXuUcW/gUL8yZnWDIt
wk6eVqqxsnen+xHflK2ZI4dK3IN9iVRxDYCq6xdy+zSpuYULuyjPF8A/fZMSu1UO
65YSanoJThFsX13cxP/vjQzMXQu5KXhYT0cSLZAPB2HyUQMYSMUd9/9oh0+vf6GJ
mGUiW4bLMuVi3x+/DDvsz1qwXlWyJMlbgrZJ53iNcOx76kY35N3/dDPS3paur2QN
zzABGA+vnDmmSWFTjJ0eDnuM7wGFd2GoJEusH3jZYu5vpHjEIUha1O+sTXNw8Vtt
0FyRBys+QB/K+v/kw0svlWfA1eakZvnbmIAnrieKQufZxq6i9zUiGKUl42ii1vfd
xWzqpTnIYMj0jfJ5A/SRCTPfsbQnO/Kk54d9VDHiYru7pAdfWaHAPynE1hGsHgg6
xPbDyW0GRiLWZ5BJThfzMOjvEG3F9pcshx1wquOSw0PaAFtqEf5BhYa63YV8ROJu
3HUfgSQyXatiyKUUqI1GMrRbdzSX9hx1G1P8rNjkPXEsnG98TSkXHy860eR3afNa
TVLc6wDQZ+lbOy5aIg6JdEqm6N6bXgsz9g5CWDygvti2I7CtIB1kz47BA/Udvd6Q
krBWBLlX8aZj9gXE9dccYCC2tDz68ORqrrVTeIFcKTxryKNGHEpvanggxzjb6ZaO
H1igivAxO2gYW/bpsF61rFdypP6DEDDZybGVIDTmgu6xp+yuQvmrXcrHEwsOw3FE
Q4JNCDkrTYmxFI+NP4YWNX4l0EqUKhUKASbQPfAP4lyfDkg/UInZgfdiZqmkUnyc
d7306lF/fXU5VtgR0TNGD/ZFnMe7bZAWqHuR99vhCk4KlkxSRnOoPA2J5j9cjr7Y
9sYIaNeBOt4l8b7ivcyUfXhCIo6ni9RAS36c6UjhOH3iJ3Bf7ptCCdfg7bIwHsCd
DTcAnmlvBxntw1wGrNUP+kCIgspNfzj/EBoWtw7NaeUFBfF1I0ZjRBvCpQ24ysE8
htAk8AHxhYK3/SpmCkvnjzYFV+FLa+hYHyKvhouY78izCoCzNnrid24sNaQ2SyH2
n/U452PpcWRhKPeIJElT/fYnNquAESV/PAw+/WOfuFHB9b6xYHFsEv/H0RMWq2Ix
U/1SIM6vLivuf5ctLXlhI4+zkvn+qznToFZRjJrotPes5CD6sbMIwMTyN7viFnBD
tZRnueZ3ZPGPL4aUfuV6pCluM3vusNbeXsVoUEB/NmBpDZ4fn6JEuoCAnn8i1tUP
sIbOW+OTeJQan0q1QLcLQ3Mh31VOhHYN450wzEC7ClAV1WYaCbewp0hw4hgsHeU+
NnVGDwZ4uslrIFxZ7TH/aDQ4ll2W1vIr2QHH1BP363O3g+DV8eaxRu/7G2vMeHWP
cnSkdpPUteYTmeA+PDK+UQI8Ajn1Pt24M5vsVufFHYnR8mv9D1pCtGx023awtkWx
ZEYIiIK0AULP+TR3mKCaLfTVXLO+s/6hXJ0PrFXRE5iANPB0dW71E5Nf9c9VUmr7
GeSoFpzivM1QMfymExAZ4HOhvr1wFoS1iGpn9r4AsMPwwk70IbGf0zf65g6p0UXo
Ie3VHBK7NfSx2I0ZvXHdWColUDJXh9utp2bqQMYWaWCJRs9+/SceaqkFGILq8dru
HSDq2Hl3dOnc5GuyIa0JTHrLeBf7+dK8eag7O+vq2K5UsNFxRCPIexlZKkse8+gS
dJolQE0+nmsfpN2nNMdYpbt4UUK8pX3ku6n2uOx1qYFEmsi0hbiBEUsJnNGBap/J
RTZ4KtFIcrOwH6f7kQmLVsq5QryyWiTvzvCN1CKg6/ZgH4wvDDspMVeEgoSgq2Tp
UVK5NxIZkeeObBfRux/4P0oJE1o61sknmOD97VkNJSsTofjtQoSvF1J4lY/T2E10
vK3SlmEeoDmaKB1lEOZAhfd+faEwpC5HDs9OfjkSkS9yf0UXZss1sbB5PRDQqvKd
lIpsbj2i8Dx3L470u2tbaouI2kAAYx/AEAn4GS/1cWT9Io8k++//TNoBuasjcBYH
RJC4hALWXyS6zdFpbgUOyRIgp0hGnnm540jzkmIvrfyzzF9JO4UnscVmvXmALlL9
uSvfRuuXXRpanJ/1L2sNlz/SNaMBiUGiyTTHYqDZAU3YDxP+UMIH1CrKHP84mTCz
WQwa29BfgQoXzy4Uq1wmPfKwsTJF2ePZ/eM3VmukfXMLwydJxv+IWwg0IUyu2AAZ
2sN/wGBW4q2k5i3UieckgI1SICGNIw+cUvxbOmiRbOn86a8kNovM2nubBjXabns+
8YJxf4Jgrmw9dmdxq6iirOOShngRUZVpHDuUv+N/+fuQP/LElugax9CIR1gzmR3e
MTblz+b+Zv8ysxMiQ+f5X9/2sfCjmBpXl4/56FcVqXtgo9xdz35p0T8rZxEqZYKJ
HoPJp4BuiPeJWRnN+EDwUsL0l87EHU/z1HSAADNJPOGBDCqHAL9z73w67i6u+j9E
DLyG44a3X6YCelawWNFuFysQxbDDA4Pd4An7GJwxOWfYiE8QkH0hxnJ4JCikVo/Q
i0kZs0dfVZg/7RadOCvy6yHZuArxwaAqHx2a018qqxWvQ9c8dpKOq3+w/x7NAprA
y3Kf/krGaBFLiyRgefPfIaP8JjrJoA3erqrcb05OynKqMbFGt9o1/hpx39BXkcjm
P08y8MKY814g4iWw2fFoMYRyPjESLojaSYW/LoXsgU0/Kq6RQ8SRAysKZbyN19Xr
Yh4fBN25/yzOroJVLXH1WRZUq+gg4Jtk20MY545DvaKLOEfwxY67+PwjBg4VVLUS
223wHRx7Y+ln+hAmIa8SmiRxZvN8gFLIL1I/yPjop5oqaXg9zPsnxhp73AGg21hV
WTi9EcorM0CJfB8CrtXWFOmqJ4hI2xqR13ap65GrI1E5C+IsJozEW7GBm7DN3DCR
vwWGph1bKUyCjV9ZogY/Mr4RVQ51CwC98Bidr2NhDww4iq7Vv/k8J21E2trTTul/
qD4a258NfKZzihnsMRUgFvFhB62U1KiJ2yw/uRuTUZGeUx5zMH8GvoE6uQq/WwLI
4XqRBK1q93ITSzYXN1dqxM33oUDipdE46qHyIzIii6lC/QUNp5fAH3qFMPMOO4GM
mWmChmsdPvGC+L44hpGzIJ2hkXSmHlOiMvOkSeKIMoUDU7Z5PIiPjTNUgSuHToRz
yduqGNddu3XRRQK3aTuEoODQufK4UhcjDT7LZxEUdPJaThnqTzeEQxHxGwXWmJEs
fnsUi+clS2UUKupMsvUbLnsZAIj8ixLCsh/qR3ZMu4q5YReo1ewSO3GmpvB2qHcJ
gzyKAdxyXiClCmeNlrZ2KO2j2r+sppLiTlf4E1pmMLOuELPllsWJAGe0pKilP6fI
C9nOaJ3pVC7DUalxJlHEkOy8/FIghZ812/0meyNHPotHTN0z4pJTRaW5sMIjzor3
oixt5nxnkhfHh3j/ahDTtE1TIgo0yadvPS4CPQfqZCiwWJh4OekcQEROJIjpUDdW
X8Qgl4Ca+CmKJLEpqR1rQX++52EoQ9c0TwJiBKqtx0lT2FMwteSE51uEHaiwUOSY
0J9CSfrLDkVCIvtiWCvLDNjoUS+5MD0OmMOJD+oq0EJclOCtNaxvGiZonWH9LYrX
PoHGcGeYkGO6nHYbzerOUmDJ4kowLj0naTAQTKV2PBFaZHcIRwud6+jiMxCRlOfw
ubaXfcVweVnziEv2JSss6A+q7SY7iT9jx0PT/Nl4pxxreCRa2PRLtVRKdrYc9tGf
enEgf+k0FdqSFPK+G5xA5LzoJiJdaW78/0YWcOu6hnZMYzIUnEFDAvybMB4vnd1y
BuAEJR80JR+WB9GdgpP/tg0BYz9WxcEuj7+2mqq8c+IzgnkYssxR42Ab9sodKPOX
YmiLXfBYbtJ4daJ0lKhAP1m3++xxaeAnBMJsybRoSK6KJ6C7tj8E+8/lOi242If2
9+2vFRDCCjAWy/og8qsJVz0QSq3aOWbhcVTpuWXCnwc3xnShYdpNlSldmj/pw9Cg
2v0yyAWm8kdb4X6govcQaMnoD1EFHyWWIjhLMgvGYY0KfBFYX6fLgm4SbJzlvQ3C
toFhaMuIJxZgu1h4seZVte8JmN5ffysar9wwQd0QxUw3pLkHt4jbzUgVjbMMY9Y5
EDIikXf0OglQtJ92Az0EUxyhGf1TEezh46KGvsDxwbJNBTJQCNG/L1P+dI6bGrIc
5VtuKSLTKB7jNS2lXuwQ4vojdBncnx5tFgrWzt0js10GCM4Abf1Xr64yrXtIUe/u
6kMxed0XJ9CSXwhT8eoDI1ojWVfOFTZS51yn8Aq5Bax266v2HDQdoBQ60OiFC1ml
27VHxnxG7SfKhtOyByJYf4c8fzKeDygWqME6XXaL2EnjiRt3h2Whl5OFgiPeCquj
ivjX39RWJcO/G/6L94s5OLFdflyqqrwfFn4F1hYRE6GK98TCrtmc/nL9voblCYju
YtiB14wku/Rt+drz6izoYSqUbX7d5xxuwB3tapbsUEm3tKXBQvkPNe8+IJmJtJH+
2ytPoxuTrCPrjL180aWRqp54FS0MGXKlj3gyKaHg1Ibbwb1sBolePSXb87Z7B5GK
fqDFh2Tl1dvtFhDeVsM7Qc4QhReXjJNHnJ5sflsnl69m+vp11QmQpV5NPYvihYJr
IedA+mAZ4R3muZer73YzQ2iBd7Olg0H3r5GgNUSyKyYrMER0O+4dGRdgZLr+gSwH
SD0rpjHdgpcr0tCc4+uMNSx84a7foW1M14qc0u+gogPGDrcFvO7OzGvVAUYec/fJ
VMvfJzpNa4VXeA8WmLdZS9EoEER2yWB7lEhYgccuNbGVl2SvdDuaZNiQG1zDpvbh
c1VbMolQoMJy/uFqUAdexLupyewMryJPRfGNxsnBK5GyrM3TvVlqa5QLw4QjnSCC
8lFXhuhnqdAQiTnLrlliSs8Sc0TlpHenFgd9ugBQ2bA6XJRJq7iCjwJTtYPXO9e6
L6AbSslbthCUPuNpYuarfVsUfKAlKTXOCDcx0oO692HsZ60iy8zX7UTMIVdIFuM9
4miae5XNDRCsVChgqb0VjC1L6h2nO4/1kECUMeMsLbV7X9tS4r1jW8C+zXto0BUy
rJLJwaEOIpbhUYtgI6gBrN2h1m/BqpLsX5ZxzWZcF2WlQIKpJ1177aqkwqzfogwf
aGvZJM9urVI90/2sZO9D8sm33TdRnsvb04VvTc0uv9dMgsmtRzNkPRnge8bQ50t6
YXldaWpaLlIpGjKdV7vnjMl3q1o5l1DNWXuEnOU5VisqM/QHTpdd/7E8IMt7+LhA
h5vXdo8PMpSoYwqP8rAQtsPB04czYAyDDvD78QXuzxqXUAxOa4NStvKafaACT6n5
7xL67PY+UMEl4VPVK8qfZCdH4TAzT59QeLWJ2BTt8MQO83JmOrL87XuGrm38XfTA
eD154WV7kMhNLQJECILooRfHPg5XTsa9InLGS4kogrTqQ19wPTLj6VFifUynYMm7
Rtra955+jImH9IlYcjmIB8YEmD/KdtnzwrmYrVmAZOF2XhjstS7oz+3XR696tUp5
QG587G6Q6Da3NxpbI2ZhOO1gTIxvdcRFyZvIwZrABAcI2FxsBe+0+5aPVAx8Wtq9
tCR9FtcycXKJRU0azkb3ekRCnMGQZJHfVEJzyJMlsxM5nT2bzX1ZJhWUVxcfVNt+
sHFlE3XRAnSGeknJIB1H41/ZUZ8iy9ZkNGJofAjqc+KIGoTnl9CefJ+D1SPWCuKR
0eak8+6Lr/nnMGnC3eU1WC9Q128H1cBV1ttFZPMYR5MWAnMXnIwMpZQ3ePeXjpde
f7O4APmNjr4p9axzlb3wVjSBf2pLYwwGgpQg9OcIJmoqEOsw3qCdM16ohu7yL1Ec
pLjyq4kGg76l4SRLfvYedUD0m0wu1/DA/cbeldRugYfAvugsNqLujpK8uh5KWgtS
q9qr9+r+uno1se0wXlWSGMG4+UM/+2wGRwelfxYpR+PCg1B0p2gKyGVwX2OEVGpy
v8qwKKVnJAlivOmTxJG+zFTGHTbtTlJvOh+mwBr/67WkDxEWO9rzzF/FE/MieABo
smXW/edli/6L6gNlT1tmPcH5poQ3qF0/0JUNLWNERxK23x6vJqMj1D7yazhH31V4
O9YVXVUEwsAYrhbS77DqV6PpDw1hcr5SBl8tYYCz5O0H3ciqgswcOkj5+0FZgARv
+ZDZ65OqZVHg4fi0qBFVNZa4IWWc3WMsMe0/1bOylNT8YcDdPTtjOq0Tzy8zcsnT
taSM5DNDxBWHeMvrTQ+4DYKNvfxzVU/kkfiTTm2vBbUKbq89P4ML980ChWu0f4nE
m8SXY/XSsxIA0qEqPtiah/e8dccYW7MXS/yoHq9G0F22q35P02Tz3g83aapl7/IT
SHJN7f1A8QffmGVBXaoFAtcF/S/VFdNiL285dpHcZnTycaftw/toeBu8M6KopkDD
fs62MsPuj0u5QdQshJUez55J1unk4/iOk0IIBSpgvuvMmpNrOQt99d2v1u+Vnwm9
h45hNDOg4iiWt+qsoA458Colt2a5pvO6CnyY6QJqr2leV32GRbC5Mrea7bVDGcpg
MCVI3bELJRsqoXj+3dgU59hk9Nj8bU2phVa86Vqo4osnirJMCYSwVYvx8b6ovzLc
CTbYzFaOb2yrds/afBnVlnhk4CCvFS4ZOAfND3I8jUsfBSsoRjYgb/BIe/md/2PU
Tc1QAE+SGJC+1KEU7YojN4FbToZimNr5Cchtq9/kNMbRuhn8+VeMK0DpX+u4AJKS
HnpDpWcmns+8G9Bkqafd+fRUhtpdvuINIeiWmIrEdeyrFoy2Fgahdo9kqwjQsH/Q
9D2e6LgLoo0Hz2DFHLK9/lrJGHSugYderN1HX+oY9o8a1NIL3y/zTkMUGkSIz/Ex
VLJis402cd4H/5vprjdVICLFFw81YUNLVWUjIbkxhyl1vShPCZ4dsHC8wgx4ISTE
ZFL3cbHjwtnCUCpuahcfLjsMOkiPoULcjOShnXFnfdXGtXdBAx7u52gZhA1TuNNP
nawmrKBf0cIxPhHJbwqKl1lQhmcQMfmTwApjwXCHdS7DlOVaUZBU+f62qG8unkh3
86E0WjrxOKvzKoB1Fh5HgCtVPZ83HZnAakurCesPJ00u/oc7urUBPWH9KNPQkGp/
ow6svsXyjWzXEutk2WKU/WFDzufRa/RixsNrooWRL1pkgOKSYC+4OzvLKQ4EHP0S
yVIL4RH94y+drNASUWH5H+WKXKDU2DmGwlnggPfPK0lfvEZ1EBC+MiDeAmR1wcpI
/kmRfkkcbNPZIWjD+zQq7ctoWJiU7vV/XO96a77D6yfeFI88pwCOEM+EX3mL9TUT
u2yPVQPzrQ6A5TGmjC11372sCma2180pGADNQzCXxq3t2Kt2A6gSC37hIFzNXvoN
ZHJvLdhqPTD4TwX51ZtqZrbaw2PaEEaCbegeVhTd9aPqfqRKys5c1jEMJC5U1Z66
jKeO1rXIlJKKZnotj/Y/Pf+dSwdKJkdWx1NBv/uhR+bI/HP4KU1aSlPEqfICARh+
F0VOXr4ue5DaaaISUtntLJbl+3SanasI/8GczYou8aWlgLBeiTGN6Sdz4vQVUQ2B
A7q3+Q+2BmcxpWzLrvcIzLl+mHPVfuLGSaPybPH3vBf7RAyTkgnlf2sUK5/H+l9B
UgfCkfVUVvLWkKPp/XpNqwPnR3a82bxV3YhIei/QUnw+Qk3MLESnG1QYBxBd/ptt
lwpOqF0Q4BM1fh5sjVTEBi2cT32Yb0ZQOMgM9ddPEp/M7VImctHQYC8NCfL5RVYG
errgbIQZ6DLPWTPBK68G7IImi5xlj2h+a/SNBUfqcsZ0tFZnrZhzAhIMyfZwdKRH
bjFmBMZ7wzzVxdEnALKuoW9+ncz9g7N1sEyqnrOosjtgdWnqxEIk4Ut6xJtb8kME
fiJzP3w8lSHKutoJWGP6SjKnueGjTGVuTX2RbGjxxvrui41R3LuUk5ps0r2Ub7pG
LK1rkysqfW/6vK6+xuXI++iIOoJY46fyv+PVYX4/lfZqabmggldOws4cZGki0Suk
B6dnmZehRBZrn/Fh8a/Shua0mCgDrM5509f1l4GXv4WojYYRWgb5Z7DIkXV6SE5d
s5QGexObVYN8qcEkB4Ep2O8gwh3oLq6id24RsHMFBVZVLdNZkZxsNkvcTfslGL0D
qSxU2lb9LOafPgtC2GhmYf1MDpm/5EkwFbDLYVhDNn27p1zEAKIFxvjG8tXYozcu
SZhiVbeDGqHBDlR2FczHUSqHuY+Ej46FESBoZeAHI/GVoePlSJodagIUKd0QGR3B
+vUOTcH10QfdJdalQ2T3I6YVhduDuJQ1aULAm5OBkpi/DVl5idshLEounwnH4H4W
2fPhJllL9q6eTWgzuAL94YnVENenEf4PCLlF2LcCK6WsptXk8FFO1sitoy+a5acg
X5RC3yJB0B9QSsyt3rCMUvmC1D0EFjQzR+9+pBQxlfPKEWWWXNINGW6YsEx9tFLl
3lr4AicnrqcfbUiVNibS/1xqF2kk6iMzUP5VtCe0D+eBJZKd599U2ZZSRVnspODn
2E0qTNlx2/dkHCKJF/ZTb0R0DkvUtXrU3U8FCXjWvL/Ns2BodBXIFe6wLh81S2U4
3DjEeighE4H9NBYv396CVBVVrONDybn5eFRVPHS4tmOwwVhMrQc35sdv0VT9LAkU
0R5MabMEIAH72+LIH3LdvICg5WLOAWcFnghGn4AtESk6ErM4a9cJvclGvRwlNKKm
1UHR/rSk86m6ZBuq2YIB8wzbs3PyBU0UQ8MAhyuPPN79zQfKUlzro1rwfm1aeXH5
rSffpMw6pfC+MuSu2pmk1e0k2wH3FIuaBNHa/K2Yj4vfIRrSBftAKwRAOwitu6/u
ogCa9fLlw54AdJB9czlniRra3lxmrIJ/TWrc6CIM9p2DC05LqhdwZVJ9cGuRILfl
/U5+JLBrFfXtS8XDjvLd6J0/YttihZpPEFJdtjIg+EKMeOm7dsVWEtNGBbbyFm13
e8OHBDBQL4y0SHfugLhdV+s5X701KOskX655nqI2I4LlWYVWv7Ot6hSeN9urGTY1
lEPKgLi1yzIWDl8MTIi9n3bybbjKee5sXcouwZmiRUaon208a+PGrqtDoP20kU2s
MBU6BATN71PE8sen2nd2TzY4a4oL+kXVR0NqGetk1mKPICpEMASQRlp+6pHV1/Hp
DcDw0+0ksekM9bS/T2iTYBu5BWu7+uX/EsMMxQnozSsUHfLW7s1xXLI8ns8X5UTC
tc13D+lpF+40W4WOTRidLwAnx4IwQnkYVBimuV2LtL7rGnjw5h3SXUrpT5fuFPk+
HvbVPTGhtRU1XdsqaRrZzsc6ODr8NoNBwpnjhguG4gOfQPtPycIQT/UzPBxx6qn4
azsfM56Ap2Vyv8AClMlCTF4E0EOj1fS/rVf2qHg2Ve5hgI0SlHoRi303xE1Upf4X
X3pRxfytfC8PC5PHjgd9JbvpFhkC8uu3+FzWyWjJfP3z2xn1fWKCUDGfEFte6/tP
wLkoOSDZMs44EZg+I6Jeaj4cWmtGRznF1agU5J702caNrYFfSCrnLeKEQ1W+hiKA
6gM7qu6z0g4FpnJMwV0aXDui2DfZIhW51eUfYXdYBVsKeaZ7vkWgiTRPhm4RYsM9
t15G/SkbZBXpbo7x34hY9ESNO+lTFBnxWsxTTTQN/7Ji47/ZN34nIVsZuch9lQks
lKfA+iSCSYiJXhcivU+Pnc6OkcsmT7NT5SuOroTgCAyOpXLObTJ+omqwQ7/PUtUr
S1PPbM0gxWYgBIdRCA+G1ZFB8P/19y4UHqfmhoOnN8kB0xaPlk3RI6InUWTzmy/S
yudsseheKgY6Al/sem/11LYAFlNbXTKXK9ovMp7d5sp8UKJnwUqIwzLgmQSoECsX
4CXPKrgtto8Yj3ORD6QTBhGuFBqSejpn4Hcg8I7B1uwSKOPhF6SjaGMKf4mavkch
KwyyxjSq8pLpcjDEtzrdrqHfE5y1nKjm1iE6x09e3ciJCakSC1wwc6cPNABK2gBn
LWTZDuWWD07ZweTwaYCN+QaV3rXfy6FxZpLjbRG+s+pbXk/1ErK8B/LNmiRaA+rD
b2elsgJDxdsneLNMpcpoEOF6hkDZZP3QEPFkzcdJl6TF4Ophqc1EcXDEz37tML6e
Ubc+8bOtnMOR01OVrUuBTChdZX1qWjC3O+CzZcB2xQkPSIrD3R1U4PCQCSToojRF
W0Eonq9nWo6Or3oajYynJfDTOI0eay7joelznAFORHrvGa9TkfC1nM2Dkw4iXHkw
tdvOlwVk3GsNqhz7AkbCpkwl15rcI7SCzVOAp1q+VSkdxeXc2ZTphFSXE4cD9FJ+
Rl+TX5JA1mP5pL3o8Vu81zaGNi7ataz5ocOI5GJG7vD3+J7kir7pQ/MP3Oqiyii2
BVbb35lMvMMhkcPvBBPrQXZGaGtbi78BSZ3wg8yl22X1sGYv2bgi6Tz2nV0UxDHe
fgBlVErp6lWyhPHtEpYgGBVeirwWSh4Ot5LxpQTbZ6aFajXg1J3ENDciu93DmJ0o
bf7IiTqZKS4YQl26YNiDCf4d2KCTupIPCn4Qq1oZvHVjYGZlSzhI1i+31shoVGH/
1HYrEDJzVasFQ6sLOoI8CH1ygTQ6NetU8/pia89inqyq+vvCBfGJ+SNWAseMopdd
h5vkK0P3YqMgMojxtM5BbUc/BR2+ZBIGgxqFmrp4JTYoRcMM7rOSgF+55wSrZAiF
usGL/qEfQx21Z9lxEQ+k89qWcCVMowHlt3au9dCxDLArrRG8TnDwtyK1olYBBdhz
uSQs4jQDvlgCv1jggBdTvHuG5f+vFlslAKvtB0JMmO7jQ6kVuw7F143jnbhGnscN
GSEOUkUSAJFLl8xvfduKrTP9ntRPpCTTm50XwMgcnzy8L1BxfUvqdVYjyr7yYyWm
PSaGuw6UWwIYaA+2uIOC27H1NMpTx2BpXQB9km9MQZV3tj5tRNGRoLavEvCv0Hdm
4RgGPJy3CjJkfFJy6VOH/Nh8ZFp4xCJaw6piwTa2Eedvi/YrWlQToBrvwWzhvFCl
QInaS/TndpG12lyuxtuwc7fy5FZF+b9DYF9Jfo2yBAUJryGr4ZzcTZMv0uFgWDbC
Yr1yQdtA4xoaTIKnzaQ8kkRENYqBtcjeN1Yt9pZ8lk2FnPmfr+g1z11HEWnzRkmQ
07rtRu6EwQPV+GvcMkZr9MTXrgV3xkx1aOdQuTK+pWmA8uEQidLSyH5tIcaxpMdV
YveAgfRO678mwsNSo45NWmqgHgWb8XoA27LEKFj9f9MvUwgMDOI5P92047bmMCAk
FRLYB7FSh4jgvcZVtJ9nlUhsJDq/0TWI8xLX2bxnGNuUIFTj9eWriCnGn0TMm0kC
AIp2Edy99EGYuGvhyIpE5bGMvv6DwhHXBgo7eGZKuCOGt1NRoSUVVNb2RmaxQEBt
bp0ID7rbT8Vb1UZ5fB8V2+8SGKDr5MYNQ28loctAh6oaYAgvXDwAQaY1B6vwYs4w
E83xiNkTtfibjuA/Aug66c+fNeDPZQgcr0ZcqHzmfFglbOe3SNNnAge1cjXYeLq5
x7fiJ4BlHbBW0zsa0HlJaL/DNBm7iemhL1Gj+evNuPbcLPM8seViiNFUIL3dzyed
2pDy0rR9lwsL6I5yeM/85gFHg74iffR5oNg7zWsx5kbFFlhN8oTWFVMRKh9Xqypf
dl8g8rwCpN0qnDe1d2icYZrcFrm1sijVeJTx595RGmUVHG8HmGcwTEVYW8PZU7xC
n7aRgJ1paHhMVsVbYUkALV/pcxdyv6c284tRzni317BNCXhm8E/YdWsie6llTX7Y
XO6nhktmyhLpamkCzs71sYVgz23SUi6+ZzauwsI4uwEWvasCjRB9emC4RZu0IQXc
0KaIOl+OExSpELMoL7pM8toQJvW8Ph4m5SMfMNkdtnxvni5F+OxnF75H9RY1cVTB
eQDmfLWFYXFa4nPd71zCmENpi28me05lppyn4ytad8bKboMffS6/pxkWZxtQ2Y+m
lgmqDv/3nQ+6lwZ+20psci7QroFkH7AwrAgeZxsHorEGAcpTfPri0mqyIak9h2RE
WGdA5aBMQnLdAuG4J1Gsju0fSrc6KnCCTQuQQdw8l8JdyNvhpONt2dtEogioUhVO
q9gk9Opwqr0u+goRULSTcdeAP1Qx7JzF6iU4MrTRSjKKXltjXOO+8OKLSIzgc3wN
Kfp873f5JZ1HRP179xA2qLSVNJ48nYTG50bbePV+UUpNgi6xlzamnt8wb1aOMJtC
94pR7A5SYmS3FT3diQa84cxfv6UGvNbF9Rlf5dC9FiqzK8CPp1ZW4L2DL+5HcHil
xqPqqNEbJldrdnzQoz0RgduIZod3q3SRudx9JPCoFmKTevkulUQlOidVlIOWgxif
31emAemdIOoUD1Ga/rMesZjKJgNEHHo+vbOJD4wUPv1OHu8ibGFyM9fgdBFg3PCy
8fU8so4mZoslaLRIDNzqFq3RkUi1eCUUNYKGnX73bJEuotnWA92xIr+d6mL2qCGr
0CTN+oJk2TNeWQm7bhtK3jBUrsl7Dpo9PZbFcTJPk8x/VOXebGqPuWZhH96kmwP6
YEjQt2cbAmtuUgt5KS/tRhmpL9FbXunG/P2dLf0F/kvnvbsMM4VbhUHct9cN5UtI
84PFonwkkAchmKEBFHrYM6UO85ND/FzgUmlbHe+Loz+6dhcoKx5PMPgzkUJYlP80
AvZ8QNXABjytbwPXCEl8WEi7JmvVImquwNTtzECKJ547okASZMNbTgqWBg5S81q1
rclxgW6ep22jIod4DAOSf9RUHlWVUpNbzlOgIC02E3H7JnidvFXb4pALtPnaDtqu
dzYlMJPM3shUBRVBXucyo8GTF33FoHy9Cn9dEfkJtw40+YULdiIppPxrLqk4evZL
zh5UyfPHK4GTHKvTkpWEaL2GaspoAIFimX/z6K4TB31zwlskOU3a/qWbYgE25ktF
5eWIWnZvisXX7a+nTR7fnMm2c0EhcgX6RuTQu9yqyXeQNIzo2DDtxczW7LUbM1oI
d/GfsJao+gx4I5tuyxLwsOhRWpQhctGgLuok+RvW2I9UExS8Hd4G/zz6KQth/zwL
xPxvJtLbb3zMHjJBuD1NlOpMHtSUXiVSzfNV9aBVLde7sOg4tToj3LsudMZkjFwN
9oerX/GssF02wysxe4a3VEjD5Qvws/Rx16RwmG8HXHIdIwmKjlcGA5/GalCj9rFm
tKLy1vQe0NO73lXDP2Hh3Ln8oapzB6Hp4ZqQvlogTLu2Zg7pZAPF16dzp8AEozas
VOzGDvHrnkgZlfn5V6ts9I4rCeXSvGFYEX0BP6QeqWpIh0UJl00Rlp4JFd7djIg5
TAcknQevmbzdFnCp2C8tIH6PKViX8IQZ8dk29u4UEoztAqvahGkzzD069otGrMbS
DPQOw0N57enBPVTiOXRa7t91WmE/t2z2KABK9ZizCyD1nf1EjKj04/dyxpQPjzGv
6XOsNYMVpxq60vDVnFYT3NQmGr+5RxvLnNE3+biAWm/iILEMNS4clj9ykbnGFCo6
TGaEWySvRiDEIDTkUsHhkHCvHeO2VU+wt/hFrf3kfQ3TTNBGH0hIIIQGyEvd5N8W
Oigp+Qh25fP8MwEhd6E6q327PY9s7ThjA6N0topym7cUYIZi5qQRO4reO11MpQZU
9bwaIvCjyorI32/U8XgG1uR9Y9UjVN3k4TDGBU1xjl+h/Xrl5kLny3Y4zloarFaE
kQNY6Slh+41OuR9zVspDq+etWP6/OgmjvIJAJvOhQ6HWFu1TTWQeRTnbFPQ4rgGW
9JITLslb/vEC3EIVPp3TDLqAHXeKDvKk35ug5J3oU1EjXyqhXcDMYFsvxEWt6F2o
uL2A9xeWkx7vw7v7lKLN7Zjp+VEuXg3xy4ecrHpsZKWyoJz21Z09a+Rb97DjmfUV
LWt4NWxVd41mWPI3l4H7b5cCbCCzcgPxLaHuip89gYCVFSerVZ61Nc+iQ9XlTcCC
j91VGFd8hUDlQZF4Ue9qpsmFFwuQHPnhsdEkFbM6sOS/WT8aUAQQBoFT0dpqyxie
8uEcBMNZsEit8WayJOWvUgjX3MKQ/ZkWR7zR9DegAeTh3x7EF93b3OKzLmpxlUPR
XTS4RorgiPX6eSoeg04jt3cnzCrQtNSLUB3NHDSRKbaixKYDdZRS3xvoaNFonwov
YmKpwo4hAIRJAMKtYzhfKyq0NjT+8Zlhgt+naXAVWQSuGqOcLwHtmQmw/vDjA59N
5aZ7v7EZnJ0ZhWY61eVEPuvfJh81R3jTrjU/q1q9iR4uwqBNlVLw9pj6wT/MRc6v
3TcYdujsgg173lF22k0H4a9QJzlEsYnaAs8WSSI8EC2XzFcgsF6XK7GnfBWpOpv4
hvd5wskv+/2gJstMxuD8Jzf00ryHacgJGmB1ofCu+uUyIqo7Ujkwtm/gmAoO2hbG
Naswn6T0rn96kFzm7I3y+zVgphqoEfp9dJqBYCIy/RgJT9a94pW3QZZZj1vYkmQz
USlEaiAuSwFEsOmhihVAAnsHjJBDaFi7p1y6ClYrxnQu/xQL6d2lqi+4uUhROht+
gQlmmU7taBZPBjWwqP0Uyg8Ww2AYF0EKpgowW3Un33j2pdrjKHPwsGiknw7zWMrv
6FDY0GNoV6EvycVr7NUZYWxGEtKJ+E/oSl7A3HVHlel65l2jttzU/gzV77vVu1vv
YdaZeNsaWYRBvdo5pnsxdxnSxGGV//bqyFXQXsX1Ys4r1l16fcYy9CU10oKtHxMH
tWhYXzY18oJ4LE6O41soPix2dzC9d61RORE18G7fJOVFd7OpOUQUFkQiohvnhCwT
9KsM8hapF/h2cE5pOPd4PRBSy+C+s5g43JUmIGb1dN/SmuvOBHXe8RAH7Y2nAlrl
TYl6c14giTy0ndeHwih5VE+K9tIgOSv6GF3MXx8F/OIWDuqbTezmYTtIsvrAOyN9
HPei1wsacLr/rEmVIriNbY5PGelodNUAt3mQAaDfT/doQoVNCLvd16/qxOnx35C8
n98X7rPlVSrcdAWPR6tg805W2Z5XpnoUxwWkvSEPyf9fh/1UUSULZsf9eR3fk3JM
cYxJpUFuo90/l3hqdxko4FxQM82Em67aluUUDxYZSaUHLCKssofLlSvLBNYI5Qnz
parOfNukQyjiDEQuH0O9aLZHlcMEKOFgxtkwFXgDZIunK9uAHij75+wl6OpOyt9v
nH/jEiJ0D0NEVCXrKAfQx5cKl+utLqpRQSFBAC6a1gubTUObPy/luuplNEbTxmns
XByxjWZ4gULdVEMtIs4Mbo+iIhvA0yPirctVbdCJV9ULW2Uh9cjnI6svGVVK3Tux
3QFxsd5KDU/5t2pM3RXfoiOjuHjnVWBMRSb1cM5ljDrMdJ8g7q9LBIdXxHbbMsXC
6KWonIIzjxmpdW+kP//zRHBZyybyQY5dhJVdkPUZtBS8jnIhdmahjt9t+duBqjv/
riDA2rZsU/9nkJppG7rH7n01vPPq49m3ZWKQgksNx19A5nJSBRziUk75LYNcUyqs
wixPkBxAVrcB8cVDoARMhSMMkaaXMhyAdIonhDyg82amum2bJGHTbz18Yw8IVTAV
Odh+jXFlQxa1yzWx2fgTcJAcA7TlG0Bv9Rc5vNpKc+vcJUdgyI9gVwE0pAgGPgJE
CT11X2z0Fsn14VpS4S+AGZLSyZB9PelFnAglAG0HbbHd9f2P3U/eg9KIhXolq0oT
z+ACH7sqyKfGvan8cjPPa9ebiT1biN5Z7i1IKLo3h46jOFouGApm8No4MrzmiNt4
70gUuSdb3y/873XejrnshM13hqI+wnu90gmd9XQjL/3QrEVw9obXmy44ZYntCPks
jr8YJZtuPNphZtAi0ym8l6dFIGpKYJ8pslHwGG1C5SY083H8MVRMqoHy9qwhufya
jL784DTnt9WFKz8M5TmlEQBk7Sg6DjoIfDTevS2Xlmguv5i4//tfFtkLblAHi+ZQ
GJMhOmjp0pgqpJ0+tNnIihHXqCrr6OZEJ+hs3foi7OAYGwgq7xBXk5Nqrq6TsGJI
h+7VUmhI5U5OHLey1ywu/yi53cu3Pkbynt0TKybL4wsLIZnvq+1P2DIZxj6Ahs0i
tDxUUW49m5yt2/A/XpcfR2ZKgYiwAGO4ex7wzxouqC9Z8GkYglkBjKcg7vz5/1bC
VWtCuKK5lIxIgZv2/UJ7DTNnFbSdD0o6a3yAPUhrGzn2pbXZ3DDyQhce4x2vnen9
cmGFmsm189eNh06ky8N/U45QEnWVBsP3ot8OPhBfP9qMLCXuHn1ZqsfauiQWY5Ov
7dV9PdozOSZMYvJ9oJbW4csTL0ERVlqvwmu6MG/tUlkxMM/x/h1sKXXUiBv4Xght
ZAN15s4eRjH4dKx+x+j3ewiejsNPd+aRc3ObmuKgKD3zm1cDFxq0FuE2mEPsXv9o
BMEHIfvIKkhueaejmJovqs6RvAXA/kzoGw/c7ZX7MdS8eEvrXIaSYBIemAxltv//
hPr1avP+B5vH189muIKd/N5gVre1cQYMJe06S4rfdRYpFxf2MTz6JOVFgyldP5Xp
ko9TmIYj0zHYJLrEqQ6Cz1uxb0SC/OP6P/N4DpckicLGFGS2Tmi5MWcNLBD/Yv5L
v9QwWQ2K9sWGvc383kFFu+oPHgX8pQagU2xRD189ooGni9c0A/Xt1FgttuuDdU+u
8VivmybEtDSDvlzgDTOof95kw/dAQBrn50Vhl4AAdRVPJsAiGD5I3XfDShVX31RH
VfBplJZe8HA9UepXYGAus7sPTLNO80ozt+07Vb8ZI3GI6q00K/maeaDpXZdG58sN
7LnwiBsQKps2jWAD99iEYv2wOwb6Y1dAYJLRF+aeL0Qk6QTf3mRtIwgWgo5PYJBk
mj8ida8ZKFuIkdvsHv7F/zm820ZbaIA20uSFxXzlDTh/UlFDj7hPUU6hnnyS8UDF
V4onw7a2rpkQ6xQChFHyWLFq2vPTV7neg/vyRq9Kb70+cUcV4lSP8r7YNZGLYb5W
chj3jT47lkfjkzjJMCcVQSKIsZZBIvOZPERkqKJqFUWI25K5vXP28uED8qkdRjhl
DlQT/Mn6KpngVZFSeqJpq95d2K7HLCs5Sur6xbb4M7MScwsDlCDacxlPDwLbR8V9
0USH1lL5HIo3Q4jhfVx/NWDpr8L0Z7QOQGpb6eNslKNpBWh5h9mNmd6z6uId1DmT
22kVy08Q80Zpt4xcXEWJZQOJe1dc18SWwGPoUeXmsmOs9Q/J0hR17uQoxJl0YKje
g8BSCw5Aw5Ro+0i1SxUv1yfI12gJoTioUcKoLhvg4snC4jzP3nC4/9FDfapkxg4M
Gcf1FPnI2cWXaZtAVRkoeV+kT6OYlQ5x8Cmv/iHHlHODn57HUouecT3ci1H+U5P6
qruA1fS0GrHn7z+IWVFzM2u2DIU/pB2qNFXYytJ9xS4Ggi/Su7okMTQXmpD7mj1A
zM7pQE0EWxnkfh/pvFLrDt/7rQ2brYhAKOsL+YqcT/Bqxhwo70aTx7x4r6MmzQ0d
uh3LF14daxSiN0w0f8o8wvvB3rIo8bSC/yKy0sD4AhCQct6MnwV38sQ00U9f6f1O
yUEdcf7kZqKf/2jGT8qqzrawRw/ZTNgMSBJyfXCRDJ1EapcIdstGV+OKdrf9b2C3
QJEy+8Pejfi8DQGJyZ5iLhOQ9FI6VpyzhgRnxvjRSWluJ5xpxSyHF67Yme1JtiiJ
XmG8gghpngtgQGLl3ruIXl0gp80FDPfJdBGqXGwH1Z/+ZuLeVH76f0wVuzNe0z6G
LuWfbhiylQvQ+dy3AZgWCKjvMsP+aL9BxOSH/IszAPjLzbtNO+8YlLz/SCbeZbOP
zCmzRwrU2QdR7hTPLzfBZ7IkSEleCRxtWUdwJNro3hNZjGLTAV4FF8htDUHk4z5W
xxQMcJs/SYGjzuQx4EAx3FLTLQYIL/eG3Jg8IQknXPOJj6WUj+kG9yyGjD4Cdrdv
u0uJ0NFDuhf4bVy+owjB/7wOaxhxkoZBtT8R8SjsHvw642fF3QYCVR1fTyrQy5Gt
UC6jWLhaFojxuOkfdyTmzog+oi5LJgSnYtTaXwF0CL2rvQu8hVFpN4F5k3iiElxx
RgIHXQZVUDgAxY+czgKQHfLDPTLnktUBKjmc/6bG96HQHcxgV5EMLDuEN88IO6GB
zdnSD3NxAhLj9CJBfY0RIrRm9Eb+jTEfSeAALiCsrdWFXQJBlQjXMSSmNolkpqKw
kgF9YUiIezpeNRsPlcH8W+3n6c8URcJN+95X8Q+PuPBFoftl97YguTtF7xHC4mC4
PaBiN2vcsVXk7+TLXMt8Qp0Xh3MPpXKxiZD7QVlEyWCLorB9bvjg5aQN5XQMlWIs
vIqhzWlGuKzbdvu9otKpx7YyBAVcVSAxaPE0P09RPW5FS3kw1AQoJIDGMn0QR2tx
vgb1vQtQsKfHmwtFeo83sb5A8wnyNh32Yxt5w5L/ujB7D+Nf3F1JzdBSK+G7HANB
k+6tILuHNHeN8v8xs1gtJUC9x+GzX/5VvBd56wDZeELWdT5dRDyQI7UXyRB0qadw
xDnhOrMD32WPWppKjJ5Ynlw/mZtiQ5jX97Hhp6oQp9kJKOArExKeErJA5sPVHFFs
d4qUg2o6OQ1brKs3vkbwWQkrURnd7naSAK+0effLrE2WJOR3ckD4XL+aFYsNehcb
p6X7kayCUs8bgafV5pMh20At3KWOvpElmxI+LLuHoMp2GyCl5XVPJX1bla1+ht0p
4aBBm2iUX2eP83FgH1lbOIqRUquRFlHSVjqHLv9Mptwosk7JtWaimMTSSJFpZvMC
O0l+PYvGzUGvb9ZJIiTGhfgawBkBtZuQT5w7Gu6Yjj2VkwaJNl6NDC66PNz4SzP1
O7ALPy/ypgZjzoLLuSiBzcieH7ziJU6Gzq/ESbNcPd6VeCyOKei33AxNso8EqjZ6
bXHv3xwD+W/paql0VB+spROZ8590+B4aIdeNIOGbTxCIvWmZ79lIlgnprLda1ira
Ru2D+TpH8LvBQ+N7NOVebvOkLEEdkVbZEgNjYQArglnYo6KENCDMRsl3JB1pZ2gb
uEwXlUM97EDsVX44NS14X795mnUVfQQsljTXOu1KkOA8GFTNeLptqZ4PGb+sUTg3
FHyaRu4FxO0AsacViusGSQQC88pDKDWlPL/PLqWOGjtiZfzTbJrTW8XxgEmXptMG
LW+roPes4+S2EQcADEjAdPpJ5OMtOFLJORgHk34lXvpvpvuoRcu5I38OaJfBBfkY
gxMTAsm+U6Pka0J2Hiu9hhRG+eB7SeakPqqF7FgXOs3bvnV6tm70mBt8G4Uh8Bm1
/LwOnBOezzTpL/z1HTJJJ/v3yTiPU67gE7zmLrYAigIEbsTK744uFrn60h9lQZwc
gAirL6ILJHXgfwoRaVJq+Mq3rBV1TEJamcs00jCw6nBEXKvNlHrXuEspBbZqrUBA
vn32j2mwWeN0zjYGRVgld7VUlk6+co71QffhBrnmjX90LpzGJim9qiFvDusCLRWt
z+8qzj04JGBOCyLKry51s07ROjRHoP1Eef+YIW1fYdKBKcjDSGFUBrAf5wPNqFd3
hDM95XveRba5lRORHSxC9vE7OjrufBfcjvsGTro6EvOjG+ZS7PB11PHb2rSqfEyG
vvA2+Yvht82aqzckVMqBHPNKfWP9fsLMe2D9xUhbudatGORcn/3zA0l8cOhGiq3d
xqa0MxsbVquUhCHUmwy5Rh+CDXHbuQnv2RSUyhB8wUnzwV4QNztJQcGvfkLdiD7z
op3SiJwdFUj+z521qj2LHnYqUKPB0au+bd1U0dCflLJhopZPnsFo1Eax5N0BkLRN
c9d01YU7dhigTTna9WlpyBmY4alpup969OggfTs3RMFRu/mJbC0sWLve94fO6XHc
y1wv4mVEo2KFQ0i7TRNRJYAOEJXNknMwrKy5vppJsHtrj4rNTKUHxPCUf5B769Ml
yNxQ2MUAoyyJio5Fnj9BLl0gFmdLWJd7UdB3FHLuDeilWAcfl1OQaAZeM3xn5Pse
EHD0qY0JZb4BRHzqorvu5/zSVC+GpHB3+6+lP778QWqjtgpTKEqVEl97xyLwT/Wx
LFnsr31HsxLnycZ4Ul4WQr7uLl1CB8Qsg543p8yaT9+eD2w/ScaP0hn++3JYUVrw
WEp5c60R3Yg6lc58z3B4IY7AfPopQsb7nGkVhYgLfCMq+bdKhi2koPRN+IjyTmB8
Eil495bi6jaH1hiEcG4BbHDeuCw8QDZN0uKdoB6pCAQcjJNtxK0xE0QYh1xbeUwR
NXSG6R7/pt1mjGlt3gxc7ym8jxHEClWRr3oI6zBoQm6ztyAMh29zSXMMlllcuPMQ
LCMxOTElG1tmrXLdx2EfCQeDzbEagvV3pzcBZQIigko3tKDGh9q4d1+bTB5a97pD
0t9iA35i+BI8a0QgfgkYkBT5JuuSPiBlCuQQO9iCDRQqiklm2sgaIuxfpdywKIX4
aWonb+sXh5Vl0h3gJSu1fgEHZH7inYVljLbHsj2VM0eWlQBw5klaWY7n/7+C1cJ1
4RKMQka63BECmIPkaISrvG3u/+xrsgZtv6sSqEHrapLP55lqDU6olFEFsbPkoyIx
pZleLK/SKOXHTfMUseZFg9ybE0wddmlRanwIOpXx8MsNQSnA+vto6JcK1OqiUpC6
VFlVpifmTbEQb1s0z84dfXDtJyeLTtYmT72hDpIsEK6TU6qLw/ISP8lWH1j8i/O4
i7De97xOQ73z/mrLFIUAlt7moWgKkK8XTakvr3wta/ihIUXQ9ySXn6aaSi5L4C3F
j7Hz8q3Ri5LaXyosI3+7TA12g9Xp24YPIcq8ZiYCSEvPyUrzpbCEBMB6B7z8V1dO
6O/PQvglslGBk2VbGysRnY7PNN7qTpJ+rko51Pb3YS/8LIXjqjuv/30TPiCiN/ms
k/iol7Pa1e8PYgacYSbDovcgxmattNec2o5Hxk8yTN4+UtqIw8fy6WvEVyx3ExmE
n+wDE8QHHP50vOXpvziK+fhMhQwNDUHz6o7zJE3eU1aXBg+c8JqX8WF/smhTBu1R
/lq/JhM3cdgKJpT8ahxQiQ0AaDMVphYJmVskbiDNxFrCwOokgy67DO4ypmEZ0WDh
txx3MHsmOTEMPRQiCyi1HZFD0PXY/d+QXPClgtMplRhrsrNshu2qFvMEE/V5QMlF
XWJilWLi+W64VSsFGwlnP56nSBmUYYUqgXlfeGmGCWXDFhpTWBaJU8d2IPobAHQY
r9kW5k88zO9CMCFpB3mnli6Z9Kuu+d5wGLWbZmPcDAdVe5kNNofJj+jj2TXsdrcW
G56ExsP74WD48Rgc9mqG6o9UwoM9vwTpyYsCKZckHVInsQBk55i2/SZJ5MaF9JEI
xUAD+IysHvY9S2PhSEeiWllH0jSF585Y0W0aLSMwnwlZ8K5tefmoMiPHsnMQCxON
X2T0+cJmFEkB9SrLmDrzYrCXm+U1se9ZSzHjZRJ3t84KufwKGP0ku2E5yOsGaylV
VgsrMbo4T7qHy/RlxCgGaXn+228H3kgJdC+UzJtVqoej/M0BrV3XHLgCDgp6MOEq
NktR8g9hCMXz34pu/j3XgHc+KwKpwH3mLaRGY4ss/R/ekBLjdPz8l6yHF77mIkJ4
/9p1UVG2cY4JRb5zhXiqhjJwUxs5b0qOrMVBEtH3wG303RSg1fksZBUC0iPhpqhT
0u6XXstZTy1azfvhtVb5sqzjguRzjqhi8inDyuyXRp/0Xg8C9rWDLZUfXZ+Sgk/+
PyPih4yGQREUkmHNkrMztywd8zY08/x4m+TcPgUqd+T9ehZ7Qd6jnk8ZSkUx5L3u
Bty+uI2lmlzVEJwYNeDJEPm3FAqQqFhPWalEnpKRDnEJ3WYxN5G9wc+n+p3A1JCi
WrhLdpvpGH/Z0ax6tyUDohkCMnuIyes/MMwFiOwmSQU04eWN8M6GiIsb+CBzqWnT
JS3wODQnTNz82uWa5xL9sy1N3Mp7Shb/zUoUCtK7V5U3FxQa4+E98DMbEb05+CUP
OmXZvP+FkKv4MbnvP5Btj/smj2aHKItT167A+McuNHYuata4cnOZH8t6pQzkFyBV
ax6u2TvOy7v2ff65q74NL6IO6awIKFCgw1dLfjYHEcHvgggqKYJ5DeYnMh0TVh/u
axfaMOuWZvSAS9zu/ha1W02JUIMJOt/ujfYfg3/zd7Sw+zeYoedj2cCODVemzCHq
T5k6ok1oq2zECIogd9t8fUFBGGiBruEbM6d7tA9dbM2QW3hZanehvDLg6o3IKXow
TZs8Y5Lj97N4SKLohiTN9t6Uccw5UcPs6l/Aom+sNFa/vCwL7eGvDsF0A34W4cEG
bINsH40N7qc7FfPVeMmvYD9NERfI26wsrc9o7w9ztojb3W1+OX/Y4DjNkYaoE14C
xgq5X3/1hF/3rKCaIt/kreJW+ImERyNhUkQFNwQBklDCN6H+aGvWEj10uVzIaCWe
UZR2tJKg4cN5u0Vg/rGNt0bRJrslbbGMRdcYTlfnKjH73y6eh3V9G7Flshs7lb4R
9k6UXgAcpobtNZEQW9Pnqr54KaFB05gsgxocf+Uf6dUvHWZWNaiix/GJQWrCrL/z
35m7nJWIhKJTPimSLjfU9KpzDtIA8fLIUvGUeQaOuSnFAX2DOEYDhBR493ic6ZBQ
cqYjYCsIm1JIc8bMp9Ow4+KuKFbQkSE28J/7rbiBXBZ5IGnkXIRGLYaxMBO7e3A5
b5o2Xls6gUrDgORq+aGjx6XZaRa9ZyQCwetzhS33gcGEm2Z4NPNRUoVT+5Bsxw2S
4sL7Rn0q8eli6zqqr8XqQ7EkjH2hYb6HCCeHoVCEUM2Gji70yLzznRI/UQh9SqF7
hi/+tJWShDXY5VLggKfx9yieXOST8i00XuqeR7IdNim3Y2AZako+MlLJJLX/5JD/
pZhKWeg9g2CTvaPh/sBbgd2zbsIfLpYtwLyNK24JPxdGDuP4RKdYrfYwUFk1QK2A
efuKbOkXdFa+HXzzi+IOKC/DtsR0Jg85U9k+wSrpQ0O8vxj/AyLo6utVChM96JD/
gX2JCRoLqgVII9sXqvtqCYYLQzEMSnBQyVYUbof0pnwBBMJV0rXqzTLk5CE2kn0E
RlHjO/ZkiI2Q3hDJHIl/eYbBnZk3j3ESRVCK16/8lwhejG9jviH+gAlFLD4jaaEo
ffQnL4V/XBqek5LkLakulFIzQMueOoc2vpvw1bsoCC2P7rsJjNBoEPJX13SPYkSG
Y/1t18pPwhBvW7rS1prrcyHGw5Cv5jpLxOcyC+1FbeuyGybUFbm1YSwl3Pr6ROwz
pB/adwFXVNyPfc6qFHcYbyvNWzvaFKRxMLyV2xoj2fNRjRmMHCKi00bmf8R5J+CC
G8AqXQ0HoUigipUb6eAD1giA1gUQJ5HaKjkDn7DV+pjyETakn0DGplXgTMFTpDkC
WoSDwF7IQaLlu36JP/0Gzg909HoM0S0hSU/6kvMfHyYduz7KU12FcGBZI/CGxY8P
WwSNCvRNxpIgT/HmNruXOOH8BQryiiyMx1BtyfkMOZpE8kHCRkJZRQZh/MNtZmWU
6OMF4nKTlwuUo7jKoDzIRSaPks97RnY8LC/aex00Q+WA5LdMMeuGWQoMxcXvemis
EAANur65tlRhgFDsSjje85skSbQTr9lMhW5oNhemnqFTH5JnzBadk2g98ByihgSN
2JxWKwGQtfon/aDVQh78qWwimdGrevKUzFLbPOhbrmee/3740LDxHTf/Gwcjr40u
KU4CeL0D4eaTiGbLbcz5dvCgU3mvuO4lAOZi3nzFDUsbkSt4I2aLlyY7JzEdWBEa
x169pcJf1xHdzZLVpwQZwnhefGOdnNYFW84dl24vMG1YRKT6kHxwMm7V+9JaNGmn
8B/VgzW4wXRf/DjO1ust8PFkjCyTbZBD0hu3Y1vKS+prJnKRgQTlxSDwVr/ja9NO
iZ9vzLxGxeasZ68PVcf6D+KQPLAQ4uqivcFecY8nwcepma3ORy44Yw9QNZNIZ6vE
f3617m5JsBju6gaTE5zQDOrqtPRb91K5rUbRD6IAmaICOrrNXBxFSeP82pFjX4Ma
Jm9fIHGFLQi7/YX7YWteJgoQoTPKvCqE5Vd78LCDZWJTfeYmQk7OtaLZoiO2lxXO
Z3ag1A2R8+aK6d6j1XNgswnBD/hLV2Uce0GKjTpF/USsxIaX5mY6tIIYEAPxK/Ei
f3vrLZmNeF6RavCeAgjhVWNZ9zU2cUJmiev+SlpTiRRErIeqf9us2NIXkDIVZFgs
yjlI3hLqKc2JK4AashptlKBB5BrhnttmToHcrIIqYy9ckBOpBWQyCbUvIseclApz
uGohygD+pDapo7J9UGeSqt4iC5t9Dj8XW7VOU7+yU0UzWZIFu9wr6brwcDpZ1nJo
Gd5ISRcVhqNknTxFEf43h/4d6XhiX5Hz6mZlQgO9Mz+/hKZenCHYL1iQ9nAPm5vS
ubSzzjd1xrKoXuwzvpMzKRQLmTOmqvSeLzongE3ZGlwukq44JC3j3JdpWFUDugHw
8jnO9KqR8OYzPT/IbBZOxoQlLjkSCrP4KjwKZrplB0DvR+/wkgK/FdElEKzHhfW7
ci5tEIY4hG/eR+GTPtS+Xvd1Z+hoTgaEfD3AgloSCAIpx4xHEK9pDvdPyigIscZc
BLvpeVkDL0YAL5CTz4i1/Ml7kB+p9C3BOvk2tYVoPyw8C2G3RUFoZcvRLOR8lQaP
KzfSb3TG9FyZdHZRw/q94MHRFCV+4z/acciALa8yk+i7N8JldozAv7Y6BMKPjzXh
7bMzlM4SU4D0zeD8otXedIzJ5rYEonIviT6l2JfI/5+q4IISv5tvVB8t1YfW3S8m
FGT0hMuUEp3777vQGtz3399yWeaa6IsK4z78hn7kWiHX88ObyYb2+HGrrptAGFln
fQw30BwGoI0UWlm/JOw0zaB4sQcCCIQXDWk553vyDy+XtPEaQnIw0bHqcIIhGqY+
mGh149rrfAOjLtkRAG9KzIYUnXlie0SfjYzpTr6/f/MhqqOX1NGQeVgrI8OHiAxR
jBGjl5BBmShRUJbb1hm2fa2RcT+s/u3MOwNs9mtY6u21pQY+VG79Si2Ahz/IvAom
a06yrdUMTVjXnj8tqJuqp2GmmrzhygBxju1E/pLEGILLZ96bZ473SpRTqyMzbWfV
6CUMBgTWBqx6lqGk8hxlCa9Fv1w8lE+XiaEWrXsHgTG+dUR/36qFcJr+1UJ6+aj3
iXtbxZ+xSFkymfsQXPkKkN43RjkfobFwERoC9Gnv884tP7XQDqcepHX/wRjWtqRJ
B00wRP4tCx/yMiyqfEF2ZRWwmc5gu1AqKwLugLUSH/NWPS0Blt1vcLUvfJFrUcgA
GXc++wXrgJcmQIPGz+sNN01U//1RR3wl9bWck+ZIkQ553nWjC4Pd1zGWAGD768c9
6FNbRPGdU+sjMuw6bGxM+KnSR0M89yEaLDxpylyjC7COsMRUPz0l5pz50ZPV7J6b
VNbgjQ8Lhv9qNK6uBlO+8vwQQzB6P4XrzeXR6hZ3ezF6mha7ndx1kx/cNSSnqiWX
8KyQ8WBD4hJy54qizK3m8jnd2mcMXOwT1O3HSoA8bO4U1TWVqB5NCos2vDO1lNDd
8iU51rtWim5FNt5/yL3sc8a0yeHOyiS1SBqdCuYIJY9GtuxZRoVzUbUYDT8TNYyi
EL0lgLQuWhWddTs3IZsyNSJ1pKCTTdHQG+18LvPrnuNG9fzU8f9NyH3hmU45fONJ
Az0m5NbBv4Q2Z1Lr8cCVipCDdR6DTob2QKPGQI+cvXU/6mZmRsh6s4jmMS8XTBYo
0+9KL8cUBQwbgpRq/apJ40ljS9EYD7MrkuWwA7Mtur1qw0asRp3RcQ+VgalmegbK
AJC6Ei2dAA8nhdU5bQzr8NglxbrirR8cfqZYXugsXa5WbGxhuiAPMVHaWUbhCcwF
FEr1BElq1HNMOx9EJk6zGHOzFbKYDsTtu1O1CNGkMed20hbH+Iic9bS2ORkLtdCk
1Qpt6taggKHfNH5kpfYxPAQcoGfFHjtEHmbvW8K9AOsIXm4RpbwKTtwJUSKKG8oP
Bpv9gOo1BP0ordMyoZGbE0XQwn5X/T3vZ2u5hYF7X4ddCOYVeltLpGzOSg5yd7bb
xtK/o/xCAqR/1IxwIYSkrcIGDSjbGbdt8JWkN0lhwG7EjgcBTKvEN9kxFIhTxESz
4qgtmTwldK/VejJ3m2EflMXZGNFyzd0h3zP8tg4QXCNMDAoKkfo+yhGHAAUtEEia
GT4yksmm7pb/3PiiJBd5RjU141nakiiWlnGUxh0HQmfMvjgfja9n9SHP4tW+w1Nd
oVhRZV8re6t+D9BLDO54p1qfvp8gfLrhmQDf/4QMJMATesmN3SxCVJ3LXIuih1SB
Saf0WZHmZDbsA67avZFGIoJyirgfUNmAqPdPW2Uq5e8Z+vuHGkFklpcSkfdd9v8L
jJcuhYRvS4eNLcBrPnBXSaqNYcygCZtMYhHb+ycqh2iINmxJKKknqkpJu2wlZzD8
X4MZBZDvNm+CrWH2W/FhhGY2iM9tKAp67bkrSReTq9iR/R4JbTUyvbQnb9+A/ipB
jE2fIriXhKiGlN1vcNy7wmILd+BIiGFZEaDEsdldUcrGa3LpkG4DphLwbtlHfdwm
VDEQj2+CjDsrJSvJLK66ekyoM2LaIPfe577p4PNrpkY6HfZ0WhzNhnC4jYfM85AC
aMf+yknWW0DzR++QqK0D6FxYfXNgfLZkoRri4rgQQuONTrFL8sg7D2x0dNFxkg3s
FGwL1btljIVfGBY5cDKKcdYwj269oEF4k/leemHzZKSVeqot9FEki3VMgFnjlyV7
mvbCkqNV+q0HTDH8wgu6y4jK6FxL8u5pGppKdC1qKlcEVxDkfD3ChBLZYH+wDNO3
zFJ6JcW/+YL05d246bO2lfIgrzPP4gIL5jgyYwpKbvVifNSlxc5117Wtx4awTNct
EChILW23P1ULt1D2nhzZWotw2J+uengOqeTNQ3/VJzAiTSwjPR7Jf2/XMMtJ871O
NQ8i8HfImeahdq8cDkih7zBTX4zeNSuh+S9HL6oZaONE1h31v8JiC6orzWqIoSsX
GWRhQICPxWWgRItmcg695IZC+oRmx3hxm+08YCXksEyI3zLucGRzqqr3qqQ5z08e
HthRAH1aba+/nxWLi4gRkBvMcyzWIxzCgCpQz1mslZTfnwenQ2WiTdAnjN+mewmS
L4Q/C7dAxtb26ZRCGtfTBuVaeu6g3Hv8FdOlcg35Fz6+VghdoaxZhehTfc5S+SIN
6ew8tDMOFQsGCcBHIRNt8KbDrTzKTZnKIymrFVB7LiyhHU/NB8ZM2onGhw5vp5gz
BlWfFN4GqJsifafery61rVudflP5GwwCwJWCrBvu+GGpMEG/1K1+1TaLCjw6BCsx
Dp/4lubhybMpOOGATuP9BB27jk/NSmVGrQIMVCnGTHfgK5GxJDj1U5QtOWmr4W52
aADgQl8Q68BwUfE9FABOBWdMVYrQH9G3VAoLzXhP9mWxFhWit2cSR622ZsSnSbyY
Zrb6x6/bK9PYtW88UGN6bN8SLbcNHWG8mPZ7W3cdUDhw17/yBJMCaMkHPeqwQqvx
cyPCsIq6H/B0FfWxP+Ty6cYU0P6jdxgWUAA2NIFz+PI=
`protect END_PROTECTED
