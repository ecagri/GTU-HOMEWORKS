`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KudbeI8SfO9g+3NJQzNUFXzOUAyVxtwNwwAGfkYRMD4yw9Wr3GJhxTVa0QloQhjk
NQHq32Ki8GAwd0sEvfNbB+S07AV7Hy289x62JzzJ72T90hLMPSOrIJcozVSlhPDt
dCRStKMoW0DqVPCKLps9HkzgQbhVWfsbS8QGCfeXfr8omkWopvGmWEM0X0hcjWuz
5IplDFy2X9D4buvEEsI61IK9LfMzJCmHWh/GVpsT9gJiUM/4YCkQ8TzFBKPW92/i
O/Fm1AbV1reUnaU3yW1yl9pVum3z5lmV320WdgC0NBQADOE3q/oppC765dxAwCt8
zP99qkxBzk8NjYbQkTxzucmt6+POX+M3QZqF99HvwxLFKh7hP6rTgNoadwLnAtGl
iEp2wBLGrNkd67wes4JoHt6ilpx+doo01xPIH3SinVZqsqlBGSMoiOAFKiQ3YBA9
m5Xkp3KoKivt6/Os8+aVQpmyfHIv4OYi/7+srHiRP+g6pK1HHVDLWavKZwBiy6B8
v29Yh//Di2xSjmhoSPZFFLXRAol8Y8L5MVT/jpJY4Iur9fCuags8hRiyC9LVYPwy
eTBEx2kIfy3V7SbGxcLeK1ymJpcgpdN+yvznYoC9SDo8+TmxZR7MRrzS296Y8XLp
r7128UFHOWwo3gtqNL1WVESfu+H4+dQCyjaUv/y8suXmvVRbB652LZWDe4/QjAT/
USx/MoH4JZ1uMSnbpkLH+yX7c5smMj4ir9C0S8fi32/eYSpeGQIhyr06JobgwOoW
JAUeqoYgSvpt6O6CuFDTjpOXkk9+HzdEI4+1+z/kDLc6W8pPoEB441MQkD5T3jEh
djJxIGjo1lyPiM7IT6E1Ad2n2LP2WyrJ6nIRB+5mpk/hm6ymNhZ/HV54WNCslLs+
DlMe2YZAOSBVEoEnjSkn9Xya6KvuAL6gfvKiUaAd0a7D7X5iRijNOcYt7WdWV2PP
c+3VHOCAlUpRR2N2iMhSl0o8z9fzbqyI3ZwqFyj1Mqcia0ycs6cbAxtABqCSW6nr
ek/IWsFbW0D1Ni0sxw5E+forjw93qEHetbhGAvlSz6xeldmMfTTMXn3kCjSam9t4
DVfS4jlAw+WjMTyU66hTUsDMzcQVXB0fCDZsteyzinisFMpwWAV6TnDt9sBjqZDu
PcC0Tww1FnTYRwquqnfjJ/U7fsUsjwJ2wel6QisNtwQlo9EZUdZYxFii2pLAop80
AYjJ+hZ7VjZnznOFGDn54xQeDgE9sgZCKIaJIYLpL9pVESTz/jsu/vCTUCxNidfK
cPH6u7EzS5AZrUKR+XLoHSdZQFjAQLQuWvzNJZfvaW9W7f99vcNP3FylSn+ipkpO
8X7t18TEmIGSrcNoS1JMbD2QSJwTV99/50av1bHgyupoh+CdjgKkroNrWxSs0hu0
XyQpax6dJMKwpX1GEgVbjnXdbMCTEziNq3MsPVxlipXgsNtHafRbapd/G/IwOI8F
pnIT5ik9Y89+9SkFKd6Hc+xnjLQ3vWXBXqOneouJdXZ+GL4ljC8gvbHX94oSjavi
nY5pS9QgvGuZqrP+AuyDEmsJKGv4mUvpWQ7cBuiEbtZmh0eaWh53HU76Ep+/sdpC
nLd1dPYrv4qnxSa6HYZ9tB/6eQWlUfqkwP29YZ2Sj0E6fdEIEgWeUPdsikZEFoPf
1H7vXZThH5YW4f20/p/+eWxba3kbsC8m5aCj8JwVLMMTta8H28inLuB/Tcbp0g5j
FpOFqGI7fmTibnipKIYtvctn23Kwoet5GzIw77ei6Qswij8+RU0IHlsITIKDYAyC
vsWn7cvRT0yn+qL4BL/Xd7Ct0NSdtc+pCMph2ONexgzK4flmyLQJ2OFTWZe2gR5Q
LNvrnAid+S5Cyo7JSlX264r7wFU7ZsOlpj2UN4YkpxYZBNSk2BeTORvFEaK2zwB8
YJ6D8vhrqbhaOez2Eet6NXMRYtSX/cP/64OovYX1PIMwRc59u0MqZ/JLRJLVWmCq
EFJebamtxMo6bpnrurzV88uXvCbEokDD/xvl1e8tYlPMxxJKaQAZIo5eqsJi+YOM
PvK5EFg5KbZK/sk3LHvQpnC6ln+EwyH6x6BLpOJ56Y71H8MuNWtjM9fB932AwK1X
C27tMhy1lz8CfsYVC4fwsEdBFIGGOipCOXmibEsdxihkhubRZoC/1funGExWn2LB
CmJ4wnwl87peamyG8UDW+j046N6r+EB1iB7bWQUHHkzS2O7NqMJFRtLsMkPmvyrg
5tplBBx39I1aSj0z8ZfrqFvq91/gTz9MyxbYIiRg3GnYbiUSvjsjpYFsK6jydhmA
81kpBcEb7WtdHK3w0n+9A2ObTlyntiIuzKmzW2s59J1fuxdKieDSQP2YSkCUi9Qt
IfwYlrpdjFCyXQLuzt99WH3sQ0qng62jNMPPaKwaYgXxoF7zkCeRrL7fRfZvfqYu
gdVB8Wt3Tu38c8leXcm4Y72zTE0yMVRFnHqOqKPWq/GoIOkDTm6euBYmBZdiZiEv
pce9NPwfIzyELZqZ203L0MlGc71vN20WJpWPjoBMRYwJb5+XsZrSz1ElJ/Mi0+Zu
WC7AOiKkk8J0vFW3RMURGR5ZMWZoPAe2RAVuEsdTDPF5AX9zjZWqfF38BNdmNhxP
PAe6HnH8tLux8u3ypTqzaxsY8zYZpuIwyq1ZDOrwrIPjOLFOe5bwnpyjeVe9y5Mw
hhFotkTaMZjUJeoa7zVKtE/7kPumvLte6wWV7Itvu7WxhiHH0jhKImw5qeR1sK6Q
oCQQc+QxRszmsS0hazSA0Ted039ZYmseP8h/+vHiJp8kaCuzkxLjT0+uvoZDs6NB
XlgOpChd7fxI0fW7T5C1AO8YAs4voLeY1c6DX6eXTWJE1Spk6bR5kD+a0jdLNABq
WUz01Z8/GUVBTSNU2kg8+9EEOENjeMI7TUA/nwV6KfliILIZEz/vH7ORqPHlTySB
Rj7V+ONpa7/woMS9Z2kHYFPsN1nC57oX5fa/WyQ5QRTrqJa3z+/yXAtEdnYggtSh
XnVxlqSwTC1GBC6gpRQSPNZ/ZDxTJS9+gXMiMU3Ep1vTHQJ8WQB11IjNlUJ3+V73
EmNjHzJRay4mKdtuRSaGrSRpi+HDhaV0BJVD8vIZOW2/rRF7To7X0HnNYK+NBU+B
9LTdmnm4U/GMLor3Cl2aFPcqZzjSdsFtO/BpHxNHqFecJTHmP4Y+3huNgaXU4tjt
TQ0Myw3lMOmxvDT3CDa7NgWjH2zf2wAypVSZHXE0JpOKdJMppzgCa1aFIXXwD3dK
MiHhXjaLJHsqAENjKuUUY4/82Ki28b8s6pOCzVl6ySBU3NXNhZYZNVMP2w1CoTuI
t8R8sls8EoAQnMcQcC4bKwTB+PCmmpLZTd+PmgoSs/Gw3SzOE6odeT7prIvKKhwX
LuURhkeJs1YVIgFyr5I8i6/K2pE3klLjaEOOj3eTsdAZ8vwqKI/w4EVmTq0076YX
CA2fT2sXnXpDE8MQCMhHXi4eMGyh6qu106aU4JzC5dA8Rc5Y0aKj1lvKNa8298eh
ywf8WCb31GrHGJ8S94ntfKXb9kZFUER6+DkV4Pm/2RpAGAm9kAR9J6bZcuJ82/qn
/95DxJCYkE6TKEoHqU2GDN4P2oJrItiKqvtZyOpSkbvGmnBiPrC55OXP7tLR65Jx
LUnI8J/egnJ+YHw9Z2vrvMA9IMCVeeFwoAw2byMhzTum1sUX1fuCTxQJAgS0SmUP
peWwUE+C+jpUTRIgvBFDXg6GvQ5FM4oy79LYZU0YEGfpQuZnlT3WEv6csUjV2knV
jncus1Elj4+hb9Cft4gpMn4qrkMQkRua+XIYmEfP+RxW69AO9wr2grsDX2GyvFua
nJ7kF+iQSrjhSd10ZBGViwMhe6gUpaxzHGzIKtQBFCvdxIi8oLJ50EdnUO5TSeFd
V6dfNOgRfBfJl5W1WGYLwrbS01v65pUTgwuvJVIncMM2jsNQU/L4aoEn8wTumBuK
IK1+0uyEMT5ErGKdyYc9U+lXo2c9ZdSJUFjN2Yp6NQaabZSfP0dqMoEwEsd/qNmp
1h2Io3QfxWSsVteLlOveMxjJd+HNbByRbSS2UE1VOV4=
`protect END_PROTECTED
