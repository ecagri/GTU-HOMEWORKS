`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7uybn1IOHGeImoXDi039HkwRGiW98GCNPt6qX4fei5rXMgPLh/nfyNGvbPa2yXwK
MVUo//wt+jgCYmteNf6E1pKL2rK7OeMRLqBg4Bt0Jm8VbpxEyYtDZ4onz7xIcA/s
61lrWqLiyrP2OMNONrLu1sOlVd7z+bVja76/LbhWx5zyc5yz0TiFW9lvZFhuFQTC
2UHQDlI5FMb8TUhheAWPqPSYHFBezAxcQRevxVfg9KWrcrKNWMUBOONRZHo4qb5D
WoSi6z5JQKY1cAOhxAzxfPvrpLAdIKb8q9pZYkoeTztbzhICAVMgbIjGlR/hy9VA
wM9q3/SZ0oq0WiX8GirXd/SYGU8906qybT69ucaV568uAjk3JgNeeOIhg6LnKxgH
7TMsNKc7fBlh2AyvihcnMeHHkuAZ7whTIBkMvkhp9/Zqr9j5z1sMEBB6nn+Y7HS6
FMfy4E/Bnwu1P3sfm4/AdMLgg7EnVoW5GMuabdtoyLqOu/Lyku35MspuNw9PXG0o
JXyEKIrkOfge/z4/uU5zjU4cCb+K01bOCQqppC3Qkii28P7US7i94Z+bXZh+IvxI
2JRemJvtYePxjxxjaRBcv64oWskiMWyTIh3hUn0sksrkwxobk8MtC1L9w8h2aqkO
IktlCQzeZiXnyrE2SenzmXD0tlgfq7kCgeLYm7ye71L4AyYOVf5iBvCx4AjurqFs
DFro6S3XUi01EfI/e3YjXcW8VzzmJjDHcRgFtmLm+U/mCgYRSAir0Hbs5Wkh+pmv
yJmNvdlfsaoxZIKWgAkF+/dT7dSpecrrX2QuusGtOlhdFiTpZLore70gc6ZzWylT
Q8mL3ZhJ4BPByPdxyJ/lwdubHKllVMcOpk+h18rgLnTANiZyzskaJ6CUyR7NNb8I
LvLJS5z3fR5LBVbUhxlTqs9M3JBssRZdjcSNl+pai+Y=
`protect END_PROTECTED
