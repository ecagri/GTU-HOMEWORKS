`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
odJ3huJNk0SNFxPxEBlicHRZUBCe3Qgp+5yyp9R/z0R4VQzeplOgknFHvmeRp68y
PJE1TXiCfWtYmfOO4HX7+FDP/L/k/H6xrnkTlRhKi6eeLrlYZpJmOutDq0AKqZJ0
dhsQdRMNV5eav3uNhbZSv66vr6CYcwaeeSsBMoZzxj35/rF3B6aoySCWElpBWmXu
98JsUaDsojZ+pVgOgZirjkQ/EupemfRSUu3mgN7W6KxqXWjwNi8JIhOI+cUheLPy
TG3ubTvctlQdFjXRHyj25Vn3TUR6NkPFqz90akw6xTexWB9u5gpt4rsYOFfUPaxH
wuEIKwfZezTOe/JxyPiM/vEB+B9SOT1YxSxAw/8mBZ9KKRBaWg2eSibMC6gQwLmg
ygnHtifOej1IPeCHGclQ77v/ScJJ3ASHyVBmu6HjX+UOeuoS8lzC4KA6NUCKG+8d
0FtENyBYyM/cOggV4++u8Ljwxpl/x9Svb/uAaspoX22NDnGOHQ9MwHuGcmjPhG71
GqLo/uHMUQA6U/Stjo/zFSVVH/Or91EyAUV2sXJeYDucmgHVA4KIFdk2+4N817gj
EIuhBiWYAohO7CNBmGGuGVKYRsOj0hdPVNICdxIhP+eMW8OKrN7JZh6WEkobXA2M
tWJca+IHhFkJEuasG/Z7WFi3hDK83qhYecyF4ukE1BfLuj56PBwu+EdbjNfqv1zc
z7b/LBOQocdELmtc4UM7WtKIunvOzJQGoN/ONEe6EaGUiDp+zXmvJNDebmlICe1F
VAT2iof851JxmY22w7xJuo/I7Q19n3vj6dUbuV/rf3eDy/IRfrtQnlczDXL7sbn2
Mj4bsR5Ccy1g8l69QVILcI1KnD2Yae0i9oVscrYikwUjylryzFjnDC7dU/L1Bal2
LipnH6XLMgYXtnGaVoBzNZIWNtuW6o4OcN7RS3e+ACztT/epNov+4y4gUXlh7TXh
6esjwTdG6K8/H3dEZnV4RzDBwEVoXcVMjAK6F8joMS9O/TnVeUCG699grRkHFMd7
L1akTrqpmjX9fyQRuQ1DVrc3WM2iHtAMqTujJp4LeC3goXIAyHHhaVQJSqLEbfmB
FH8p5xam1k8kP+zI76FlcuYZ7MqHK2X1ABcr2J39sblmeB8NBbpxNvve8aN2AW+Y
erTj17772M2J35rsV1XG0Ib/WQxezHS1oGkno2+qkasViZNacLm+N64xZGsm5Mr6
cmTUZeKyBhD7J+4JtttTuyg9xry/2HVLBS/0hJKKj4flS8Mu6SoDju4AU2QGQMMb
whEXYzae0YK1fTOiQENjYi1hAq/Kmqb9y8hqwWL/RQfsgJbU7BfzOTwdQZU1bFn/
ZWAIk4yVNAYtr1e0GYBv6BnlfAgLbpcFHZhr/vCpj2rSHwgjNFAuETjjqLgsYTLY
MY2Mb81/zG4BHgF83rAPWCpOITPfw+LGnmJo9SryXCm2vdkG2+I7T06AtOSkcVP4
`protect END_PROTECTED
